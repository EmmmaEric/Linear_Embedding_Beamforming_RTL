
module memory_rom_28(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h35ebbe2a;
    11'b00000000001: data <= 32'h3107bae4;
    11'b00000000010: data <= 32'hb4453b55;
    11'b00000000011: data <= 32'hbcf03da4;
    11'b00000000100: data <= 32'hbed1b4aa;
    11'b00000000101: data <= 32'hbc50c032;
    11'b00000000110: data <= 32'hb615bf25;
    11'b00000000111: data <= 32'hb8712546;
    11'b00000001000: data <= 32'hba313c73;
    11'b00000001001: data <= 32'h30233b6e;
    11'b00000001010: data <= 32'h3d4a3a7c;
    11'b00000001011: data <= 32'h3b1d3d8d;
    11'b00000001100: data <= 32'hbc2e3e78;
    11'b00000001101: data <= 32'hc0013a59;
    11'b00000001110: data <= 32'hb868b137;
    11'b00000001111: data <= 32'h3e75b4dd;
    11'b00000010000: data <= 32'h4034b2c8;
    11'b00000010001: data <= 32'h3c46b9ca;
    11'b00000010010: data <= 32'h37f7bc78;
    11'b00000010011: data <= 32'h3bc9b29f;
    11'b00000010100: data <= 32'h3c4d3d02;
    11'b00000010101: data <= 32'ha4563c7b;
    11'b00000010110: data <= 32'hbcb5bb7b;
    11'b00000010111: data <= 32'hbcebc126;
    11'b00000011000: data <= 32'hb984bfc3;
    11'b00000011001: data <= 32'hb854b270;
    11'b00000011010: data <= 32'hb79635b7;
    11'b00000011011: data <= 32'h338bb4f0;
    11'b00000011100: data <= 32'h3adeb4c1;
    11'b00000011101: data <= 32'h22e13c1a;
    11'b00000011110: data <= 32'hbf3a4019;
    11'b00000011111: data <= 32'hc0b03df9;
    11'b00000100000: data <= 32'hb9cf33c5;
    11'b00000100001: data <= 32'h3c6fb449;
    11'b00000100010: data <= 32'h3ca6b040;
    11'b00000100011: data <= 32'h32aeb222;
    11'b00000100100: data <= 32'h35e9b21c;
    11'b00000100101: data <= 32'h3ed63914;
    11'b00000100110: data <= 32'h40503e79;
    11'b00000100111: data <= 32'h39fe3c86;
    11'b00000101000: data <= 32'hbb51ba68;
    11'b00000101001: data <= 32'hbc67c024;
    11'b00000101010: data <= 32'hb3aebdad;
    11'b00000101011: data <= 32'h3425b4c6;
    11'b00000101100: data <= 32'h340eb8c9;
    11'b00000101101: data <= 32'h3779bea4;
    11'b00000101110: data <= 32'h38f8bd39;
    11'b00000101111: data <= 32'hb4103974;
    11'b00000110000: data <= 32'hbf0b4018;
    11'b00000110001: data <= 32'hc0563d35;
    11'b00000110010: data <= 32'hbbe1b480;
    11'b00000110011: data <= 32'h2dfcba0e;
    11'b00000110100: data <= 32'hb436b071;
    11'b00000110101: data <= 32'hbb003522;
    11'b00000110110: data <= 32'h2d3936e3;
    11'b00000110111: data <= 32'h3fe73bad;
    11'b00000111000: data <= 32'h40bd3ecb;
    11'b00000111001: data <= 32'h38e03dc1;
    11'b00000111010: data <= 32'hbc802e7f;
    11'b00000111011: data <= 32'hbb31ba51;
    11'b00000111100: data <= 32'h37d0b735;
    11'b00000111101: data <= 32'h3c82b1ae;
    11'b00000111110: data <= 32'h3a5dbcc4;
    11'b00000111111: data <= 32'h3918c0aa;
    11'b00001000000: data <= 32'h3a9fbe5c;
    11'b00001000001: data <= 32'h362a3924;
    11'b00001000010: data <= 32'hba563efe;
    11'b00001000011: data <= 32'hbdde3819;
    11'b00001000100: data <= 32'hbc67bcf1;
    11'b00001000101: data <= 32'hba6bbd69;
    11'b00001000110: data <= 32'hbd51b354;
    11'b00001000111: data <= 32'hbe1535e7;
    11'b00001001000: data <= 32'hb0043155;
    11'b00001001001: data <= 32'h3eed361c;
    11'b00001001010: data <= 32'h3ee73d43;
    11'b00001001011: data <= 32'hb3893f2b;
    11'b00001001100: data <= 32'hbe873cd9;
    11'b00001001101: data <= 32'hba6d381e;
    11'b00001001110: data <= 32'h3b0b3666;
    11'b00001001111: data <= 32'h3d2d2c49;
    11'b00001010000: data <= 32'h38d8bc91;
    11'b00001010001: data <= 32'h3821c008;
    11'b00001010010: data <= 32'h3d49bc26;
    11'b00001010011: data <= 32'h3e4a3b96;
    11'b00001010100: data <= 32'h38873dc7;
    11'b00001010101: data <= 32'hb8deb276;
    11'b00001010110: data <= 32'hbbd0bf36;
    11'b00001010111: data <= 32'hbc39bdf1;
    11'b00001011000: data <= 32'hbdc3b3c7;
    11'b00001011001: data <= 32'hbd75ae04;
    11'b00001011010: data <= 32'hacd2bb58;
    11'b00001011011: data <= 32'h3d10bade;
    11'b00001011100: data <= 32'h3a8638e7;
    11'b00001011101: data <= 32'hbc423fab;
    11'b00001011110: data <= 32'hbfde3f57;
    11'b00001011111: data <= 32'hba813c41;
    11'b00001100000: data <= 32'h390c3903;
    11'b00001100001: data <= 32'h380533a1;
    11'b00001100010: data <= 32'hb5feb8e4;
    11'b00001100011: data <= 32'h2a55bc5a;
    11'b00001100100: data <= 32'h3ef0b0de;
    11'b00001100101: data <= 32'h411f3d48;
    11'b00001100110: data <= 32'h3df53d52;
    11'b00001100111: data <= 32'haeffb49a;
    11'b00001101000: data <= 32'hb9b2bdc0;
    11'b00001101001: data <= 32'hb8d3bae3;
    11'b00001101010: data <= 32'hb95ea45b;
    11'b00001101011: data <= 32'hb900b9c5;
    11'b00001101100: data <= 32'h315cc055;
    11'b00001101101: data <= 32'h3b89c012;
    11'b00001101110: data <= 32'h35d3a08d;
    11'b00001101111: data <= 32'hbc9d3ef0;
    11'b00001110000: data <= 32'hbeda3e84;
    11'b00001110001: data <= 32'hba3038ce;
    11'b00001110010: data <= 32'habfd314a;
    11'b00001110011: data <= 32'hba843353;
    11'b00001110100: data <= 32'hbe89a97f;
    11'b00001110101: data <= 32'hb865b51e;
    11'b00001110110: data <= 32'h3f1e34d2;
    11'b00001110111: data <= 32'h417e3d66;
    11'b00001111000: data <= 32'h3dc23d7f;
    11'b00001111001: data <= 32'hb3e434e5;
    11'b00001111010: data <= 32'hb7e2b454;
    11'b00001111011: data <= 32'h311e3490;
    11'b00001111100: data <= 32'h34ec3705;
    11'b00001111101: data <= 32'h2879bc3e;
    11'b00001111110: data <= 32'h3503c19a;
    11'b00001111111: data <= 32'h3b64c0e0;
    11'b00010000000: data <= 32'h39b6b179;
    11'b00010000001: data <= 32'hb4e23d8d;
    11'b00010000010: data <= 32'hbaba3a88;
    11'b00010000011: data <= 32'hb857b6e1;
    11'b00010000100: data <= 32'hb970b840;
    11'b00010000101: data <= 32'hbf573083;
    11'b00010000110: data <= 32'hc0db3202;
    11'b00010000111: data <= 32'hbb72b518;
    11'b00010001000: data <= 32'h3dcdb0c1;
    11'b00010001001: data <= 32'h402b3a87;
    11'b00010001010: data <= 32'h386c3d86;
    11'b00010001011: data <= 32'hbaa13c7c;
    11'b00010001100: data <= 32'hb67f3bdc;
    11'b00010001101: data <= 32'h39933d3e;
    11'b00010001110: data <= 32'h39b53b44;
    11'b00010001111: data <= 32'ha518bb1c;
    11'b00010010000: data <= 32'h2c6ac0ef;
    11'b00010010001: data <= 32'h3c5abf84;
    11'b00010010010: data <= 32'h3e6631b0;
    11'b00010010011: data <= 32'h3bf43c5f;
    11'b00010010100: data <= 32'h32cea29a;
    11'b00010010101: data <= 32'hb0b6bcd5;
    11'b00010010110: data <= 32'hba30ba6e;
    11'b00010010111: data <= 32'hbfbb3305;
    11'b00010011000: data <= 32'hc09c274c;
    11'b00010011001: data <= 32'hbb08bc69;
    11'b00010011010: data <= 32'h3be3bd48;
    11'b00010011011: data <= 32'h3c54ade8;
    11'b00010011100: data <= 32'hb7623ccb;
    11'b00010011101: data <= 32'hbd383e33;
    11'b00010011110: data <= 32'hb5a83e14;
    11'b00010011111: data <= 32'h39c23e75;
    11'b00010100000: data <= 32'h32dd3c83;
    11'b00010100001: data <= 32'hbb5cb575;
    11'b00010100010: data <= 32'hb8ccbddf;
    11'b00010100011: data <= 32'h3caebab3;
    11'b00010100100: data <= 32'h40ba3981;
    11'b00010100101: data <= 32'h3fa03b8e;
    11'b00010100110: data <= 32'h3aa7b56d;
    11'b00010100111: data <= 32'h331fbc82;
    11'b00010101000: data <= 32'hb46fb45c;
    11'b00010101001: data <= 32'hbc703914;
    11'b00010101010: data <= 32'hbdc5b42b;
    11'b00010101011: data <= 32'hb815c036;
    11'b00010101100: data <= 32'h392dc0f8;
    11'b00010101101: data <= 32'h36babaf9;
    11'b00010101110: data <= 32'hba973ad5;
    11'b00010101111: data <= 32'hbca43d12;
    11'b00010110000: data <= 32'hb0a73c12;
    11'b00010110001: data <= 32'h35c93c49;
    11'b00010110010: data <= 32'hbac33c12;
    11'b00010110011: data <= 32'hc0553359;
    11'b00010110100: data <= 32'hbd8cb825;
    11'b00010110101: data <= 32'h3c03afc9;
    11'b00010110110: data <= 32'h40e13ac2;
    11'b00010110111: data <= 32'h3f543ac6;
    11'b00010111000: data <= 32'h3947ac7a;
    11'b00010111001: data <= 32'h360db334;
    11'b00010111010: data <= 32'h37cd3ad6;
    11'b00010111011: data <= 32'h25ee3d32;
    11'b00010111100: data <= 32'hb849b58b;
    11'b00010111101: data <= 32'hb30bc135;
    11'b00010111110: data <= 32'h3829c1c0;
    11'b00010111111: data <= 32'h3766bc31;
    11'b00011000000: data <= 32'hb3f73830;
    11'b00011000001: data <= 32'hb51a3719;
    11'b00011000010: data <= 32'h34e0b089;
    11'b00011000011: data <= 32'h27a130d4;
    11'b00011000100: data <= 32'hbed23a36;
    11'b00011000101: data <= 32'hc1ec384e;
    11'b00011000110: data <= 32'hbf55b35f;
    11'b00011000111: data <= 32'h391cb4a6;
    11'b00011001000: data <= 32'h3eff35c6;
    11'b00011001001: data <= 32'h3ab23917;
    11'b00011001010: data <= 32'haf743703;
    11'b00011001011: data <= 32'h350c3ac7;
    11'b00011001100: data <= 32'h3c4f3f95;
    11'b00011001101: data <= 32'h398a3f87;
    11'b00011001110: data <= 32'hb4e1ad7e;
    11'b00011001111: data <= 32'hb63cc071;
    11'b00011010000: data <= 32'h37b3c076;
    11'b00011010001: data <= 32'h3c1db857;
    11'b00011010010: data <= 32'h3ace35d0;
    11'b00011010011: data <= 32'h3a11b6c3;
    11'b00011010100: data <= 32'h3addbca4;
    11'b00011010101: data <= 32'h2cd8b687;
    11'b00011010110: data <= 32'hbef13a08;
    11'b00011010111: data <= 32'hc18e3875;
    11'b00011011000: data <= 32'hbeacb98a;
    11'b00011011001: data <= 32'h3480bcfa;
    11'b00011011010: data <= 32'h39bcb88f;
    11'b00011011011: data <= 32'hb65c342f;
    11'b00011011100: data <= 32'hbb01396f;
    11'b00011011101: data <= 32'h33d03d31;
    11'b00011011110: data <= 32'h3d014055;
    11'b00011011111: data <= 32'h38144015;
    11'b00011100000: data <= 32'hbbc1363d;
    11'b00011100001: data <= 32'hbc48bcc5;
    11'b00011100010: data <= 32'h359ebbec;
    11'b00011100011: data <= 32'h3e4333ba;
    11'b00011100100: data <= 32'h3ea135aa;
    11'b00011100101: data <= 32'h3d7fbaff;
    11'b00011100110: data <= 32'h3ce7bd8e;
    11'b00011100111: data <= 32'h385ab020;
    11'b00011101000: data <= 32'hbb0a3ca7;
    11'b00011101001: data <= 32'hbef737cd;
    11'b00011101010: data <= 32'hbc2dbdc3;
    11'b00011101011: data <= 32'h2dd9c092;
    11'b00011101100: data <= 32'haa48bd7a;
    11'b00011101101: data <= 32'hbc3fb072;
    11'b00011101110: data <= 32'hbc003604;
    11'b00011101111: data <= 32'h36c13a11;
    11'b00011110000: data <= 32'h3c6f3dec;
    11'b00011110001: data <= 32'hb4633ed2;
    11'b00011110010: data <= 32'hc0263a83;
    11'b00011110011: data <= 32'hbf93b105;
    11'b00011110100: data <= 32'h2cec24c6;
    11'b00011110101: data <= 32'h3e493979;
    11'b00011110110: data <= 32'h3e253507;
    11'b00011110111: data <= 32'h3c5fba7a;
    11'b00011111000: data <= 32'h3ccbba36;
    11'b00011111001: data <= 32'h3cb53ab8;
    11'b00011111010: data <= 32'h35343f7d;
    11'b00011111011: data <= 32'hb86e3865;
    11'b00011111100: data <= 32'hb743bf4a;
    11'b00011111101: data <= 32'h2a80c13e;
    11'b00011111110: data <= 32'hb243bde6;
    11'b00011111111: data <= 32'hba4eb569;
    11'b00100000000: data <= 32'hb569b57e;
    11'b00100000001: data <= 32'h3b56b771;
    11'b00100000010: data <= 32'h3ba234c1;
    11'b00100000011: data <= 32'hbbd93ca5;
    11'b00100000100: data <= 32'hc19d3c0a;
    11'b00100000101: data <= 32'hc09c34d2;
    11'b00100000110: data <= 32'hb2cf312c;
    11'b00100000111: data <= 32'h3b993683;
    11'b00100001000: data <= 32'h37b82c83;
    11'b00100001001: data <= 32'h2d01b800;
    11'b00100001010: data <= 32'h3aba2f16;
    11'b00100001011: data <= 32'h3e8c3f3e;
    11'b00100001100: data <= 32'h3c9540e9;
    11'b00100001101: data <= 32'h9b7a3a56;
    11'b00100001110: data <= 32'hb630bde4;
    11'b00100001111: data <= 32'h8334bfae;
    11'b00100010000: data <= 32'h3128ba13;
    11'b00100010001: data <= 32'h2e3fb337;
    11'b00100010010: data <= 32'h3943bc4d;
    11'b00100010011: data <= 32'h3e00be7a;
    11'b00100010100: data <= 32'h3c25b8ac;
    11'b00100010101: data <= 32'hbc053afc;
    11'b00100010110: data <= 32'hc1253c0d;
    11'b00100010111: data <= 32'hbfdd2a47;
    11'b00100011000: data <= 32'hb547b868;
    11'b00100011001: data <= 32'h29d3b6cf;
    11'b00100011010: data <= 32'hbb02b5ae;
    11'b00100011011: data <= 32'hbc01b580;
    11'b00100011100: data <= 32'h37b33827;
    11'b00100011101: data <= 32'h3f0f4013;
    11'b00100011110: data <= 32'h3cab40f7;
    11'b00100011111: data <= 32'hb6733c47;
    11'b00100100000: data <= 32'hbb8eb874;
    11'b00100100001: data <= 32'hb20ab882;
    11'b00100100010: data <= 32'h3894356e;
    11'b00100100011: data <= 32'h3a9d2c5d;
    11'b00100100100: data <= 32'h3cf1bdd3;
    11'b00100100101: data <= 32'h3f22c016;
    11'b00100100110: data <= 32'h3d6eb8bb;
    11'b00100100111: data <= 32'hb3c63c83;
    11'b00100101000: data <= 32'hbdb93bf8;
    11'b00100101001: data <= 32'hbc2ab859;
    11'b00100101010: data <= 32'hb2c9bded;
    11'b00100101011: data <= 32'hb90dbcc1;
    11'b00100101100: data <= 32'hbeecb9bc;
    11'b00100101101: data <= 32'hbdbcb871;
    11'b00100101110: data <= 32'h378d2a31;
    11'b00100101111: data <= 32'h3ea53d0a;
    11'b00100110000: data <= 32'h38763f7c;
    11'b00100110001: data <= 32'hbd763cc5;
    11'b00100110010: data <= 32'hbee83610;
    11'b00100110011: data <= 32'hb768390b;
    11'b00100110100: data <= 32'h38ed3c70;
    11'b00100110101: data <= 32'h39f933ff;
    11'b00100110110: data <= 32'h3b0dbda5;
    11'b00100110111: data <= 32'h3e12be79;
    11'b00100111000: data <= 32'h3ed6328c;
    11'b00100111001: data <= 32'h3adb3f25;
    11'b00100111010: data <= 32'hac223c58;
    11'b00100111011: data <= 32'haef2bb4e;
    11'b00100111100: data <= 32'h1882bf50;
    11'b00100111101: data <= 32'hba34bcf3;
    11'b00100111110: data <= 32'hbe9eb9c9;
    11'b00100111111: data <= 32'hbbcebc1d;
    11'b00101000000: data <= 32'h3b2dbc4a;
    11'b00101000001: data <= 32'h3e36add9;
    11'b00101000010: data <= 32'hae243bd2;
    11'b00101000011: data <= 32'hc02b3c6c;
    11'b00101000100: data <= 32'hc0323a80;
    11'b00101000101: data <= 32'hb8de3bd7;
    11'b00101000110: data <= 32'h324d3c48;
    11'b00101000111: data <= 32'hb2e12e97;
    11'b00101001000: data <= 32'hb49bbc9e;
    11'b00101001001: data <= 32'h3a89ba8e;
    11'b00101001010: data <= 32'h3f7b3c8b;
    11'b00101001011: data <= 32'h3e8840af;
    11'b00101001100: data <= 32'h39973ced;
    11'b00101001101: data <= 32'h337eb9c3;
    11'b00101001110: data <= 32'h2d55bcd3;
    11'b00101001111: data <= 32'hb788b62b;
    11'b00101010000: data <= 32'hbb17b495;
    11'b00101010001: data <= 32'ha9dcbdd5;
    11'b00101010010: data <= 32'h3dd9c056;
    11'b00101010011: data <= 32'h3e53bcc2;
    11'b00101010100: data <= 32'hb3673614;
    11'b00101010101: data <= 32'hbfa73b7f;
    11'b00101010110: data <= 32'hbe9338d1;
    11'b00101010111: data <= 32'hb6e5369a;
    11'b00101011000: data <= 32'hb6aa3564;
    11'b00101011001: data <= 32'hbe08b4e2;
    11'b00101011010: data <= 32'hbe58bbde;
    11'b00101011011: data <= 32'h2fb9b57e;
    11'b00101011100: data <= 32'h3f273da9;
    11'b00101011101: data <= 32'h3eb9408f;
    11'b00101011110: data <= 32'h377f3d03;
    11'b00101011111: data <= 32'hb1f6acc3;
    11'b00101100000: data <= 32'hace22d53;
    11'b00101100001: data <= 32'hacb23b6f;
    11'b00101100010: data <= 32'hb03435c9;
    11'b00101100011: data <= 32'h3891be64;
    11'b00101100100: data <= 32'h3ebdc135;
    11'b00101100101: data <= 32'h3ec4bd8c;
    11'b00101100110: data <= 32'h349d374a;
    11'b00101100111: data <= 32'hbab63af1;
    11'b00101101000: data <= 32'hb814293e;
    11'b00101101001: data <= 32'h2a3db809;
    11'b00101101010: data <= 32'hbaa2b72d;
    11'b00101101011: data <= 32'hc0b9b90f;
    11'b00101101100: data <= 32'hc074bc22;
    11'b00101101101: data <= 32'haf1ab8d5;
    11'b00101101110: data <= 32'h3e6539a7;
    11'b00101101111: data <= 32'h3c703de8;
    11'b00101110000: data <= 32'hb7203c13;
    11'b00101110001: data <= 32'hbbbe38ad;
    11'b00101110010: data <= 32'hb5593d12;
    11'b00101110011: data <= 32'h2d5b3fb6;
    11'b00101110100: data <= 32'ha8e33a77;
    11'b00101110101: data <= 32'h3495bdba;
    11'b00101110110: data <= 32'h3d03c06f;
    11'b00101110111: data <= 32'h3ed2b960;
    11'b00101111000: data <= 32'h3c6f3c55;
    11'b00101111001: data <= 32'h38183b97;
    11'b00101111010: data <= 32'h3957b66b;
    11'b00101111011: data <= 32'h388abbe8;
    11'b00101111100: data <= 32'hba8cb888;
    11'b00101111101: data <= 32'hc0a5b80c;
    11'b00101111110: data <= 32'hbf89bccc;
    11'b00101111111: data <= 32'h33f3bdcf;
    11'b00110000000: data <= 32'h3deab8fc;
    11'b00110000001: data <= 32'h36a53545;
    11'b00110000010: data <= 32'hbd0f38c1;
    11'b00110000011: data <= 32'hbd9e3aa3;
    11'b00110000100: data <= 32'hb6183e9e;
    11'b00110000101: data <= 32'hac634013;
    11'b00110000110: data <= 32'hb9f03a26;
    11'b00110000111: data <= 32'hbad2bc9b;
    11'b00110001000: data <= 32'h34d3bd9b;
    11'b00110001001: data <= 32'h3e07353c;
    11'b00110001010: data <= 32'h3eac3ecc;
    11'b00110001011: data <= 32'h3d3d3c1b;
    11'b00110001100: data <= 32'h3cc9b6e8;
    11'b00110001101: data <= 32'h3a70b8d1;
    11'b00110001110: data <= 32'hb77a33e8;
    11'b00110001111: data <= 32'hbe3a315c;
    11'b00110010000: data <= 32'hbb5bbd0f;
    11'b00110010001: data <= 32'h3ae8c09f;
    11'b00110010010: data <= 32'h3dddbf04;
    11'b00110010011: data <= 32'h2e3fb7d0;
    11'b00110010100: data <= 32'hbd3b32f7;
    11'b00110010101: data <= 32'hbbfd385c;
    11'b00110010110: data <= 32'h215b3c6a;
    11'b00110010111: data <= 32'hb5383d3b;
    11'b00110011000: data <= 32'hbf283546;
    11'b00110011001: data <= 32'hc05cbba9;
    11'b00110011010: data <= 32'hb922ba40;
    11'b00110011011: data <= 32'h3cac3a62;
    11'b00110011100: data <= 32'h3e6f3eca;
    11'b00110011101: data <= 32'h3c6f3ae8;
    11'b00110011110: data <= 32'h3a94afd4;
    11'b00110011111: data <= 32'h3929370a;
    11'b00110100000: data <= 32'hab403e59;
    11'b00110100001: data <= 32'hb98c3c52;
    11'b00110100010: data <= 32'hb047bc6e;
    11'b00110100011: data <= 32'h3ca1c137;
    11'b00110100100: data <= 32'h3db4bff5;
    11'b00110100101: data <= 32'h34eab808;
    11'b00110100110: data <= 32'hb7a62ecd;
    11'b00110100111: data <= 32'h30e9a830;
    11'b00110101000: data <= 32'h3a1d2efc;
    11'b00110101001: data <= 32'hb69e3616;
    11'b00110101010: data <= 32'hc0f5acfb;
    11'b00110101011: data <= 32'hc1bdbb26;
    11'b00110101100: data <= 32'hbc0aba1a;
    11'b00110101101: data <= 32'h3b1b3546;
    11'b00110101110: data <= 32'h3c073b19;
    11'b00110101111: data <= 32'h309a35b8;
    11'b00110110000: data <= 32'hac793232;
    11'b00110110001: data <= 32'h34ea3dc6;
    11'b00110110010: data <= 32'h31c44149;
    11'b00110110011: data <= 32'hb5b03ed6;
    11'b00110110100: data <= 32'hb1deba66;
    11'b00110110101: data <= 32'h39e8c058;
    11'b00110110110: data <= 32'h3cbabcfb;
    11'b00110110111: data <= 32'h3a38324a;
    11'b00110111000: data <= 32'h396c3417;
    11'b00110111001: data <= 32'h3d97b83c;
    11'b00110111010: data <= 32'h3e05b8ac;
    11'b00110111011: data <= 32'hb2c4289d;
    11'b00110111100: data <= 32'hc0bd22df;
    11'b00110111101: data <= 32'hc109baa1;
    11'b00110111110: data <= 32'hb8f6bd0f;
    11'b00110111111: data <= 32'h3a80ba5a;
    11'b00111000000: data <= 32'h345cb546;
    11'b00111000001: data <= 32'hbad4b52a;
    11'b00111000010: data <= 32'hb9c3327a;
    11'b00111000011: data <= 32'h32853ef5;
    11'b00111000100: data <= 32'h3337418a;
    11'b00111000101: data <= 32'hb9d23ebe;
    11'b00111000110: data <= 32'hbc6eb840;
    11'b00111000111: data <= 32'hb46fbd48;
    11'b00111001000: data <= 32'h39a6ae2f;
    11'b00111001001: data <= 32'h3c3f3c0b;
    11'b00111001010: data <= 32'h3d783683;
    11'b00111001011: data <= 32'h3fe0b9c8;
    11'b00111001100: data <= 32'h3f40b813;
    11'b00111001101: data <= 32'h315b3905;
    11'b00111001110: data <= 32'hbe4539e5;
    11'b00111001111: data <= 32'hbdb9b8e0;
    11'b00111010000: data <= 32'h3181bf48;
    11'b00111010001: data <= 32'h3b10bf32;
    11'b00111010010: data <= 32'hb1aabcda;
    11'b00111010011: data <= 32'hbcbeba9b;
    11'b00111010100: data <= 32'hb856b10a;
    11'b00111010101: data <= 32'h38ff3c97;
    11'b00111010110: data <= 32'h33de3fca;
    11'b00111010111: data <= 32'hbdd23c65;
    11'b00111011000: data <= 32'hc096b6be;
    11'b00111011001: data <= 32'hbd37b8c0;
    11'b00111011010: data <= 32'h320a3923;
    11'b00111011011: data <= 32'h3b063cf7;
    11'b00111011100: data <= 32'h3c7733a0;
    11'b00111011101: data <= 32'h3e24b966;
    11'b00111011110: data <= 32'h3e2e32a3;
    11'b00111011111: data <= 32'h38093f41;
    11'b00111100000: data <= 32'hb8f13efa;
    11'b00111100001: data <= 32'hb660b364;
    11'b00111100010: data <= 32'h399fbfc9;
    11'b00111100011: data <= 32'h3ae9bfe5;
    11'b00111100100: data <= 32'hb29cbcd3;
    11'b00111100101: data <= 32'hb973bb09;
    11'b00111100110: data <= 32'h3719b979;
    11'b00111100111: data <= 32'h3de62d3a;
    11'b00111101000: data <= 32'h36913a60;
    11'b00111101001: data <= 32'hbfbd3747;
    11'b00111101010: data <= 32'hc1d2b679;
    11'b00111101011: data <= 32'hbebeb5cd;
    11'b00111101100: data <= 32'hadc737f1;
    11'b00111101101: data <= 32'h34b038e5;
    11'b00111101110: data <= 32'h2dadb5bc;
    11'b00111101111: data <= 32'h3731b90a;
    11'b00111110000: data <= 32'h3bd73bc3;
    11'b00111110001: data <= 32'h39644194;
    11'b00111110010: data <= 32'hae0a40d6;
    11'b00111110011: data <= 32'hb02e3045;
    11'b00111110100: data <= 32'h37bdbdf2;
    11'b00111110101: data <= 32'h385cbcae;
    11'b00111110110: data <= 32'ha3f8b582;
    11'b00111110111: data <= 32'h32bbb835;
    11'b00111111000: data <= 32'h3e68bc6a;
    11'b00111111001: data <= 32'h4096ba2c;
    11'b00111111010: data <= 32'h39cb3097;
    11'b00111111011: data <= 32'hbf0a3536;
    11'b00111111100: data <= 32'hc101b4a5;
    11'b00111111101: data <= 32'hbcaeb8b4;
    11'b00111111110: data <= 32'h1cbfb580;
    11'b00111111111: data <= 32'hb5deb811;
    11'b01000000000: data <= 32'hbc30bc90;
    11'b01000000001: data <= 32'hb7f9ba44;
    11'b01000000010: data <= 32'h391d3ca6;
    11'b01000000011: data <= 32'h39e741ba;
    11'b01000000100: data <= 32'hb279409f;
    11'b01000000101: data <= 32'hba0d3466;
    11'b01000000110: data <= 32'hb6b7b991;
    11'b01000000111: data <= 32'ha9f32e82;
    11'b01000001000: data <= 32'h2c1b3a03;
    11'b01000001001: data <= 32'h3a16b014;
    11'b01000001010: data <= 32'h403fbd25;
    11'b01000001011: data <= 32'h411fbb8b;
    11'b01000001100: data <= 32'h3c1c36d0;
    11'b01000001101: data <= 32'hbbfc3b53;
    11'b01000001110: data <= 32'hbd3829c3;
    11'b01000001111: data <= 32'haf70bb43;
    11'b01000010000: data <= 32'h352abcb4;
    11'b01000010001: data <= 32'hba45bd64;
    11'b01000010010: data <= 32'hbe6ebe9b;
    11'b01000010011: data <= 32'hb918bc7e;
    11'b01000010100: data <= 32'h3b3538ac;
    11'b01000010101: data <= 32'h3ae63fc6;
    11'b01000010110: data <= 32'hb9663df5;
    11'b01000010111: data <= 32'hbef730ab;
    11'b01000011000: data <= 32'hbd9ca438;
    11'b01000011001: data <= 32'hb8eb3c36;
    11'b01000011010: data <= 32'hb1123d38;
    11'b01000011011: data <= 32'h37e4af18;
    11'b01000011100: data <= 32'h3e70bd4b;
    11'b01000011101: data <= 32'h4030b7d2;
    11'b01000011110: data <= 32'h3c953d8b;
    11'b01000011111: data <= 32'hae843f7d;
    11'b01000100000: data <= 32'hacc03811;
    11'b01000100001: data <= 32'h39efbb84;
    11'b01000100010: data <= 32'h381dbd37;
    11'b01000100011: data <= 32'hbafebd1a;
    11'b01000100100: data <= 32'hbd77be36;
    11'b01000100101: data <= 32'h2e88bddd;
    11'b01000100110: data <= 32'h3ec1b6dd;
    11'b01000100111: data <= 32'h3c8938e0;
    11'b01000101000: data <= 32'hbc0e3824;
    11'b01000101001: data <= 32'hc08fac86;
    11'b01000101010: data <= 32'hbef03405;
    11'b01000101011: data <= 32'hba583cad;
    11'b01000101100: data <= 32'hb8d73b8f;
    11'b01000101101: data <= 32'hb7dbb902;
    11'b01000101110: data <= 32'h35b4bd95;
    11'b01000101111: data <= 32'h3cd92e49;
    11'b01000110000: data <= 32'h3c444084;
    11'b01000110001: data <= 32'h36f34105;
    11'b01000110010: data <= 32'h373f3a97;
    11'b01000110011: data <= 32'h3a86b887;
    11'b01000110100: data <= 32'h34d8b839;
    11'b01000110101: data <= 32'hba6ab444;
    11'b01000110110: data <= 32'hb96dbb3a;
    11'b01000110111: data <= 32'h3c85be88;
    11'b01000111000: data <= 32'h40f7bd1a;
    11'b01000111001: data <= 32'h3dcab4c6;
    11'b01000111010: data <= 32'hbafd2ca9;
    11'b01000111011: data <= 32'hbf85ae1b;
    11'b01000111100: data <= 32'hbc5f3057;
    11'b01000111101: data <= 32'hb6f8386f;
    11'b01000111110: data <= 32'hbc19a587;
    11'b01000111111: data <= 32'hbe6fbd8f;
    11'b01001000000: data <= 32'hbab3be5d;
    11'b01001000001: data <= 32'h384b3464;
    11'b01001000010: data <= 32'h3ba840a4;
    11'b01001000011: data <= 32'h36b9409a;
    11'b01001000100: data <= 32'h2c7839f5;
    11'b01001000101: data <= 32'h2e1620b8;
    11'b01001000110: data <= 32'hb44739c7;
    11'b01001000111: data <= 32'hba633c43;
    11'b01001001000: data <= 32'hb20eb116;
    11'b01001001001: data <= 32'h3e81be74;
    11'b01001001010: data <= 32'h415abe15;
    11'b01001001011: data <= 32'h3e4fb456;
    11'b01001001100: data <= 32'hb4b23725;
    11'b01001001101: data <= 32'hb99e3284;
    11'b01001001110: data <= 32'h31eead5f;
    11'b01001001111: data <= 32'h3358b1a1;
    11'b01001010000: data <= 32'hbcdeba8a;
    11'b01001010001: data <= 32'hc072bf6b;
    11'b01001010010: data <= 32'hbcf6bf40;
    11'b01001010011: data <= 32'h3864b11f;
    11'b01001010100: data <= 32'h3c143daa;
    11'b01001010101: data <= 32'h2b7b3d16;
    11'b01001010110: data <= 32'hba363472;
    11'b01001010111: data <= 32'hba963740;
    11'b01001011000: data <= 32'hba833edb;
    11'b01001011001: data <= 32'hbba63f91;
    11'b01001011010: data <= 32'hb5b2307d;
    11'b01001011011: data <= 32'h3c7ebe3a;
    11'b01001011100: data <= 32'h400ebcb5;
    11'b01001011101: data <= 32'h3d85382a;
    11'b01001011110: data <= 32'h35de3d42;
    11'b01001011111: data <= 32'h387a3948;
    11'b01001100000: data <= 32'h3d4ab02b;
    11'b01001100001: data <= 32'h39dfb5c1;
    11'b01001100010: data <= 32'hbcbaba08;
    11'b01001100011: data <= 32'hc02cbe6c;
    11'b01001100100: data <= 32'hb991bf7d;
    11'b01001100101: data <= 32'h3ce0bb94;
    11'b01001100110: data <= 32'h3d272b6e;
    11'b01001100111: data <= 32'hb41624b1;
    11'b01001101000: data <= 32'hbd52b470;
    11'b01001101001: data <= 32'hbca33884;
    11'b01001101010: data <= 32'hbb083fb6;
    11'b01001101011: data <= 32'hbca93f00;
    11'b01001101100: data <= 32'hbc88b331;
    11'b01001101101: data <= 32'hb0b0be79;
    11'b01001101110: data <= 32'h3af0b928;
    11'b01001101111: data <= 32'h3b8e3d78;
    11'b01001110000: data <= 32'h39c23fcc;
    11'b01001110001: data <= 32'h3cb63b2f;
    11'b01001110010: data <= 32'h3e902b5d;
    11'b01001110011: data <= 32'h39af339a;
    11'b01001110100: data <= 32'hbc553443;
    11'b01001110101: data <= 32'hbde5b98e;
    11'b01001110110: data <= 32'h3460beb8;
    11'b01001110111: data <= 32'h3ffebe5c;
    11'b01001111000: data <= 32'h3e38bb79;
    11'b01001111001: data <= 32'hb3f7b994;
    11'b01001111010: data <= 32'hbc4db843;
    11'b01001111011: data <= 32'hb8193665;
    11'b01001111100: data <= 32'hb48d3d9c;
    11'b01001111101: data <= 32'hbcf33b03;
    11'b01001111110: data <= 32'hc013bbac;
    11'b01001111111: data <= 32'hbdacbf2b;
    11'b01010000000: data <= 32'hae70b61b;
    11'b01010000001: data <= 32'h387d3e2d;
    11'b01010000010: data <= 32'h39043ef6;
    11'b01010000011: data <= 32'h3b2838e9;
    11'b01010000100: data <= 32'h3c3234f9;
    11'b01010000101: data <= 32'h322a3d1b;
    11'b01010000110: data <= 32'hbc4c3ead;
    11'b01010000111: data <= 32'hbb8535ae;
    11'b01010001000: data <= 32'h3ad1bd65;
    11'b01010001001: data <= 32'h4066bee7;
    11'b01010001010: data <= 32'h3e11bc0c;
    11'b01010001011: data <= 32'h2999b7d8;
    11'b01010001100: data <= 32'hae52b51b;
    11'b01010001101: data <= 32'h3aa631c0;
    11'b01010001110: data <= 32'h39853951;
    11'b01010001111: data <= 32'hbc5f2709;
    11'b01010010000: data <= 32'hc108bdc2;
    11'b01010010001: data <= 32'hbfb7bf8a;
    11'b01010010010: data <= 32'hb4b3b88d;
    11'b01010010011: data <= 32'h37f53a9d;
    11'b01010010100: data <= 32'h3420393b;
    11'b01010010101: data <= 32'h2c8cb107;
    11'b01010010110: data <= 32'h2f0b3679;
    11'b01010010111: data <= 32'hb5f64039;
    11'b01010011000: data <= 32'hbc934136;
    11'b01010011001: data <= 32'hbb393b2b;
    11'b01010011010: data <= 32'h382cbc7a;
    11'b01010011011: data <= 32'h3e07bd6e;
    11'b01010011100: data <= 32'h3c1fb447;
    11'b01010011101: data <= 32'h35a335cc;
    11'b01010011110: data <= 32'h3bf630cc;
    11'b01010011111: data <= 32'h402a2d17;
    11'b01010100000: data <= 32'h3de13526;
    11'b01010100001: data <= 32'hbab8ac20;
    11'b01010100010: data <= 32'hc0aabca9;
    11'b01010100011: data <= 32'hbdcdbebc;
    11'b01010100100: data <= 32'h3526bc0e;
    11'b01010100101: data <= 32'h3a15b5b7;
    11'b01010100110: data <= 32'had80b9bd;
    11'b01010100111: data <= 32'hb8cbbc10;
    11'b01010101000: data <= 32'hb5c8341b;
    11'b01010101001: data <= 32'hb6ed4084;
    11'b01010101010: data <= 32'hbc844119;
    11'b01010101011: data <= 32'hbd703904;
    11'b01010101100: data <= 32'hb892bc98;
    11'b01010101101: data <= 32'h336eba75;
    11'b01010101110: data <= 32'h345a3947;
    11'b01010101111: data <= 32'h36943c71;
    11'b01010110000: data <= 32'h3e1b3669;
    11'b01010110001: data <= 32'h41022d82;
    11'b01010110010: data <= 32'h3e5a3906;
    11'b01010110011: data <= 32'hb9633a3c;
    11'b01010110100: data <= 32'hbed1b0cb;
    11'b01010110101: data <= 32'hb6eebca5;
    11'b01010110110: data <= 32'h3cc2bd59;
    11'b01010110111: data <= 32'h3c34bcfb;
    11'b01010111000: data <= 32'hb30cbe39;
    11'b01010111001: data <= 32'hb8cfbdd9;
    11'b01010111010: data <= 32'h2f2ca47c;
    11'b01010111011: data <= 32'h33ee3eda;
    11'b01010111100: data <= 32'hbb0b3ea0;
    11'b01010111101: data <= 32'hbfb8b15c;
    11'b01010111110: data <= 32'hbee6bd67;
    11'b01010111111: data <= 32'hbafeb703;
    11'b01011000000: data <= 32'hb5973c3b;
    11'b01011000001: data <= 32'h31383c47;
    11'b01011000010: data <= 32'h3cdc2abf;
    11'b01011000011: data <= 32'h3fb32902;
    11'b01011000100: data <= 32'h3c2e3d54;
    11'b01011000101: data <= 32'hb981401b;
    11'b01011000110: data <= 32'hbc5f3c31;
    11'b01011000111: data <= 32'h355eb868;
    11'b01011001000: data <= 32'h3e37bd15;
    11'b01011001001: data <= 32'h3bccbd23;
    11'b01011001010: data <= 32'hb257bd92;
    11'b01011001011: data <= 32'h2a6fbd11;
    11'b01011001100: data <= 32'h3d47b35f;
    11'b01011001101: data <= 32'h3d7e3b59;
    11'b01011001110: data <= 32'hb6d23931;
    11'b01011001111: data <= 32'hc055ba6f;
    11'b01011010000: data <= 32'hc05ebdb8;
    11'b01011010001: data <= 32'hbc94b638;
    11'b01011010010: data <= 32'hb7c23934;
    11'b01011010011: data <= 32'hb3433003;
    11'b01011010100: data <= 32'h3599baeb;
    11'b01011010101: data <= 32'h3ae0b22e;
    11'b01011010110: data <= 32'h355a3f96;
    11'b01011010111: data <= 32'hba2341db;
    11'b01011011000: data <= 32'hbad63ec9;
    11'b01011011001: data <= 32'h34c1b238;
    11'b01011011010: data <= 32'h3c0bbac1;
    11'b01011011011: data <= 32'h35adb80a;
    11'b01011011100: data <= 32'hb30ab72f;
    11'b01011011101: data <= 32'h3ad5b964;
    11'b01011011110: data <= 32'h4101b4e1;
    11'b01011011111: data <= 32'h40933690;
    11'b01011100000: data <= 32'h1fb3348c;
    11'b01011100001: data <= 32'hbf89b986;
    11'b01011100010: data <= 32'hbeb0bc78;
    11'b01011100011: data <= 32'hb797b815;
    11'b01011100100: data <= 32'hb026b36e;
    11'b01011100101: data <= 32'hb853bcaf;
    11'b01011100110: data <= 32'hb743bf87;
    11'b01011100111: data <= 32'h3067b88e;
    11'b01011101000: data <= 32'h2ea23f9b;
    11'b01011101001: data <= 32'hb95d41ad;
    11'b01011101010: data <= 32'hbc043da6;
    11'b01011101011: data <= 32'hb7d1b465;
    11'b01011101100: data <= 32'hb1c4b50b;
    11'b01011101101: data <= 32'hb8a0383f;
    11'b01011101110: data <= 32'hb6e43832;
    11'b01011101111: data <= 32'h3cd6b3e3;
    11'b01011110000: data <= 32'h41c8b593;
    11'b01011110001: data <= 32'h40dd36f9;
    11'b01011110010: data <= 32'h31803a90;
    11'b01011110011: data <= 32'hbd07334f;
    11'b01011110100: data <= 32'hb883b6a7;
    11'b01011110101: data <= 32'h38bcb843;
    11'b01011110110: data <= 32'h3561bb4f;
    11'b01011110111: data <= 32'hb993bfec;
    11'b01011111000: data <= 32'hb9a6c0cb;
    11'b01011111001: data <= 32'h34eabb2a;
    11'b01011111010: data <= 32'h395c3d55;
    11'b01011111011: data <= 32'hb4053f79;
    11'b01011111100: data <= 32'hbd06372e;
    11'b01011111101: data <= 32'hbda2b91f;
    11'b01011111110: data <= 32'hbd092b17;
    11'b01011111111: data <= 32'hbd3e3c9a;
    11'b01100000000: data <= 32'hba4d3a3f;
    11'b01100000001: data <= 32'h3ac2b761;
    11'b01100000010: data <= 32'h407fb85d;
    11'b01100000011: data <= 32'h3f053a8b;
    11'b01100000100: data <= 32'h22e83f5d;
    11'b01100000101: data <= 32'hb93c3d96;
    11'b01100000110: data <= 32'h366a357c;
    11'b01100000111: data <= 32'h3cfab4d6;
    11'b01100001000: data <= 32'h3694baf0;
    11'b01100001001: data <= 32'hba64bf15;
    11'b01100001010: data <= 32'hb5eac039;
    11'b01100001011: data <= 32'h3cfdbbf7;
    11'b01100001100: data <= 32'h3f093869;
    11'b01100001101: data <= 32'h3604397d;
    11'b01100001110: data <= 32'hbd1fb777;
    11'b01100001111: data <= 32'hbf01bb1b;
    11'b01100010000: data <= 32'hbdfe326c;
    11'b01100010001: data <= 32'hbda13c2e;
    11'b01100010010: data <= 32'hbc6e2f43;
    11'b01100010011: data <= 32'ha31bbd51;
    11'b01100010100: data <= 32'h3c1fbbb6;
    11'b01100010101: data <= 32'h3a403c86;
    11'b01100010110: data <= 32'hb3e64123;
    11'b01100010111: data <= 32'hb591400e;
    11'b01100011000: data <= 32'h393339b5;
    11'b01100011001: data <= 32'h3be82ede;
    11'b01100011010: data <= 32'hb090ad20;
    11'b01100011011: data <= 32'hbc08b992;
    11'b01100011100: data <= 32'h310ebd1d;
    11'b01100011101: data <= 32'h4085bb15;
    11'b01100011110: data <= 32'h4155916d;
    11'b01100011111: data <= 32'h3afe2a65;
    11'b01100100000: data <= 32'hbbaab933;
    11'b01100100001: data <= 32'hbcd8b951;
    11'b01100100010: data <= 32'hb9c33423;
    11'b01100100011: data <= 32'hbac83746;
    11'b01100100100: data <= 32'hbcfcbbf3;
    11'b01100100101: data <= 32'hbabdc0b2;
    11'b01100100110: data <= 32'h2b0dbdcc;
    11'b01100100111: data <= 32'h33ce3c2d;
    11'b01100101000: data <= 32'hb44840db;
    11'b01100101001: data <= 32'hb5603ea2;
    11'b01100101010: data <= 32'h3150378c;
    11'b01100101011: data <= 32'h1df137c1;
    11'b01100101100: data <= 32'hbc513bc4;
    11'b01100101101: data <= 32'hbd753819;
    11'b01100101110: data <= 32'h35f8b855;
    11'b01100101111: data <= 32'h4128ba45;
    11'b01100110000: data <= 32'h4180af37;
    11'b01100110001: data <= 32'h3b6a347c;
    11'b01100110010: data <= 32'hb72b28f6;
    11'b01100110011: data <= 32'hada72849;
    11'b01100110100: data <= 32'h387e3689;
    11'b01100110101: data <= 32'hace9a9c1;
    11'b01100110110: data <= 32'hbcf1bedb;
    11'b01100110111: data <= 32'hbcd3c1a9;
    11'b01100111000: data <= 32'had0fbedf;
    11'b01100111001: data <= 32'h38753867;
    11'b01100111010: data <= 32'h30353dc1;
    11'b01100111011: data <= 32'hb66b3800;
    11'b01100111100: data <= 32'hb84db1e7;
    11'b01100111101: data <= 32'hbbbd396b;
    11'b01100111110: data <= 32'hbf393eb8;
    11'b01100111111: data <= 32'hbee13c45;
    11'b01101000000: data <= 32'h28c8b7b0;
    11'b01101000001: data <= 32'h3fa3bb7a;
    11'b01101000010: data <= 32'h3f9e2d33;
    11'b01101000011: data <= 32'h38043c3a;
    11'b01101000100: data <= 32'ha5fa3c53;
    11'b01101000101: data <= 32'h3b983a74;
    11'b01101000110: data <= 32'h3e073989;
    11'b01101000111: data <= 32'h34b4251f;
    11'b01101001000: data <= 32'hbd0cbde2;
    11'b01101001001: data <= 32'hbc31c0d0;
    11'b01101001010: data <= 32'h38c5be58;
    11'b01101001011: data <= 32'h3dfeac21;
    11'b01101001100: data <= 32'h3a45323d;
    11'b01101001101: data <= 32'hb532b99e;
    11'b01101001110: data <= 32'hba83b9f5;
    11'b01101001111: data <= 32'hbca939be;
    11'b01101010000: data <= 32'hbf343ef4;
    11'b01101010001: data <= 32'hbf6c396f;
    11'b01101010010: data <= 32'hb967bcb4;
    11'b01101010011: data <= 32'h3919bd82;
    11'b01101010100: data <= 32'h3939342a;
    11'b01101010101: data <= 32'had2f3eb5;
    11'b01101010110: data <= 32'h30e43ea7;
    11'b01101010111: data <= 32'h3d653c74;
    11'b01101011000: data <= 32'h3e2c3bc6;
    11'b01101011001: data <= 32'hab9c3988;
    11'b01101011010: data <= 32'hbdf0b596;
    11'b01101011011: data <= 32'hb96cbd41;
    11'b01101011100: data <= 32'h3ddcbc9c;
    11'b01101011101: data <= 32'h40b1b776;
    11'b01101011110: data <= 32'h3d04b89f;
    11'b01101011111: data <= 32'hacc2bcc3;
    11'b01101100000: data <= 32'hb5a3ba04;
    11'b01101100001: data <= 32'hb5863a2a;
    11'b01101100010: data <= 32'hbc073d45;
    11'b01101100011: data <= 32'hbebcb40b;
    11'b01101100100: data <= 32'hbd5ec03f;
    11'b01101100101: data <= 32'hb765bf74;
    11'b01101100110: data <= 32'hb26d3214;
    11'b01101100111: data <= 32'hb5da3e4c;
    11'b01101101000: data <= 32'h304e3d04;
    11'b01101101001: data <= 32'h3c293963;
    11'b01101101010: data <= 32'h3a1b3c44;
    11'b01101101011: data <= 32'hbb463e53;
    11'b01101101100: data <= 32'hbf733bc4;
    11'b01101101101: data <= 32'hb7e9b411;
    11'b01101101110: data <= 32'h3f23ba0b;
    11'b01101101111: data <= 32'h40cab826;
    11'b01101110000: data <= 32'h3c97b830;
    11'b01101110001: data <= 32'h3232b9dd;
    11'b01101110010: data <= 32'h38f8b138;
    11'b01101110011: data <= 32'h3c273ba3;
    11'b01101110100: data <= 32'h2d5e3b20;
    11'b01101110101: data <= 32'hbd6bbb86;
    11'b01101110110: data <= 32'hbe78c126;
    11'b01101110111: data <= 32'hba28c007;
    11'b01101111000: data <= 32'hb0bbaef4;
    11'b01101111001: data <= 32'haee239b7;
    11'b01101111010: data <= 32'h2ea31bd8;
    11'b01101111011: data <= 32'h3716b4ae;
    11'b01101111100: data <= 32'hb0a23b74;
    11'b01101111101: data <= 32'hbe70405b;
    11'b01101111110: data <= 32'hc04a3ec7;
    11'b01101111111: data <= 32'hb97b2e08;
    11'b01110000000: data <= 32'h3ce3b9d2;
    11'b01110000001: data <= 32'h3ddcb58e;
    11'b01110000010: data <= 32'h36e82fbe;
    11'b01110000011: data <= 32'h34b032c5;
    11'b01110000100: data <= 32'h3e2238a9;
    11'b01110000101: data <= 32'h404b3cd2;
    11'b01110000110: data <= 32'h3a1f3ae6;
    11'b01110000111: data <= 32'hbca6ba3e;
    11'b01110001000: data <= 32'hbdd8c02a;
    11'b01110001001: data <= 32'hb3c9be7c;
    11'b01110001010: data <= 32'h3947b69d;
    11'b01110001011: data <= 32'h380eb666;
    11'b01110001100: data <= 32'h31bebd6f;
    11'b01110001101: data <= 32'h2fe0bcbb;
    11'b01110001110: data <= 32'hb66a39be;
    11'b01110001111: data <= 32'hbe36406e;
    11'b01110010000: data <= 32'hc01d3dde;
    11'b01110010001: data <= 32'hbc73b6ed;
    11'b01110010010: data <= 32'h2cf7bc72;
    11'b01110010011: data <= 32'h2b77b206;
    11'b01110010100: data <= 32'hb7e939ea;
    11'b01110010101: data <= 32'h31e53a98;
    11'b01110010110: data <= 32'h3f8e3adb;
    11'b01110010111: data <= 32'h40b53d3b;
    11'b01110011000: data <= 32'h38ee3d23;
    11'b01110011001: data <= 32'hbd313302;
    11'b01110011010: data <= 32'hbc79babf;
    11'b01110011011: data <= 32'h38b0bab9;
    11'b01110011100: data <= 32'h3e0cb810;
    11'b01110011101: data <= 32'h3babbc71;
    11'b01110011110: data <= 32'h34d4c00e;
    11'b01110011111: data <= 32'h360fbdba;
    11'b01110100000: data <= 32'h34e43931;
    11'b01110100001: data <= 32'hb90a3f48;
    11'b01110100010: data <= 32'hbe3038d5;
    11'b01110100011: data <= 32'hbdd8bd6b;
    11'b01110100100: data <= 32'hbb8fbe59;
    11'b01110100101: data <= 32'hbbe6b195;
    11'b01110100110: data <= 32'hbc3d3a5e;
    11'b01110100111: data <= 32'h1d853824;
    11'b01110101000: data <= 32'h3e6534ef;
    11'b01110101001: data <= 32'h3eae3c5c;
    11'b01110101010: data <= 32'hb1ad3f6d;
    11'b01110101011: data <= 32'hbea93dce;
    11'b01110101100: data <= 32'hbb1936a4;
    11'b01110101101: data <= 32'h3c17b011;
    11'b01110101110: data <= 32'h3e97b5bd;
    11'b01110101111: data <= 32'h3a25bc41;
    11'b01110110000: data <= 32'h34adbec6;
    11'b01110110001: data <= 32'h3c33bb7c;
    11'b01110110010: data <= 32'h3e613a80;
    11'b01110110011: data <= 32'h39483d7f;
    11'b01110110100: data <= 32'hbb02b12d;
    11'b01110110101: data <= 32'hbdfcbf86;
    11'b01110110110: data <= 32'hbcfbbeb8;
    11'b01110110111: data <= 32'hbc55b395;
    11'b01110111000: data <= 32'hbb8132d5;
    11'b01110111001: data <= 32'hac2fb91b;
    11'b01110111010: data <= 32'h3c02bacd;
    11'b01110111011: data <= 32'h39c238c9;
    11'b01110111100: data <= 32'hbb82405e;
    11'b01110111101: data <= 32'hbfa6404e;
    11'b01110111110: data <= 32'hbb163b80;
    11'b01110111111: data <= 32'h39a82d77;
    11'b01111000000: data <= 32'h3a81af71;
    11'b01111000001: data <= 32'hb012b6e3;
    11'b01111000010: data <= 32'h2870b9f1;
    11'b01111000011: data <= 32'h3eb4b0b9;
    11'b01111000100: data <= 32'h41583c32;
    11'b01111000101: data <= 32'h3e263cc9;
    11'b01111000110: data <= 32'hb735b2fa;
    11'b01111000111: data <= 32'hbcecbdf0;
    11'b01111001000: data <= 32'hb9dfbc81;
    11'b01111001001: data <= 32'hb4e6b249;
    11'b01111001010: data <= 32'hb4efb8dc;
    11'b01111001011: data <= 32'h2067bfd9;
    11'b01111001100: data <= 32'h3898bfd0;
    11'b01111001101: data <= 32'h34772ee2;
    11'b01111001110: data <= 32'hbbd94025;
    11'b01111001111: data <= 32'hbec53fc1;
    11'b01111010000: data <= 32'hbbed379f;
    11'b01111010001: data <= 32'hb0a9b46d;
    11'b01111010010: data <= 32'hb86629c8;
    11'b01111010011: data <= 32'hbd1e342c;
    11'b01111010100: data <= 32'hb632257c;
    11'b01111010101: data <= 32'h3f63334a;
    11'b01111010110: data <= 32'h41c73c37;
    11'b01111010111: data <= 32'h3df53d50;
    11'b01111011000: data <= 32'hb82937f7;
    11'b01111011001: data <= 32'hbafab4bb;
    11'b01111011010: data <= 32'h308eaf4a;
    11'b01111011011: data <= 32'h394e2a51;
    11'b01111011100: data <= 32'h33b5bc6a;
    11'b01111011101: data <= 32'h2c34c148;
    11'b01111011110: data <= 32'h38a2c0ae;
    11'b01111011111: data <= 32'h39baacde;
    11'b01111100000: data <= 32'haf943e8f;
    11'b01111100001: data <= 32'hbbac3c30;
    11'b01111100010: data <= 32'hbbddb83c;
    11'b01111100011: data <= 32'hbb73bab6;
    11'b01111100100: data <= 32'hbe6b2e32;
    11'b01111100101: data <= 32'hc00a3838;
    11'b01111100110: data <= 32'hb9dba85f;
    11'b01111100111: data <= 32'h3df6b3eb;
    11'b01111101000: data <= 32'h4060390a;
    11'b01111101001: data <= 32'h392d3e2d;
    11'b01111101010: data <= 32'hbba53de8;
    11'b01111101011: data <= 32'hb8f73bc4;
    11'b01111101100: data <= 32'h3a023a77;
    11'b01111101101: data <= 32'h3c1f36a9;
    11'b01111101110: data <= 32'h305fbbae;
    11'b01111101111: data <= 32'hafc9c09a;
    11'b01111110000: data <= 32'h3b40bf57;
    11'b01111110001: data <= 32'h3ef9301b;
    11'b01111110010: data <= 32'h3cb33cb9;
    11'b01111110011: data <= 32'haab5307b;
    11'b01111110100: data <= 32'hba06bd0f;
    11'b01111110101: data <= 32'hbc69bc1e;
    11'b01111110110: data <= 32'hbed731be;
    11'b01111110111: data <= 32'hbfbc3444;
    11'b01111111000: data <= 32'hba66bb68;
    11'b01111111001: data <= 32'h3b0abd9b;
    11'b01111111010: data <= 32'h3c80af12;
    11'b01111111011: data <= 32'hb4d43e46;
    11'b01111111100: data <= 32'hbd3d400a;
    11'b01111111101: data <= 32'hb80d3e0f;
    11'b01111111110: data <= 32'h39d73c6c;
    11'b01111111111: data <= 32'h375139a0;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    