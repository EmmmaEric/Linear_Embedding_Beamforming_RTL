
module memory_rom_39(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbd3a3b21;
    11'b00000000001: data <= 32'hb9b13870;
    11'b00000000010: data <= 32'h3a43b7e4;
    11'b00000000011: data <= 32'h3f6db3dd;
    11'b00000000100: data <= 32'h3c683d4f;
    11'b00000000101: data <= 32'hb899408f;
    11'b00000000110: data <= 32'hbb613e6c;
    11'b00000000111: data <= 32'h366835f8;
    11'b00000001000: data <= 32'h3d46b4dc;
    11'b00000001001: data <= 32'h385eba22;
    11'b00000001010: data <= 32'hb704bde6;
    11'b00000001011: data <= 32'h339cbe8a;
    11'b00000001100: data <= 32'h3f58b843;
    11'b00000001101: data <= 32'h401339e0;
    11'b00000001110: data <= 32'h35683810;
    11'b00000001111: data <= 32'hbd8cbaa6;
    11'b00000010000: data <= 32'hbed8bd04;
    11'b00000010001: data <= 32'hbd24b24b;
    11'b00000010010: data <= 32'hbc793805;
    11'b00000010011: data <= 32'hbafbb781;
    11'b00000010100: data <= 32'h2469be93;
    11'b00000010101: data <= 32'h3a0fbad9;
    11'b00000010110: data <= 32'h34543dc6;
    11'b00000010111: data <= 32'hba534178;
    11'b00000011000: data <= 32'hba5d3fb9;
    11'b00000011001: data <= 32'h3405383b;
    11'b00000011010: data <= 32'h38cb2a81;
    11'b00000011011: data <= 32'hb5ca2cca;
    11'b00000011100: data <= 32'hbac4b576;
    11'b00000011101: data <= 32'h3915ba2c;
    11'b00000011110: data <= 32'h4160b557;
    11'b00000011111: data <= 32'h4187371e;
    11'b00000100000: data <= 32'h39f2350f;
    11'b00000100001: data <= 32'hbbeab83a;
    11'b00000100010: data <= 32'hbbbbb97b;
    11'b00000100011: data <= 32'hb4a49f1d;
    11'b00000100100: data <= 32'hb64dada9;
    11'b00000100101: data <= 32'hbac5be56;
    11'b00000100110: data <= 32'hb84dc14a;
    11'b00000100111: data <= 32'h320dbd88;
    11'b00000101000: data <= 32'h30fd3cac;
    11'b00000101001: data <= 32'hb86a408f;
    11'b00000101010: data <= 32'hba2e3cf9;
    11'b00000101011: data <= 32'hb65b2b77;
    11'b00000101100: data <= 32'hb89b3435;
    11'b00000101101: data <= 32'hbdc63b5c;
    11'b00000101110: data <= 32'hbd6a3895;
    11'b00000101111: data <= 32'h38ceb53b;
    11'b00000110000: data <= 32'h4150b5bb;
    11'b00000110001: data <= 32'h4104376f;
    11'b00000110010: data <= 32'h38a23af2;
    11'b00000110011: data <= 32'hb8943812;
    11'b00000110100: data <= 32'h2d5e3474;
    11'b00000110101: data <= 32'h3ae83590;
    11'b00000110110: data <= 32'h33e9b5a0;
    11'b00000110111: data <= 32'hba8fc002;
    11'b00000111000: data <= 32'hb92bc1b3;
    11'b00000111001: data <= 32'h37d4be11;
    11'b00000111010: data <= 32'h3b49392d;
    11'b00000111011: data <= 32'h311c3ccb;
    11'b00000111100: data <= 32'hb93e2820;
    11'b00000111101: data <= 32'hbba0b8fe;
    11'b00000111110: data <= 32'hbd813551;
    11'b00000111111: data <= 32'hc00d3d3b;
    11'b00001000000: data <= 32'hbecb393d;
    11'b00001000001: data <= 32'h2eb8b9c0;
    11'b00001000010: data <= 32'h3ef9ba4d;
    11'b00001000011: data <= 32'h3dd23891;
    11'b00001000100: data <= 32'h24073e96;
    11'b00001000101: data <= 32'hb5113e34;
    11'b00001000110: data <= 32'h3a853c42;
    11'b00001000111: data <= 32'h3d8a39fb;
    11'b00001001000: data <= 32'h3377a4f3;
    11'b00001001001: data <= 32'hbc1abdab;
    11'b00001001010: data <= 32'hb6f0c045;
    11'b00001001011: data <= 32'h3d61bcd0;
    11'b00001001100: data <= 32'h400f3184;
    11'b00001001101: data <= 32'h3bbf315c;
    11'b00001001110: data <= 32'hb5f2baf7;
    11'b00001001111: data <= 32'hbb51bb6e;
    11'b00001010000: data <= 32'hbcd236b9;
    11'b00001010001: data <= 32'hbee53ca6;
    11'b00001010010: data <= 32'hbec0ace4;
    11'b00001010011: data <= 32'hb87fbef6;
    11'b00001010100: data <= 32'h3844bdea;
    11'b00001010101: data <= 32'h35513828;
    11'b00001010110: data <= 32'hb77d3fef;
    11'b00001010111: data <= 32'hb31b3f4b;
    11'b00001011000: data <= 32'h3b283c9a;
    11'b00001011001: data <= 32'h3bc03bda;
    11'b00001011010: data <= 32'hb83739f4;
    11'b00001011011: data <= 32'hbe12b1f7;
    11'b00001011100: data <= 32'hb398bbf6;
    11'b00001011101: data <= 32'h4015b9d5;
    11'b00001011110: data <= 32'h4166ab9e;
    11'b00001011111: data <= 32'h3d62b399;
    11'b00001100000: data <= 32'ha8d7bb0e;
    11'b00001100001: data <= 32'hb300b83f;
    11'b00001100010: data <= 32'hafff3980;
    11'b00001100011: data <= 32'hb9fd3a5b;
    11'b00001100100: data <= 32'hbd8fbc05;
    11'b00001100101: data <= 32'hbc27c15d;
    11'b00001100110: data <= 32'hb361c009;
    11'b00001100111: data <= 32'haec333fc;
    11'b00001101000: data <= 32'hb6d83e2a;
    11'b00001101001: data <= 32'hb0633c3c;
    11'b00001101010: data <= 32'h37bd3763;
    11'b00001101011: data <= 32'h1ddf3b85;
    11'b00001101100: data <= 32'hbe2f3e00;
    11'b00001101101: data <= 32'hc0253b40;
    11'b00001101110: data <= 32'hb523b316;
    11'b00001101111: data <= 32'h3ff5b833;
    11'b00001110000: data <= 32'h40c1acf4;
    11'b00001110001: data <= 32'h3c032c95;
    11'b00001110010: data <= 32'h3106ad40;
    11'b00001110011: data <= 32'h39f435bf;
    11'b00001110100: data <= 32'h3cc53c77;
    11'b00001110101: data <= 32'h3318390a;
    11'b00001110110: data <= 32'hbc6fbd7f;
    11'b00001110111: data <= 32'hbca0c1aa;
    11'b00001111000: data <= 32'hb181c008;
    11'b00001111001: data <= 32'h362fadcc;
    11'b00001111010: data <= 32'h321f384b;
    11'b00001111011: data <= 32'h2c7eb4da;
    11'b00001111100: data <= 32'h2c64b858;
    11'b00001111101: data <= 32'hb9b239e8;
    11'b00001111110: data <= 32'hc02b3f7b;
    11'b00001111111: data <= 32'hc0a93ce5;
    11'b00010000000: data <= 32'hb978b53c;
    11'b00010000001: data <= 32'h3c8abaad;
    11'b00010000010: data <= 32'h3cbeac0d;
    11'b00010000011: data <= 32'h30323967;
    11'b00010000100: data <= 32'h30583ac8;
    11'b00010000101: data <= 32'h3dc03c73;
    11'b00010000110: data <= 32'h3fc53deb;
    11'b00010000111: data <= 32'h381f3b0d;
    11'b00010001000: data <= 32'hbca7ba9d;
    11'b00010001001: data <= 32'hbc1bbff9;
    11'b00010001010: data <= 32'h37c1bdad;
    11'b00010001011: data <= 32'h3d74b4b1;
    11'b00010001100: data <= 32'h3bc4b71e;
    11'b00010001101: data <= 32'h35d0bdb8;
    11'b00010001110: data <= 32'h2d29bcb3;
    11'b00010001111: data <= 32'hb87d3921;
    11'b00010010000: data <= 32'hbeba3f2a;
    11'b00010010001: data <= 32'hc02439a8;
    11'b00010010010: data <= 32'hbc62bcb4;
    11'b00010010011: data <= 32'ha503bdf7;
    11'b00010010100: data <= 32'hb0fab11a;
    11'b00010010101: data <= 32'hb9903be6;
    11'b00010010110: data <= 32'h23423c78;
    11'b00010010111: data <= 32'h3e423c7d;
    11'b00010011000: data <= 32'h3f033e0c;
    11'b00010011001: data <= 32'ha9903dad;
    11'b00010011010: data <= 32'hbe6d358f;
    11'b00010011011: data <= 32'hbb30b929;
    11'b00010011100: data <= 32'h3c73b8bc;
    11'b00010011101: data <= 32'h4004b482;
    11'b00010011110: data <= 32'h3d2ebb06;
    11'b00010011111: data <= 32'h3860beb6;
    11'b00010100000: data <= 32'h38b8bc0a;
    11'b00010100001: data <= 32'h377a3ab6;
    11'b00010100010: data <= 32'hb81a3e04;
    11'b00010100011: data <= 32'hbdb1af8b;
    11'b00010100100: data <= 32'hbd3dc024;
    11'b00010100101: data <= 32'hba5abffd;
    11'b00010100110: data <= 32'hbab9b54f;
    11'b00010100111: data <= 32'hbb64397e;
    11'b00010101000: data <= 32'h0b383659;
    11'b00010101001: data <= 32'h3cf3342c;
    11'b00010101010: data <= 32'h3b653c8d;
    11'b00010101011: data <= 32'hbbee3f9f;
    11'b00010101100: data <= 32'hc0483dbe;
    11'b00010101101: data <= 32'hbb743622;
    11'b00010101110: data <= 32'h3c9fad59;
    11'b00010101111: data <= 32'h3ee0b14d;
    11'b00010110000: data <= 32'h3a70b932;
    11'b00010110001: data <= 32'h3707bc2a;
    11'b00010110010: data <= 32'h3d2ab2fd;
    11'b00010110011: data <= 32'h3f153d06;
    11'b00010110100: data <= 32'h39b73d52;
    11'b00010110101: data <= 32'hba77b851;
    11'b00010110110: data <= 32'hbd06c07d;
    11'b00010110111: data <= 32'hba75bf81;
    11'b00010111000: data <= 32'hb84fb68a;
    11'b00010111001: data <= 32'hb6ffacd6;
    11'b00010111010: data <= 32'h3228bb95;
    11'b00010111011: data <= 32'h3ac8bbfd;
    11'b00010111100: data <= 32'h322f38a7;
    11'b00010111101: data <= 32'hbe2f4025;
    11'b00010111110: data <= 32'hc0a03f41;
    11'b00010111111: data <= 32'hbc4e37e4;
    11'b00011000000: data <= 32'h3826b310;
    11'b00011000001: data <= 32'h3860afb9;
    11'b00011000010: data <= 32'hb500ae1e;
    11'b00011000011: data <= 32'h2b24b05c;
    11'b00011000100: data <= 32'h3f093855;
    11'b00011000101: data <= 32'h41233e42;
    11'b00011000110: data <= 32'h3cfc3da7;
    11'b00011000111: data <= 32'hb92bb1b8;
    11'b00011001000: data <= 32'hbc47bdb7;
    11'b00011001001: data <= 32'hb2debc32;
    11'b00011001010: data <= 32'h3605b40c;
    11'b00011001011: data <= 32'h3550ba8d;
    11'b00011001100: data <= 32'h3753c03b;
    11'b00011001101: data <= 32'h39edbf8e;
    11'b00011001110: data <= 32'h3212333c;
    11'b00011001111: data <= 32'hbcaf3f9d;
    11'b00011010000: data <= 32'hbf663d77;
    11'b00011010001: data <= 32'hbc95b424;
    11'b00011010010: data <= 32'hb64dbabd;
    11'b00011010011: data <= 32'hbaa7b292;
    11'b00011010100: data <= 32'hbda934a0;
    11'b00011010101: data <= 32'hb5ce340e;
    11'b00011010110: data <= 32'h3f0e38ad;
    11'b00011010111: data <= 32'h40e73db5;
    11'b00011011000: data <= 32'h3a8d3e8c;
    11'b00011011001: data <= 32'hbc163a0f;
    11'b00011011010: data <= 32'hbb77aa31;
    11'b00011011011: data <= 32'h372c2c21;
    11'b00011011100: data <= 32'h3c6c2da7;
    11'b00011011101: data <= 32'h398dbc67;
    11'b00011011110: data <= 32'h3816c0e0;
    11'b00011011111: data <= 32'h3bcebf90;
    11'b00011100000: data <= 32'h3bef3518;
    11'b00011100001: data <= 32'h25783e68;
    11'b00011100010: data <= 32'hbb4f3849;
    11'b00011100011: data <= 32'hbc07bcd1;
    11'b00011100100: data <= 32'hbbf0bd89;
    11'b00011100101: data <= 32'hbe61b48e;
    11'b00011100110: data <= 32'hbf6432f9;
    11'b00011100111: data <= 32'hb836b422;
    11'b00011101000: data <= 32'h3da1b49f;
    11'b00011101001: data <= 32'h3e8f3a37;
    11'b00011101010: data <= 32'hb0bb3f0b;
    11'b00011101011: data <= 32'hbe593e9a;
    11'b00011101100: data <= 32'hbb3d3c3e;
    11'b00011101101: data <= 32'h396a3a85;
    11'b00011101110: data <= 32'h3c04366f;
    11'b00011101111: data <= 32'h3289ba92;
    11'b00011110000: data <= 32'h30d3bf5a;
    11'b00011110001: data <= 32'h3d48bc76;
    11'b00011110010: data <= 32'h402d3a01;
    11'b00011110011: data <= 32'h3d503d90;
    11'b00011110100: data <= 32'ha67ba808;
    11'b00011110101: data <= 32'hb9aabe2f;
    11'b00011110110: data <= 32'hbb6ebd1d;
    11'b00011110111: data <= 32'hbd63b07f;
    11'b00011111000: data <= 32'hbdadb298;
    11'b00011111001: data <= 32'hb578bd92;
    11'b00011111010: data <= 32'h3bf4be80;
    11'b00011111011: data <= 32'h3a66acc6;
    11'b00011111100: data <= 32'hbacb3e90;
    11'b00011111101: data <= 32'hbf273fb3;
    11'b00011111110: data <= 32'hbaeb3cf6;
    11'b00011111111: data <= 32'h359e3a42;
    11'b00100000000: data <= 32'h293b37d6;
    11'b00100000001: data <= 32'hbbdeb402;
    11'b00100000010: data <= 32'hb84ebadb;
    11'b00100000011: data <= 32'h3de1b369;
    11'b00100000100: data <= 32'h41853c6a;
    11'b00100000101: data <= 32'h3fc73d4e;
    11'b00100000110: data <= 32'h34a32a23;
    11'b00100000111: data <= 32'hb6efbb78;
    11'b00100001000: data <= 32'hb509b648;
    11'b00100001001: data <= 32'hb633351e;
    11'b00100001010: data <= 32'hb86eb8e7;
    11'b00100001011: data <= 32'ha68ac0d5;
    11'b00100001100: data <= 32'h3a39c139;
    11'b00100001101: data <= 32'h3861b90a;
    11'b00100001110: data <= 32'hb9643d57;
    11'b00100001111: data <= 32'hbd233dc5;
    11'b00100010000: data <= 32'hb923378f;
    11'b00100010001: data <= 32'hb2fc2e73;
    11'b00100010010: data <= 32'hbcbb35bb;
    11'b00100010011: data <= 32'hc06332cd;
    11'b00100010100: data <= 32'hbccbb40c;
    11'b00100010101: data <= 32'h3d291fc4;
    11'b00100010110: data <= 32'h412e3b96;
    11'b00100010111: data <= 32'h3e1d3d1f;
    11'b00100011000: data <= 32'haea03926;
    11'b00100011001: data <= 32'hb53d3488;
    11'b00100011010: data <= 32'h36793ab3;
    11'b00100011011: data <= 32'h382f3b80;
    11'b00100011100: data <= 32'h9ca8b959;
    11'b00100011101: data <= 32'h28a8c158;
    11'b00100011110: data <= 32'h3a36c14e;
    11'b00100011111: data <= 32'h3c14b88b;
    11'b00100100000: data <= 32'h35893c24;
    11'b00100100001: data <= 32'hb36c3889;
    11'b00100100010: data <= 32'hb26cb8f9;
    11'b00100100011: data <= 32'hb86eb8eb;
    11'b00100100100: data <= 32'hbf7833ee;
    11'b00100100101: data <= 32'hc1633572;
    11'b00100100110: data <= 32'hbdc7b73e;
    11'b00100100111: data <= 32'h3b33b97b;
    11'b00100101000: data <= 32'h3ef43232;
    11'b00100101001: data <= 32'h37153c5d;
    11'b00100101010: data <= 32'hba963cfb;
    11'b00100101011: data <= 32'hb5833d35;
    11'b00100101100: data <= 32'h3a603ebc;
    11'b00100101101: data <= 32'h39b03d8e;
    11'b00100101110: data <= 32'hb4e0b508;
    11'b00100101111: data <= 32'hb686c010;
    11'b00100110000: data <= 32'h3a7abf28;
    11'b00100110001: data <= 32'h3f3a9ece;
    11'b00100110010: data <= 32'h3e353afe;
    11'b00100110011: data <= 32'h3a37b04c;
    11'b00100110100: data <= 32'h34a2bcec;
    11'b00100110101: data <= 32'hb5f2b9a5;
    11'b00100110110: data <= 32'hbe4f3734;
    11'b00100110111: data <= 32'hc06d32c9;
    11'b00100111000: data <= 32'hbcaabd13;
    11'b00100111001: data <= 32'h3843bfa1;
    11'b00100111010: data <= 32'h3a4bba5b;
    11'b00100111011: data <= 32'hb80939db;
    11'b00100111100: data <= 32'hbce73d6d;
    11'b00100111101: data <= 32'hb4603dbf;
    11'b00100111110: data <= 32'h39f43e8f;
    11'b00100111111: data <= 32'h2c2e3db8;
    11'b00101000000: data <= 32'hbd78333b;
    11'b00101000001: data <= 32'hbcf5bbab;
    11'b00101000010: data <= 32'h397db975;
    11'b00101000011: data <= 32'h408e3866;
    11'b00101000100: data <= 32'h403d3a72;
    11'b00101000101: data <= 32'h3c7db4d4;
    11'b00101000110: data <= 32'h3896bb76;
    11'b00101000111: data <= 32'h339f295f;
    11'b00101001000: data <= 32'hb8533c32;
    11'b00101001001: data <= 32'hbc9d2e53;
    11'b00101001010: data <= 32'hb936c01f;
    11'b00101001011: data <= 32'h3560c1af;
    11'b00101001100: data <= 32'h3507bdad;
    11'b00101001101: data <= 32'hb91f35bd;
    11'b00101001110: data <= 32'hbb033ac2;
    11'b00101001111: data <= 32'h2cc938d3;
    11'b00101010000: data <= 32'h37a53a61;
    11'b00101010001: data <= 32'hbb3e3c77;
    11'b00101010010: data <= 32'hc10b3939;
    11'b00101010011: data <= 32'hc002b125;
    11'b00101010100: data <= 32'h3620b06b;
    11'b00101010101: data <= 32'h4014388e;
    11'b00101010110: data <= 32'h3e943941;
    11'b00101010111: data <= 32'h38dda0cc;
    11'b00101011000: data <= 32'h3839232c;
    11'b00101011001: data <= 32'h3b563cd8;
    11'b00101011010: data <= 32'h384f3f33;
    11'b00101011011: data <= 32'hb4ee32fc;
    11'b00101011100: data <= 32'hb64fc06e;
    11'b00101011101: data <= 32'h3428c1aa;
    11'b00101011110: data <= 32'h37ddbd1e;
    11'b00101011111: data <= 32'h2e1a3165;
    11'b00101100000: data <= 32'h2eb3187a;
    11'b00101100001: data <= 32'h3958b91d;
    11'b00101100010: data <= 32'h35c2b25c;
    11'b00101100011: data <= 32'hbdd23a5f;
    11'b00101100100: data <= 32'hc1f73a9a;
    11'b00101100101: data <= 32'hc070ad2e;
    11'b00101100110: data <= 32'h2ac3b844;
    11'b00101100111: data <= 32'h3cd0ae29;
    11'b00101101000: data <= 32'h36d934ec;
    11'b00101101001: data <= 32'hb5f33575;
    11'b00101101010: data <= 32'h34bf3af6;
    11'b00101101011: data <= 32'h3d4f400f;
    11'b00101101100: data <= 32'h3be7408a;
    11'b00101101101: data <= 32'hb4d23885;
    11'b00101101110: data <= 32'hb9cdbe46;
    11'b00101101111: data <= 32'h307cbf6c;
    11'b00101110000: data <= 32'h3c04b7c7;
    11'b00101110001: data <= 32'h3c7332e0;
    11'b00101110010: data <= 32'h3c5fb997;
    11'b00101110011: data <= 32'h3ce7bdf7;
    11'b00101110100: data <= 32'h38bab8d4;
    11'b00101110101: data <= 32'hbc8c3adf;
    11'b00101110110: data <= 32'hc0d03aa8;
    11'b00101110111: data <= 32'hbefab8e4;
    11'b00101111000: data <= 32'haff5be2d;
    11'b00101111001: data <= 32'h3431bc41;
    11'b00101111010: data <= 32'hb9f9b11c;
    11'b00101111011: data <= 32'hbc5e3597;
    11'b00101111100: data <= 32'h32743ba0;
    11'b00101111101: data <= 32'h3d8b3fa7;
    11'b00101111110: data <= 32'h390c4051;
    11'b00101111111: data <= 32'hbc853b8e;
    11'b00110000000: data <= 32'hbe1eb810;
    11'b00110000001: data <= 32'hafb3b849;
    11'b00110000010: data <= 32'h3d4b363a;
    11'b00110000011: data <= 32'h3e69355e;
    11'b00110000100: data <= 32'h3d8fbba3;
    11'b00110000101: data <= 32'h3da5bdec;
    11'b00110000110: data <= 32'h3c52af0e;
    11'b00110000111: data <= 32'haf023da8;
    11'b00110001000: data <= 32'hbc9b3af8;
    11'b00110001001: data <= 32'hbb57bcdc;
    11'b00110001010: data <= 32'haf66c0c1;
    11'b00110001011: data <= 32'hb46cbea5;
    11'b00110001100: data <= 32'hbcabb7dd;
    11'b00110001101: data <= 32'hbc13add1;
    11'b00110001110: data <= 32'h37c42fa6;
    11'b00110001111: data <= 32'h3d1b3b30;
    11'b00110010000: data <= 32'hafc63e36;
    11'b00110010001: data <= 32'hc0533ca2;
    11'b00110010010: data <= 32'hc0903562;
    11'b00110010011: data <= 32'hb6f734a9;
    11'b00110010100: data <= 32'h3c6c39ab;
    11'b00110010101: data <= 32'h3c763475;
    11'b00110010110: data <= 32'h39d7ba85;
    11'b00110010111: data <= 32'h3c6bba32;
    11'b00110011000: data <= 32'h3e353b52;
    11'b00110011001: data <= 32'h3c014054;
    11'b00110011010: data <= 32'ha7af3c31;
    11'b00110011011: data <= 32'hb56fbd5a;
    11'b00110011100: data <= 32'hac53c0ae;
    11'b00110011101: data <= 32'hb3b2bda0;
    11'b00110011110: data <= 32'hb987b769;
    11'b00110011111: data <= 32'hb29ab9f9;
    11'b00110100000: data <= 32'h3c54bc95;
    11'b00110100001: data <= 32'h3d04b5d5;
    11'b00110100010: data <= 32'hb8c83b2f;
    11'b00110100011: data <= 32'hc12b3cb4;
    11'b00110100100: data <= 32'hc0d43854;
    11'b00110100101: data <= 32'hb8c63177;
    11'b00110100110: data <= 32'h36ce33af;
    11'b00110100111: data <= 32'hafc6ac55;
    11'b00110101000: data <= 32'hb804b8b5;
    11'b00110101001: data <= 32'h3849a7d8;
    11'b00110101010: data <= 32'h3f213ebc;
    11'b00110101011: data <= 32'h3e3a412b;
    11'b00110101100: data <= 32'h343b3d1f;
    11'b00110101101: data <= 32'hb708ba7d;
    11'b00110101110: data <= 32'hb14cbd5e;
    11'b00110101111: data <= 32'h302ab612;
    11'b00110110000: data <= 32'h31b3ad96;
    11'b00110110001: data <= 32'h39c1bd05;
    11'b00110110010: data <= 32'h3e7bc02e;
    11'b00110110011: data <= 32'h3db3bc43;
    11'b00110110100: data <= 32'hb5c5398f;
    11'b00110110101: data <= 32'hbff23c88;
    11'b00110110110: data <= 32'hbeed3114;
    11'b00110110111: data <= 32'hb76eb946;
    11'b00110111000: data <= 32'hb525b92c;
    11'b00110111001: data <= 32'hbd82b84d;
    11'b00110111010: data <= 32'hbe1bb895;
    11'b00110111011: data <= 32'h30a22df6;
    11'b00110111100: data <= 32'h3f0b3e31;
    11'b00110111101: data <= 32'h3d624099;
    11'b00110111110: data <= 32'hb5b13d87;
    11'b00110111111: data <= 32'hbc8c2bff;
    11'b00111000000: data <= 32'hb70e2a96;
    11'b00111000001: data <= 32'h36923a6c;
    11'b00111000010: data <= 32'h395a35aa;
    11'b00111000011: data <= 32'h3bfebd9b;
    11'b00111000100: data <= 32'h3eb0c070;
    11'b00111000101: data <= 32'h3eb7ba75;
    11'b00111000110: data <= 32'h37ed3c74;
    11'b00111000111: data <= 32'hb9513cbf;
    11'b00111001000: data <= 32'hb8cdb5ee;
    11'b00111001001: data <= 32'haf7dbdd2;
    11'b00111001010: data <= 32'hb9cdbce7;
    11'b00111001011: data <= 32'hbfbdba3b;
    11'b00111001100: data <= 32'hbedabaa2;
    11'b00111001101: data <= 32'h341bb8bb;
    11'b00111001110: data <= 32'h3e9e379f;
    11'b00111001111: data <= 32'h398a3d9c;
    11'b00111010000: data <= 32'hbd443d01;
    11'b00111010001: data <= 32'hbf783a06;
    11'b00111010010: data <= 32'hb9a03c0b;
    11'b00111010011: data <= 32'h352e3da2;
    11'b00111010100: data <= 32'h34d93810;
    11'b00111010101: data <= 32'h34b3bcfc;
    11'b00111010110: data <= 32'h3c66be84;
    11'b00111010111: data <= 32'h3f412f4e;
    11'b00111011000: data <= 32'h3dc33f54;
    11'b00111011001: data <= 32'h38b03d5d;
    11'b00111011010: data <= 32'h349eb897;
    11'b00111011011: data <= 32'h31d4be0a;
    11'b00111011100: data <= 32'hb936bb7e;
    11'b00111011101: data <= 32'hbe59b828;
    11'b00111011110: data <= 32'hbc26bcae;
    11'b00111011111: data <= 32'h3a6fbec1;
    11'b00111100000: data <= 32'h3e86bb46;
    11'b00111100001: data <= 32'h31ca36b5;
    11'b00111100010: data <= 32'hbf333bd4;
    11'b00111100011: data <= 32'hbfe73b26;
    11'b00111100100: data <= 32'hb9643c20;
    11'b00111100101: data <= 32'hace23c76;
    11'b00111100110: data <= 32'hba2e3394;
    11'b00111100111: data <= 32'hbc36bc20;
    11'b00111101000: data <= 32'h3247bb1b;
    11'b00111101001: data <= 32'h3ee83b57;
    11'b00111101010: data <= 32'h3fa1407a;
    11'b00111101011: data <= 32'h3c1e3db3;
    11'b00111101100: data <= 32'h3676b497;
    11'b00111101101: data <= 32'h323fb949;
    11'b00111101110: data <= 32'hb4b33238;
    11'b00111101111: data <= 32'hba0931ee;
    11'b00111110000: data <= 32'haeb1bd62;
    11'b00111110001: data <= 32'h3d5cc10c;
    11'b00111110010: data <= 32'h3ecabf10;
    11'b00111110011: data <= 32'h330ca8e1;
    11'b00111110100: data <= 32'hbd5a3a41;
    11'b00111110101: data <= 32'hbcd0381f;
    11'b00111110110: data <= 32'hb3513446;
    11'b00111110111: data <= 32'hb7ce3410;
    11'b00111111000: data <= 32'hbfa1b37c;
    11'b00111111001: data <= 32'hc079bb9a;
    11'b00111111010: data <= 32'hb7c0b8e1;
    11'b00111111011: data <= 32'h3e063b3d;
    11'b00111111100: data <= 32'h3ebc3f8a;
    11'b00111111101: data <= 32'h37ff3cf6;
    11'b00111111110: data <= 32'hb35c342a;
    11'b00111111111: data <= 32'hac9238d9;
    11'b01000000000: data <= 32'h25533e29;
    11'b01000000001: data <= 32'hb0db3b90;
    11'b01000000010: data <= 32'h348bbd03;
    11'b01000000011: data <= 32'h3d62c13e;
    11'b01000000100: data <= 32'h3ecdbe7a;
    11'b01000000101: data <= 32'h3a253466;
    11'b01000000110: data <= 32'hb0ab3a71;
    11'b01000000111: data <= 32'h2ddaa72c;
    11'b01000001000: data <= 32'h3755b8ce;
    11'b01000001001: data <= 32'hb8f5b6ad;
    11'b01000001010: data <= 32'hc0d5b73f;
    11'b01000001011: data <= 32'hc11dbbff;
    11'b01000001100: data <= 32'hb82fbc0d;
    11'b01000001101: data <= 32'h3d5ba894;
    11'b01000001110: data <= 32'h3c193aa6;
    11'b01000001111: data <= 32'hb7f43a13;
    11'b01000010000: data <= 32'hbc1f393b;
    11'b01000010001: data <= 32'hb5493e06;
    11'b01000010010: data <= 32'h2e25409a;
    11'b01000010011: data <= 32'hb44c3d30;
    11'b01000010100: data <= 32'hb4a3bc00;
    11'b01000010101: data <= 32'h3915c00e;
    11'b01000010110: data <= 32'h3df5b98c;
    11'b01000010111: data <= 32'h3d9b3c25;
    11'b01000011000: data <= 32'h3c243bbb;
    11'b01000011001: data <= 32'h3ca0b5a5;
    11'b01000011010: data <= 32'h3c02baf6;
    11'b01000011011: data <= 32'hb687b422;
    11'b01000011100: data <= 32'hc020ad2d;
    11'b01000011101: data <= 32'hbfa3bc0f;
    11'b01000011110: data <= 32'h2896bf2d;
    11'b01000011111: data <= 32'h3d4abd5e;
    11'b01000100000: data <= 32'h36c9b57f;
    11'b01000100001: data <= 32'hbca53259;
    11'b01000100010: data <= 32'hbd1138ec;
    11'b01000100011: data <= 32'hb2f13e10;
    11'b01000100100: data <= 32'ha05a4024;
    11'b01000100101: data <= 32'hbc243c37;
    11'b01000100110: data <= 32'hbe32ba42;
    11'b01000100111: data <= 32'hb775bce4;
    11'b01000101000: data <= 32'h3c523426;
    11'b01000101001: data <= 32'h3e9a3e45;
    11'b01000101010: data <= 32'h3dda3bf5;
    11'b01000101011: data <= 32'h3d7cb536;
    11'b01000101100: data <= 32'h3c5fb508;
    11'b01000101101: data <= 32'ha71d3a3a;
    11'b01000101110: data <= 32'hbcbf3a8c;
    11'b01000101111: data <= 32'hbadebac8;
    11'b01000110000: data <= 32'h3981c0c2;
    11'b01000110001: data <= 32'h3d6fc05a;
    11'b01000110010: data <= 32'h33b2bb7e;
    11'b01000110011: data <= 32'hbbcfb02c;
    11'b01000110100: data <= 32'hb8c631e9;
    11'b01000110101: data <= 32'h369039c7;
    11'b01000110110: data <= 32'hac9e3c81;
    11'b01000110111: data <= 32'hbf9b37b5;
    11'b01000111000: data <= 32'hc169b98b;
    11'b01000111001: data <= 32'hbd41ba10;
    11'b01000111010: data <= 32'h3962380a;
    11'b01000111011: data <= 32'h3d5a3d4e;
    11'b01000111100: data <= 32'h3b4e392f;
    11'b01000111101: data <= 32'h398cafb6;
    11'b01000111110: data <= 32'h3a013964;
    11'b01000111111: data <= 32'h34864030;
    11'b01001000000: data <= 32'hb6e73f16;
    11'b01001000001: data <= 32'hb362b826;
    11'b01001000010: data <= 32'h3a8fc0b5;
    11'b01001000011: data <= 32'h3cebc008;
    11'b01001000100: data <= 32'h3764b8f9;
    11'b01001000101: data <= 32'hac49ac6f;
    11'b01001000110: data <= 32'h394db5ad;
    11'b01001000111: data <= 32'h3d3cb44a;
    11'b01001001000: data <= 32'h2cac33a3;
    11'b01001001001: data <= 32'hc0813007;
    11'b01001001010: data <= 32'hc209b924;
    11'b01001001011: data <= 32'hbd94badc;
    11'b01001001100: data <= 32'h37f3b0d4;
    11'b01001001101: data <= 32'h395d3515;
    11'b01001001110: data <= 32'hb1d4aaca;
    11'b01001001111: data <= 32'hb4bea882;
    11'b01001010000: data <= 32'h359c3d8d;
    11'b01001010001: data <= 32'h36cc41b5;
    11'b01001010010: data <= 32'hb464406b;
    11'b01001010011: data <= 32'hb82bb28e;
    11'b01001010100: data <= 32'h3178beeb;
    11'b01001010101: data <= 32'h3a69bc0c;
    11'b01001010110: data <= 32'h3a2134c5;
    11'b01001010111: data <= 32'h3b3f3340;
    11'b01001011000: data <= 32'h3ef1b9c3;
    11'b01001011001: data <= 32'h3ff1ba3f;
    11'b01001011010: data <= 32'h36642f91;
    11'b01001011011: data <= 32'hbf6336a6;
    11'b01001011100: data <= 32'hc09eb752;
    11'b01001011101: data <= 32'hb9b5bd35;
    11'b01001011110: data <= 32'h38c8bcec;
    11'b01001011111: data <= 32'h29dabaf3;
    11'b01001100000: data <= 32'hbc3fba4e;
    11'b01001100001: data <= 32'hba6fb3bc;
    11'b01001100010: data <= 32'h35c43d47;
    11'b01001100011: data <= 32'h37e9412a;
    11'b01001100100: data <= 32'hb9aa3f8d;
    11'b01001100101: data <= 32'hbe27acfc;
    11'b01001100110: data <= 32'hbb85bb43;
    11'b01001100111: data <= 32'h31f53038;
    11'b01001101000: data <= 32'h3a633c5e;
    11'b01001101001: data <= 32'h3ceb360a;
    11'b01001101010: data <= 32'h3fb9bab3;
    11'b01001101011: data <= 32'h4018b85d;
    11'b01001101100: data <= 32'h39cf3b37;
    11'b01001101101: data <= 32'hbb9e3d41;
    11'b01001101110: data <= 32'hbc5dac45;
    11'b01001101111: data <= 32'h31ffbe86;
    11'b01001110000: data <= 32'h3a2bbfbf;
    11'b01001110001: data <= 32'hb40dbdda;
    11'b01001110010: data <= 32'hbcb9bc92;
    11'b01001110011: data <= 32'hb658b954;
    11'b01001110100: data <= 32'h3bc43803;
    11'b01001110101: data <= 32'h39453dfa;
    11'b01001110110: data <= 32'hbd283c59;
    11'b01001110111: data <= 32'hc117b041;
    11'b01001111000: data <= 32'hbf3ab5a6;
    11'b01001111001: data <= 32'hb4d53955;
    11'b01001111010: data <= 32'h37093c7c;
    11'b01001111011: data <= 32'h39252c6b;
    11'b01001111100: data <= 32'h3c8dbad4;
    11'b01001111101: data <= 32'h3e083083;
    11'b01001111110: data <= 32'h3b2a4019;
    11'b01001111111: data <= 32'hb01c4099;
    11'b01010000000: data <= 32'hb2143647;
    11'b01010000001: data <= 32'h38cfbe05;
    11'b01010000010: data <= 32'h39a5bee5;
    11'b01010000011: data <= 32'hb3a5bc40;
    11'b01010000100: data <= 32'hb8aabb6d;
    11'b01010000101: data <= 32'h396fbc53;
    11'b01010000110: data <= 32'h3fa3b855;
    11'b01010000111: data <= 32'h3bca35a3;
    11'b01010001000: data <= 32'hbdfa3716;
    11'b01010001001: data <= 32'hc194b195;
    11'b01010001010: data <= 32'hbf55b443;
    11'b01010001011: data <= 32'hb605353a;
    11'b01010001100: data <= 32'hb0463509;
    11'b01010001101: data <= 32'hb7f3b95e;
    11'b01010001110: data <= 32'had75bbbe;
    11'b01010001111: data <= 32'h3a91395a;
    11'b01010010000: data <= 32'h3b5d4175;
    11'b01010010001: data <= 32'h3216416e;
    11'b01010010010: data <= 32'hb1353946;
    11'b01010010011: data <= 32'h319abb7e;
    11'b01010010100: data <= 32'h33feb965;
    11'b01010010101: data <= 32'hb0e62c29;
    11'b01010010110: data <= 32'h3171b5b8;
    11'b01010010111: data <= 32'h3ea3bd40;
    11'b01010011000: data <= 32'h4130bcc4;
    11'b01010011001: data <= 32'h3d3dad52;
    11'b01010011010: data <= 32'hbc6737c6;
    11'b01010011011: data <= 32'hc0112443;
    11'b01010011100: data <= 32'hbbc4b7c4;
    11'b01010011101: data <= 32'ha5fdb80a;
    11'b01010011110: data <= 32'hb8f8ba20;
    11'b01010011111: data <= 32'hbdf9bdc4;
    11'b01010100000: data <= 32'hbb39bcf5;
    11'b01010100001: data <= 32'h387e388e;
    11'b01010100010: data <= 32'h3bbd40d0;
    11'b01010100011: data <= 32'ha5de407d;
    11'b01010100100: data <= 32'hbb48388c;
    11'b01010100101: data <= 32'hba7fb3d1;
    11'b01010100110: data <= 32'hb6b53893;
    11'b01010100111: data <= 32'hb3933ca4;
    11'b01010101000: data <= 32'h36bb2d17;
    11'b01010101001: data <= 32'h3f39bd83;
    11'b01010101010: data <= 32'h4117bca8;
    11'b01010101011: data <= 32'h3dd9369e;
    11'b01010101100: data <= 32'hb5193cf3;
    11'b01010101101: data <= 32'hb9c5377b;
    11'b01010101110: data <= 32'h3317b945;
    11'b01010101111: data <= 32'h3726bc64;
    11'b01010110000: data <= 32'hbabcbd3e;
    11'b01010110001: data <= 32'hbf3abeec;
    11'b01010110010: data <= 32'hba5dbe2b;
    11'b01010110011: data <= 32'h3bffb121;
    11'b01010110100: data <= 32'h3cbe3cf2;
    11'b01010110101: data <= 32'hb6bb3cac;
    11'b01010110110: data <= 32'hbf1232d6;
    11'b01010110111: data <= 32'hbe8132c9;
    11'b01010111000: data <= 32'hbb143d26;
    11'b01010111001: data <= 32'hb8423e03;
    11'b01010111010: data <= 32'haef0a72a;
    11'b01010111011: data <= 32'h3b82bdbb;
    11'b01010111100: data <= 32'h3f07b96b;
    11'b01010111101: data <= 32'h3d5d3d87;
    11'b01010111110: data <= 32'h364c4053;
    11'b01010111111: data <= 32'h35953b85;
    11'b01011000000: data <= 32'h3baeb84d;
    11'b01011000001: data <= 32'h38e6bb41;
    11'b01011000010: data <= 32'hbac3bac8;
    11'b01011000011: data <= 32'hbdaabd36;
    11'b01011000100: data <= 32'h2cbcbec3;
    11'b01011000101: data <= 32'h3f77bc5a;
    11'b01011000110: data <= 32'h3e2aac1a;
    11'b01011000111: data <= 32'hb8a33213;
    11'b01011001000: data <= 32'hbffeadbd;
    11'b01011001001: data <= 32'hbe6634a9;
    11'b01011001010: data <= 32'hba513ca3;
    11'b01011001011: data <= 32'hbb013b6f;
    11'b01011001100: data <= 32'hbc8eb970;
    11'b01011001101: data <= 32'hb6e1be6b;
    11'b01011001110: data <= 32'h39e1b3a1;
    11'b01011001111: data <= 32'h3c514008;
    11'b01011010000: data <= 32'h396d4112;
    11'b01011010001: data <= 32'h38b63c56;
    11'b01011010010: data <= 32'h3a5db0e0;
    11'b01011010011: data <= 32'h34542a0e;
    11'b01011010100: data <= 32'hba96369c;
    11'b01011010101: data <= 32'hba4cb683;
    11'b01011010110: data <= 32'h3bd7be7c;
    11'b01011010111: data <= 32'h4108beb8;
    11'b01011011000: data <= 32'h3f34b9af;
    11'b01011011001: data <= 32'hb515ab63;
    11'b01011011010: data <= 32'hbd45a9dd;
    11'b01011011011: data <= 32'hb8f2303c;
    11'b01011011100: data <= 32'hb03537ae;
    11'b01011011101: data <= 32'hbc40aa36;
    11'b01011011110: data <= 32'hc01fbdb0;
    11'b01011011111: data <= 32'hbdd1bf60;
    11'b01011100000: data <= 32'h3116b418;
    11'b01011100001: data <= 32'h3b863efe;
    11'b01011100010: data <= 32'h38173fda;
    11'b01011100011: data <= 32'h243639bd;
    11'b01011100100: data <= 32'hab533408;
    11'b01011100101: data <= 32'hb5e83cda;
    11'b01011100110: data <= 32'hbb4f3ed8;
    11'b01011100111: data <= 32'hb80735e0;
    11'b01011101000: data <= 32'h3ca4bddb;
    11'b01011101001: data <= 32'h40c6beb7;
    11'b01011101010: data <= 32'h3edeb67b;
    11'b01011101011: data <= 32'h32683833;
    11'b01011101100: data <= 32'had8435cf;
    11'b01011101101: data <= 32'h3a2d9e0d;
    11'b01011101110: data <= 32'h3984ae69;
    11'b01011101111: data <= 32'hbc1fb8dd;
    11'b01011110000: data <= 32'hc0c2be9e;
    11'b01011110001: data <= 32'hbe34bfd4;
    11'b01011110010: data <= 32'h3643ba09;
    11'b01011110011: data <= 32'h3c5f393c;
    11'b01011110100: data <= 32'h31403994;
    11'b01011110101: data <= 32'hba4e1fdb;
    11'b01011110110: data <= 32'hbae836f2;
    11'b01011110111: data <= 32'hba673fab;
    11'b01011111000: data <= 32'hbc48408a;
    11'b01011111001: data <= 32'hbab93805;
    11'b01011111010: data <= 32'h35debdb0;
    11'b01011111011: data <= 32'h3db4bcfc;
    11'b01011111100: data <= 32'h3cfd379c;
    11'b01011111101: data <= 32'h39023daa;
    11'b01011111110: data <= 32'h3bae3a88;
    11'b01011111111: data <= 32'h3ef426ab;
    11'b01100000000: data <= 32'h3c8aab4a;
    11'b01100000001: data <= 32'hbb36b2c3;
    11'b01100000010: data <= 32'hc014bc4f;
    11'b01100000011: data <= 32'hba61bf1c;
    11'b01100000100: data <= 32'h3cc7bd93;
    11'b01100000101: data <= 32'h3dbeb8e6;
    11'b01100000110: data <= 32'ha943b826;
    11'b01100000111: data <= 32'hbc7db8e4;
    11'b01100001000: data <= 32'hbb293584;
    11'b01100001001: data <= 32'hb8ae3f55;
    11'b01100001010: data <= 32'hbc7c3f5b;
    11'b01100001011: data <= 32'hbe60aac5;
    11'b01100001100: data <= 32'hbbb0be4f;
    11'b01100001101: data <= 32'h3133ba59;
    11'b01100001110: data <= 32'h391e3cb1;
    11'b01100001111: data <= 32'h39a73f59;
    11'b01100010000: data <= 32'h3cf23af8;
    11'b01100010001: data <= 32'h3efc3132;
    11'b01100010010: data <= 32'h3b6d3923;
    11'b01100010011: data <= 32'hbace3c04;
    11'b01100010100: data <= 32'hbdb02b07;
    11'b01100010101: data <= 32'h305bbd62;
    11'b01100010110: data <= 32'h3f89bf02;
    11'b01100010111: data <= 32'h3e8abd25;
    11'b01100011000: data <= 32'h249cbbbd;
    11'b01100011001: data <= 32'hb958b9fc;
    11'b01100011010: data <= 32'h28de3047;
    11'b01100011011: data <= 32'h34ba3cba;
    11'b01100011100: data <= 32'hbb8a3af2;
    11'b01100011101: data <= 32'hc086ba8e;
    11'b01100011110: data <= 32'hc002bf20;
    11'b01100011111: data <= 32'hb920b93b;
    11'b01100100000: data <= 32'h34593c69;
    11'b01100100001: data <= 32'h374b3d43;
    11'b01100100010: data <= 32'h399e34dc;
    11'b01100100011: data <= 32'h3b7e32d1;
    11'b01100100100: data <= 32'h348f3e2f;
    11'b01100100101: data <= 32'hbb6440a1;
    11'b01100100110: data <= 32'hbc183c4f;
    11'b01100100111: data <= 32'h37bebb4e;
    11'b01100101000: data <= 32'h3f3fbe86;
    11'b01100101001: data <= 32'h3d83bc18;
    11'b01100101010: data <= 32'h328ab775;
    11'b01100101011: data <= 32'h34d9b5de;
    11'b01100101100: data <= 32'h3dbea279;
    11'b01100101101: data <= 32'h3d843833;
    11'b01100101110: data <= 32'hb8c8317f;
    11'b01100101111: data <= 32'hc0dbbc76;
    11'b01100110000: data <= 32'hc04abf06;
    11'b01100110001: data <= 32'hb83cbacf;
    11'b01100110010: data <= 32'h35b4342c;
    11'b01100110011: data <= 32'h2e252a2f;
    11'b01100110100: data <= 32'hb0adb966;
    11'b01100110101: data <= 32'h26702b12;
    11'b01100110110: data <= 32'hb2d34023;
    11'b01100110111: data <= 32'hbbd641d7;
    11'b01100111000: data <= 32'hbc633d7d;
    11'b01100111001: data <= 32'hac6fba0d;
    11'b01100111010: data <= 32'h3adabcae;
    11'b01100111011: data <= 32'h3925aff1;
    11'b01100111100: data <= 32'h346337ef;
    11'b01100111101: data <= 32'h3c9630cc;
    11'b01100111110: data <= 32'h40e8aa20;
    11'b01100111111: data <= 32'h400b358b;
    11'b01101000000: data <= 32'hb4df3579;
    11'b01101000001: data <= 32'hc012b87b;
    11'b01101000010: data <= 32'hbd91bd4e;
    11'b01101000011: data <= 32'h34f0bc86;
    11'b01101000100: data <= 32'h39fbba50;
    11'b01101000101: data <= 32'hb0d4bce4;
    11'b01101000110: data <= 32'hb94bbe1d;
    11'b01101000111: data <= 32'hb2e4b3ec;
    11'b01101001000: data <= 32'ha8b33fa1;
    11'b01101001001: data <= 32'hba784102;
    11'b01101001010: data <= 32'hbdff3a92;
    11'b01101001011: data <= 32'hbcafbb7e;
    11'b01101001100: data <= 32'hb766b985;
    11'b01101001101: data <= 32'hb34d39c1;
    11'b01101001110: data <= 32'h2e203c6c;
    11'b01101001111: data <= 32'h3d483426;
    11'b01101010000: data <= 32'h40fcae48;
    11'b01101010001: data <= 32'h3f7539b8;
    11'b01101010010: data <= 32'hb3e43d4f;
    11'b01101010011: data <= 32'hbd9438f8;
    11'b01101010100: data <= 32'hb57cb8e6;
    11'b01101010101: data <= 32'h3ca9bcc3;
    11'b01101010110: data <= 32'h3c0fbd58;
    11'b01101010111: data <= 32'hb3bfbee3;
    11'b01101011000: data <= 32'hb815bf0e;
    11'b01101011001: data <= 32'h37cdb80e;
    11'b01101011010: data <= 32'h3b0b3cea;
    11'b01101011011: data <= 32'hb57b3dc9;
    11'b01101011100: data <= 32'hbf5fadb8;
    11'b01101011101: data <= 32'hc022bcdd;
    11'b01101011110: data <= 32'hbd54b6ee;
    11'b01101011111: data <= 32'hb9f93b60;
    11'b01101100000: data <= 32'hb4093a7f;
    11'b01101100001: data <= 32'h3a02b53f;
    11'b01101100010: data <= 32'h3e7fb537;
    11'b01101100011: data <= 32'h3c6d3d1f;
    11'b01101100100: data <= 32'hb65140f2;
    11'b01101100101: data <= 32'hbb433ee4;
    11'b01101100110: data <= 32'h33ff24d3;
    11'b01101100111: data <= 32'h3d45bb5e;
    11'b01101101000: data <= 32'h3a11bc18;
    11'b01101101001: data <= 32'hb50cbcc3;
    11'b01101101010: data <= 32'h2fb8bd3b;
    11'b01101101011: data <= 32'h3ed6b8b8;
    11'b01101101100: data <= 32'h4019380f;
    11'b01101101101: data <= 32'h33ae3842;
    11'b01101101110: data <= 32'hbf3db8dd;
    11'b01101101111: data <= 32'hc047bcdc;
    11'b01101110000: data <= 32'hbce1b659;
    11'b01101110001: data <= 32'hb91836a1;
    11'b01101110010: data <= 32'hb896b453;
    11'b01101110011: data <= 32'hb0bcbd94;
    11'b01101110100: data <= 32'h3833ba01;
    11'b01101110101: data <= 32'h36493e41;
    11'b01101110110: data <= 32'hb7ff41fc;
    11'b01101110111: data <= 32'hba3a4017;
    11'b01101111000: data <= 32'h2551328e;
    11'b01101111001: data <= 32'h3878b763;
    11'b01101111010: data <= 32'hab8aad0b;
    11'b01101111011: data <= 32'hb83dac88;
    11'b01101111100: data <= 32'h398fb8b8;
    11'b01101111101: data <= 32'h4142b873;
    11'b01101111110: data <= 32'h417f3112;
    11'b01101111111: data <= 32'h38f13648;
    11'b01110000000: data <= 32'hbd82b42a;
    11'b01110000001: data <= 32'hbd5bb9c1;
    11'b01110000010: data <= 32'hb416b62d;
    11'b01110000011: data <= 32'hac67b57e;
    11'b01110000100: data <= 32'hb9f1bdbc;
    11'b01110000101: data <= 32'hba6dc0a9;
    11'b01110000110: data <= 32'ha03fbcc4;
    11'b01110000111: data <= 32'h35933d44;
    11'b01110001000: data <= 32'hb497410e;
    11'b01110001001: data <= 32'hbb2d3d9a;
    11'b01110001010: data <= 32'hba2eaf8f;
    11'b01110001011: data <= 32'hb921ab15;
    11'b01110001100: data <= 32'hbc223b0a;
    11'b01110001101: data <= 32'hbb2c3a7f;
    11'b01110001110: data <= 32'h39ebb3fc;
    11'b01110001111: data <= 32'h413bb8f3;
    11'b01110010000: data <= 32'h4111342e;
    11'b01110010001: data <= 32'h389c3c3e;
    11'b01110010010: data <= 32'hba5a3a4d;
    11'b01110010011: data <= 32'hb21c2f0e;
    11'b01110010100: data <= 32'h3ad5b2e8;
    11'b01110010101: data <= 32'h36f0b9c5;
    11'b01110010110: data <= 32'hba8bbf83;
    11'b01110010111: data <= 32'hbb25c119;
    11'b01110011000: data <= 32'h3600bd9c;
    11'b01110011001: data <= 32'h3c753964;
    11'b01110011010: data <= 32'h34b13d87;
    11'b01110011011: data <= 32'hbbd83426;
    11'b01110011100: data <= 32'hbddab90b;
    11'b01110011101: data <= 32'hbdd13134;
    11'b01110011110: data <= 32'hbe4f3d33;
    11'b01110011111: data <= 32'hbd043ab1;
    11'b01110100000: data <= 32'h3196b954;
    11'b01110100001: data <= 32'h3eadbb97;
    11'b01110100010: data <= 32'h3e4b3868;
    11'b01110100011: data <= 32'h32973fe3;
    11'b01110100100: data <= 32'hb5ca3f4f;
    11'b01110100101: data <= 32'h38c63a72;
    11'b01110100110: data <= 32'h3d4a2fdd;
    11'b01110100111: data <= 32'h35e7b607;
    11'b01110101000: data <= 32'hbbc9bd1e;
    11'b01110101001: data <= 32'hb855bfb4;
    11'b01110101010: data <= 32'h3d5dbd25;
    11'b01110101011: data <= 32'h406d2312;
    11'b01110101100: data <= 32'h3bc534ac;
    11'b01110101101: data <= 32'hba95b894;
    11'b01110101110: data <= 32'hbdddbabd;
    11'b01110101111: data <= 32'hbd233417;
    11'b01110110000: data <= 32'hbd603c44;
    11'b01110110001: data <= 32'hbda526d4;
    11'b01110110010: data <= 32'hb952be9b;
    11'b01110110011: data <= 32'h3699bdf4;
    11'b01110110100: data <= 32'h386b394e;
    11'b01110110101: data <= 32'hb03140c6;
    11'b01110110110: data <= 32'hb2814033;
    11'b01110110111: data <= 32'h39123b55;
    11'b01110111000: data <= 32'h3acf3779;
    11'b01110111001: data <= 32'hb59f382b;
    11'b01110111010: data <= 32'hbd40a524;
    11'b01110111011: data <= 32'hb193bb52;
    11'b01110111100: data <= 32'h403fbc08;
    11'b01110111101: data <= 32'h41beb566;
    11'b01110111110: data <= 32'h3d4aae94;
    11'b01110111111: data <= 32'hb735b83b;
    11'b01111000000: data <= 32'hb986b777;
    11'b01111000001: data <= 32'hb24b3642;
    11'b01111000010: data <= 32'hb8103858;
    11'b01111000011: data <= 32'hbd58bbcb;
    11'b01111000100: data <= 32'hbd34c11b;
    11'b01111000101: data <= 32'hb5ccbfcc;
    11'b01111000110: data <= 32'h320b36bf;
    11'b01111000111: data <= 32'hac543fae;
    11'b01111001000: data <= 32'hb2aa3d66;
    11'b01111001001: data <= 32'h2df335bb;
    11'b01111001010: data <= 32'hb12a3925;
    11'b01111001011: data <= 32'hbd2f3dca;
    11'b01111001100: data <= 32'hbef73c5c;
    11'b01111001101: data <= 32'hb1abb3d4;
    11'b01111001110: data <= 32'h402bbb1e;
    11'b01111001111: data <= 32'h4123b53e;
    11'b01111010000: data <= 32'h3c5834d4;
    11'b01111010001: data <= 32'hac9034e4;
    11'b01111010010: data <= 32'h36c13543;
    11'b01111010011: data <= 32'h3c813942;
    11'b01111010100: data <= 32'h35433431;
    11'b01111010101: data <= 32'hbcd0bd7a;
    11'b01111010110: data <= 32'hbdd6c169;
    11'b01111010111: data <= 32'hb3e4c006;
    11'b01111011000: data <= 32'h39b6aae4;
    11'b01111011001: data <= 32'h376a3a71;
    11'b01111011010: data <= 32'hb191201d;
    11'b01111011011: data <= 32'hb750b7c5;
    11'b01111011100: data <= 32'hbb393910;
    11'b01111011101: data <= 32'hbf303fa6;
    11'b01111011110: data <= 32'hc0023d87;
    11'b01111011111: data <= 32'hb8f2b64c;
    11'b01111100000: data <= 32'h3ca5bc95;
    11'b01111100001: data <= 32'h3db2b13f;
    11'b01111100010: data <= 32'h36543c26;
    11'b01111100011: data <= 32'h2fe03cff;
    11'b01111100100: data <= 32'h3cf23c01;
    11'b01111100101: data <= 32'h3f733ba8;
    11'b01111100110: data <= 32'h3875383e;
    11'b01111100111: data <= 32'hbd05ba46;
    11'b01111101000: data <= 32'hbcebbfb0;
    11'b01111101001: data <= 32'h3821be65;
    11'b01111101010: data <= 32'h3ec5b7a0;
    11'b01111101011: data <= 32'h3c85b4c8;
    11'b01111101100: data <= 32'h9ca1bc5e;
    11'b01111101101: data <= 32'hb7c6bc0f;
    11'b01111101110: data <= 32'hb9e038ba;
    11'b01111101111: data <= 32'hbdba3f2b;
    11'b01111110000: data <= 32'hbf9a3a5d;
    11'b01111110001: data <= 32'hbceebced;
    11'b01111110010: data <= 32'hae7cbeb6;
    11'b01111110011: data <= 32'h306aaea0;
    11'b01111110100: data <= 32'hb47b3db8;
    11'b01111110101: data <= 32'h2f6a3e0b;
    11'b01111110110: data <= 32'h3d7f3c0d;
    11'b01111110111: data <= 32'h3e873c59;
    11'b01111111000: data <= 32'h23303ce9;
    11'b01111111001: data <= 32'hbe51379e;
    11'b01111111010: data <= 32'hbb8cb93c;
    11'b01111111011: data <= 32'h3cf2bbc1;
    11'b01111111100: data <= 32'h40a6b912;
    11'b01111111101: data <= 32'h3da7ba3d;
    11'b01111111110: data <= 32'h329cbd3a;
    11'b01111111111: data <= 32'h2fddbacd;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    