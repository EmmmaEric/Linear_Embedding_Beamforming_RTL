
module memory_rom_51(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3e4cb007;
    11'b00000000001: data <= 32'h3b5db08b;
    11'b00000000010: data <= 32'hbb202a7e;
    11'b00000000011: data <= 32'hbefbb964;
    11'b00000000100: data <= 32'hb5a3bebd;
    11'b00000000101: data <= 32'h3e61bede;
    11'b00000000110: data <= 32'h3e74bbb2;
    11'b00000000111: data <= 32'hb034b831;
    11'b00000001000: data <= 32'hbd2cb633;
    11'b00000001001: data <= 32'hbaf13610;
    11'b00000001010: data <= 32'hb56e3df3;
    11'b00000001011: data <= 32'hbbe73d53;
    11'b00000001100: data <= 32'hbf6cb660;
    11'b00000001101: data <= 32'hbdc0be8a;
    11'b00000001110: data <= 32'hac88b92a;
    11'b00000001111: data <= 32'h3a5c3d7e;
    11'b00000010000: data <= 32'h3b063fc4;
    11'b00000010001: data <= 32'h3c123a9a;
    11'b00000010010: data <= 32'h3ce42ee5;
    11'b00000010011: data <= 32'h386f3a88;
    11'b00000010100: data <= 32'hba633db5;
    11'b00000010101: data <= 32'hbc60368a;
    11'b00000010110: data <= 32'h36eebd75;
    11'b00000010111: data <= 32'h4007c001;
    11'b00000011000: data <= 32'h3ea9bd3f;
    11'b00000011001: data <= 32'h2c43b8bd;
    11'b00000011010: data <= 32'hb809b57a;
    11'b00000011011: data <= 32'h355a2e5c;
    11'b00000011100: data <= 32'h38ab39a6;
    11'b00000011101: data <= 32'hbb273618;
    11'b00000011110: data <= 32'hc0fcbbfe;
    11'b00000011111: data <= 32'hc06ebefb;
    11'b00000100000: data <= 32'hb834b961;
    11'b00000100001: data <= 32'h38c43b67;
    11'b00000100010: data <= 32'h381d3c56;
    11'b00000100011: data <= 32'h3402312e;
    11'b00000100100: data <= 32'h34cd3402;
    11'b00000100101: data <= 32'ha6633f0f;
    11'b00000100110: data <= 32'hba834126;
    11'b00000100111: data <= 32'hbad93ca0;
    11'b00000101000: data <= 32'h3681bc40;
    11'b00000101001: data <= 32'h3e5abee6;
    11'b00000101010: data <= 32'h3d33b9d5;
    11'b00000101011: data <= 32'h36283064;
    11'b00000101100: data <= 32'h38e62b84;
    11'b00000101101: data <= 32'h3ec7ae31;
    11'b00000101110: data <= 32'h3df23119;
    11'b00000101111: data <= 32'hb9181a2d;
    11'b00000110000: data <= 32'hc0f4bbc0;
    11'b00000110001: data <= 32'hbff5be88;
    11'b00000110010: data <= 32'haf2cbc3d;
    11'b00000110011: data <= 32'h39ffb184;
    11'b00000110100: data <= 32'h2d37b45e;
    11'b00000110101: data <= 32'hb8a1b9d0;
    11'b00000110110: data <= 32'hb65130e1;
    11'b00000110111: data <= 32'hb433403b;
    11'b00000111000: data <= 32'hba8f41a0;
    11'b00000111001: data <= 32'hbcb03c83;
    11'b00000111010: data <= 32'hb7f3bbe1;
    11'b00000111011: data <= 32'h36fbbc91;
    11'b00000111100: data <= 32'h38ba3441;
    11'b00000111101: data <= 32'h38283c0c;
    11'b00000111110: data <= 32'h3d5b366a;
    11'b00000111111: data <= 32'h40cbb0b8;
    11'b00001000000: data <= 32'h3f5533f4;
    11'b00001000001: data <= 32'hb66338a1;
    11'b00001000010: data <= 32'hbf99b0a7;
    11'b00001000011: data <= 32'hbc18bcc9;
    11'b00001000100: data <= 32'h3a25bdc9;
    11'b00001000101: data <= 32'h3c33bccc;
    11'b00001000110: data <= 32'hb146bd49;
    11'b00001000111: data <= 32'hbabebd5c;
    11'b00001001000: data <= 32'hb354b03c;
    11'b00001001001: data <= 32'h328d3ed7;
    11'b00001001010: data <= 32'hb924402d;
    11'b00001001011: data <= 32'hbeff36e4;
    11'b00001001100: data <= 32'hbecbbc88;
    11'b00001001101: data <= 32'hba3cb92e;
    11'b00001001110: data <= 32'haf143b57;
    11'b00001001111: data <= 32'h354b3d13;
    11'b00001010000: data <= 32'h3cf133d2;
    11'b00001010001: data <= 32'h4022b1ab;
    11'b00001010010: data <= 32'h3dd93af0;
    11'b00001010011: data <= 32'hb5453f28;
    11'b00001010100: data <= 32'hbcc63c39;
    11'b00001010101: data <= 32'hac59b8b4;
    11'b00001010110: data <= 32'h3d76bdfa;
    11'b00001010111: data <= 32'h3c6fbdef;
    11'b00001011000: data <= 32'hb24dbdc3;
    11'b00001011001: data <= 32'hb60dbd5b;
    11'b00001011010: data <= 32'h3a68b6a9;
    11'b00001011011: data <= 32'h3cf83b1a;
    11'b00001011100: data <= 32'hb3b33bfe;
    11'b00001011101: data <= 32'hc03ab55d;
    11'b00001011110: data <= 32'hc0cabd14;
    11'b00001011111: data <= 32'hbd40b7ab;
    11'b00001100000: data <= 32'hb68b3a32;
    11'b00001100001: data <= 32'hacd038b6;
    11'b00001100010: data <= 32'h36ebb830;
    11'b00001100011: data <= 32'h3c25b59a;
    11'b00001100100: data <= 32'h39e33e12;
    11'b00001100101: data <= 32'hb63541af;
    11'b00001100110: data <= 32'hba5b3fa2;
    11'b00001100111: data <= 32'h3210b03a;
    11'b00001101000: data <= 32'h3c7dbc86;
    11'b00001101001: data <= 32'h3943baeb;
    11'b00001101010: data <= 32'hb215b91b;
    11'b00001101011: data <= 32'h36d7ba90;
    11'b00001101100: data <= 32'h401db881;
    11'b00001101101: data <= 32'h408b32c9;
    11'b00001101110: data <= 32'h331635bf;
    11'b00001101111: data <= 32'hbfddb7f5;
    11'b00001110000: data <= 32'hc041bc63;
    11'b00001110001: data <= 32'hbae7b88f;
    11'b00001110010: data <= 32'hb1b29d9b;
    11'b00001110011: data <= 32'hb773b93f;
    11'b00001110100: data <= 32'hb800be36;
    11'b00001110101: data <= 32'h2ea7b990;
    11'b00001110110: data <= 32'h34cc3eca;
    11'b00001110111: data <= 32'hb5d14212;
    11'b00001111000: data <= 32'hbab33f86;
    11'b00001111001: data <= 32'hb650ad50;
    11'b00001111010: data <= 32'h2e0bb88f;
    11'b00001111011: data <= 32'hb26832e4;
    11'b00001111100: data <= 32'hb55e3729;
    11'b00001111101: data <= 32'h3b91b47c;
    11'b00001111110: data <= 32'h416cb8ec;
    11'b00001111111: data <= 32'h41502b50;
    11'b00010000000: data <= 32'h37bd38f4;
    11'b00010000001: data <= 32'hbd8831fb;
    11'b00010000010: data <= 32'hbc5ab823;
    11'b00010000011: data <= 32'h325cb93b;
    11'b00010000100: data <= 32'h34f7ba5e;
    11'b00010000101: data <= 32'hb987be9e;
    11'b00010000110: data <= 32'hbbd2c07d;
    11'b00010000111: data <= 32'ha8efbc3e;
    11'b00010001000: data <= 32'h38e03d02;
    11'b00010001001: data <= 32'habac407e;
    11'b00010001010: data <= 32'hbc6a3c22;
    11'b00010001011: data <= 32'hbd58b664;
    11'b00010001100: data <= 32'hbc45aef3;
    11'b00010001101: data <= 32'hbc123c37;
    11'b00010001110: data <= 32'hb94c3c02;
    11'b00010001111: data <= 32'h3a26b42e;
    11'b00010010000: data <= 32'h40a7b9f7;
    11'b00010010001: data <= 32'h405a35e8;
    11'b00010010010: data <= 32'h36a13e35;
    11'b00010010011: data <= 32'hb9b03d4f;
    11'b00010010100: data <= 32'h28213385;
    11'b00010010101: data <= 32'h3c54b817;
    11'b00010010110: data <= 32'h387abbc2;
    11'b00010010111: data <= 32'hba5ebeeb;
    11'b00010011000: data <= 32'hba74c05c;
    11'b00010011001: data <= 32'h399ebcfc;
    11'b00010011010: data <= 32'h3e4b3750;
    11'b00010011011: data <= 32'h38023c0a;
    11'b00010011100: data <= 32'hbcf09cfe;
    11'b00010011101: data <= 32'hbf8eb9ea;
    11'b00010011110: data <= 32'hbe452eb3;
    11'b00010011111: data <= 32'hbd343cc0;
    11'b00010100000: data <= 32'hbc1538f4;
    11'b00010100001: data <= 32'ha591bb80;
    11'b00010100010: data <= 32'h3cadbc52;
    11'b00010100011: data <= 32'h3cc93a0f;
    11'b00010100100: data <= 32'h30b940dd;
    11'b00010100101: data <= 32'hb4ab404e;
    11'b00010100110: data <= 32'h386639d0;
    11'b00010100111: data <= 32'h3c94b070;
    11'b00010101000: data <= 32'h3319b578;
    11'b00010101001: data <= 32'hbb8bba8f;
    11'b00010101010: data <= 32'hb480bdc1;
    11'b00010101011: data <= 32'h3f0cbcc4;
    11'b00010101100: data <= 32'h4129b306;
    11'b00010101101: data <= 32'h3c2c3013;
    11'b00010101110: data <= 32'hbc15b7af;
    11'b00010101111: data <= 32'hbe56b9a3;
    11'b00010110000: data <= 32'hbc1f30df;
    11'b00010110001: data <= 32'hbb1b3994;
    11'b00010110010: data <= 32'hbceab68a;
    11'b00010110011: data <= 32'hbb8dbfc9;
    11'b00010110100: data <= 32'h220fbe2b;
    11'b00010110101: data <= 32'h37153a8b;
    11'b00010110110: data <= 32'h1e4d411f;
    11'b00010110111: data <= 32'hb304401d;
    11'b00010111000: data <= 32'h34273920;
    11'b00010111001: data <= 32'h35a93464;
    11'b00010111010: data <= 32'hb8e139cf;
    11'b00010111011: data <= 32'hbcee378b;
    11'b00010111100: data <= 32'h2cc4b8aa;
    11'b00010111101: data <= 32'h40a8bc36;
    11'b00010111110: data <= 32'h41d7b76a;
    11'b00010111111: data <= 32'h3ce32e06;
    11'b00011000000: data <= 32'hb856ab1d;
    11'b00011000001: data <= 32'hb867b155;
    11'b00011000010: data <= 32'h32f93356;
    11'b00011000011: data <= 32'hae292ed9;
    11'b00011000100: data <= 32'hbd00bd33;
    11'b00011000101: data <= 32'hbdf0c13a;
    11'b00011000110: data <= 32'hb6b2bf84;
    11'b00011000111: data <= 32'h378436e0;
    11'b00011001000: data <= 32'h33cf3f10;
    11'b00011001001: data <= 32'hb51f3c2e;
    11'b00011001010: data <= 32'hb7392978;
    11'b00011001011: data <= 32'hb971383b;
    11'b00011001100: data <= 32'hbdaf3e6f;
    11'b00011001101: data <= 32'hbe553d3a;
    11'b00011001110: data <= 32'hae1bb42c;
    11'b00011001111: data <= 32'h3fb4bc59;
    11'b00011010000: data <= 32'h4098b4f1;
    11'b00011010001: data <= 32'h3b393a32;
    11'b00011010010: data <= 32'hac503b75;
    11'b00011010011: data <= 32'h38d338bb;
    11'b00011010100: data <= 32'h3d80371a;
    11'b00011010101: data <= 32'h3790a67f;
    11'b00011010110: data <= 32'hbce9bd61;
    11'b00011010111: data <= 32'hbdd2c0e0;
    11'b00011011000: data <= 32'h2af7bf6c;
    11'b00011011001: data <= 32'h3d05b204;
    11'b00011011010: data <= 32'h3a7c3807;
    11'b00011011011: data <= 32'hb574b420;
    11'b00011011100: data <= 32'hbb55b905;
    11'b00011011101: data <= 32'hbc8d38b4;
    11'b00011011110: data <= 32'hbe853f78;
    11'b00011011111: data <= 32'hbf243cd0;
    11'b00011100000: data <= 32'hb9e8b9d9;
    11'b00011100001: data <= 32'h39f6bdab;
    11'b00011100010: data <= 32'h3c45ab14;
    11'b00011100011: data <= 32'h34d53e1a;
    11'b00011100100: data <= 32'h31a13ecf;
    11'b00011100101: data <= 32'h3cea3c29;
    11'b00011100110: data <= 32'h3ee839bd;
    11'b00011100111: data <= 32'h35ed37e3;
    11'b00011101000: data <= 32'hbd66b6a1;
    11'b00011101001: data <= 32'hbc50bddf;
    11'b00011101010: data <= 32'h3b9ebde6;
    11'b00011101011: data <= 32'h4061b967;
    11'b00011101100: data <= 32'h3d5ab797;
    11'b00011101101: data <= 32'hb16fbc22;
    11'b00011101110: data <= 32'hb96fbae3;
    11'b00011101111: data <= 32'hb8a238af;
    11'b00011110000: data <= 32'hbc113e1e;
    11'b00011110001: data <= 32'hbec335d7;
    11'b00011110010: data <= 32'hbddfbe99;
    11'b00011110011: data <= 32'hb7eabf89;
    11'b00011110100: data <= 32'h1dfd998d;
    11'b00011110101: data <= 32'hb06c3eb8;
    11'b00011110110: data <= 32'h31683e57;
    11'b00011110111: data <= 32'h3c5d3a55;
    11'b00011111000: data <= 32'h3c9c3aea;
    11'b00011111001: data <= 32'hb5943d83;
    11'b00011111010: data <= 32'hbea03b98;
    11'b00011111011: data <= 32'hba2db4dd;
    11'b00011111100: data <= 32'h3e05bc0c;
    11'b00011111101: data <= 32'h4103ba79;
    11'b00011111110: data <= 32'h3d92b93f;
    11'b00011111111: data <= 32'h2db5bad2;
    11'b00100000000: data <= 32'h3222b76f;
    11'b00100000001: data <= 32'h39dd3970;
    11'b00100000010: data <= 32'h2ccd3c17;
    11'b00100000011: data <= 32'hbd7cb7a4;
    11'b00100000100: data <= 32'hbf7cc096;
    11'b00100000101: data <= 32'hbc43c045;
    11'b00100000110: data <= 32'hb39db317;
    11'b00100000111: data <= 32'had163c15;
    11'b00100001000: data <= 32'h2ccd381e;
    11'b00100001001: data <= 32'h37d5adcc;
    11'b00100001010: data <= 32'h326b3a39;
    11'b00100001011: data <= 32'hbc894035;
    11'b00100001100: data <= 32'hbfd63fac;
    11'b00100001101: data <= 32'hba973502;
    11'b00100001110: data <= 32'h3cd8ba9b;
    11'b00100001111: data <= 32'h3f56b91f;
    11'b00100010000: data <= 32'h3a82aea3;
    11'b00100010001: data <= 32'h338124ad;
    11'b00100010010: data <= 32'h3cba341e;
    11'b00100010011: data <= 32'h40093b0a;
    11'b00100010100: data <= 32'h3baa3a95;
    11'b00100010101: data <= 32'hbc5bb8d5;
    11'b00100010110: data <= 32'hbf35c029;
    11'b00100010111: data <= 32'hb9dcbf8b;
    11'b00100011000: data <= 32'h364fb844;
    11'b00100011001: data <= 32'h36e6ad10;
    11'b00100011010: data <= 32'h2be2bb4b;
    11'b00100011011: data <= 32'h1c02bc5b;
    11'b00100011100: data <= 32'hb4f5385a;
    11'b00100011101: data <= 32'hbd474097;
    11'b00100011110: data <= 32'hbfe83fd8;
    11'b00100011111: data <= 32'hbcc6280c;
    11'b00100100000: data <= 32'h31f3bc47;
    11'b00100100001: data <= 32'h37ceb673;
    11'b00100100010: data <= 32'hafc03906;
    11'b00100100011: data <= 32'h31223a7c;
    11'b00100100100: data <= 32'h3ee03992;
    11'b00100100101: data <= 32'h410b3c0f;
    11'b00100100110: data <= 32'h3c533c70;
    11'b00100100111: data <= 32'hbc5d31cf;
    11'b00100101000: data <= 32'hbdc0bc05;
    11'b00100101001: data <= 32'h2f56bcb3;
    11'b00100101010: data <= 32'h3d48b981;
    11'b00100101011: data <= 32'h3ba4bb9b;
    11'b00100101100: data <= 32'h3074bf63;
    11'b00100101101: data <= 32'h2b36be55;
    11'b00100101110: data <= 32'h2f823617;
    11'b00100101111: data <= 32'hb8f33fd8;
    11'b00100110000: data <= 32'hbe483ccb;
    11'b00100110001: data <= 32'hbe5abac5;
    11'b00100110010: data <= 32'hbb7bbe20;
    11'b00100110011: data <= 32'hb9ecb4b5;
    11'b00100110100: data <= 32'hbadf3b5e;
    11'b00100110101: data <= 32'haa533a77;
    11'b00100110110: data <= 32'h3e473616;
    11'b00100110111: data <= 32'h40183b0e;
    11'b00100111000: data <= 32'h37003eae;
    11'b00100111001: data <= 32'hbd853dad;
    11'b00100111010: data <= 32'hbc69353d;
    11'b00100111011: data <= 32'h3a1db629;
    11'b00100111100: data <= 32'h3ef0b89f;
    11'b00100111101: data <= 32'h3bb7bc6a;
    11'b00100111110: data <= 32'h310cbf27;
    11'b00100111111: data <= 32'h3902bd37;
    11'b00101000000: data <= 32'h3d343706;
    11'b00101000001: data <= 32'h39193dc7;
    11'b00101000010: data <= 32'hbb3f34bd;
    11'b00101000011: data <= 32'hbedabe48;
    11'b00101000100: data <= 32'hbdd8bf08;
    11'b00101000101: data <= 32'hbc84b50c;
    11'b00101000110: data <= 32'hbbb53843;
    11'b00101000111: data <= 32'hb2b1b04e;
    11'b00101001000: data <= 32'h3bbfb93c;
    11'b00101001001: data <= 32'h3c473720;
    11'b00101001010: data <= 32'hb6864030;
    11'b00101001011: data <= 32'hbeb640a7;
    11'b00101001100: data <= 32'hbbfe3c71;
    11'b00101001101: data <= 32'h39a922b9;
    11'b00101001110: data <= 32'h3cbfb4df;
    11'b00101001111: data <= 32'h33f9b870;
    11'b00101010000: data <= 32'ha8e1bb6a;
    11'b00101010001: data <= 32'h3d37b862;
    11'b00101010010: data <= 32'h41073928;
    11'b00101010011: data <= 32'h3ecf3c84;
    11'b00101010100: data <= 32'hb5d8a877;
    11'b00101010101: data <= 32'hbdfbbdec;
    11'b00101010110: data <= 32'hbc81bd95;
    11'b00101010111: data <= 32'hb852b4e4;
    11'b00101011000: data <= 32'hb742b414;
    11'b00101011001: data <= 32'hb2eabdee;
    11'b00101011010: data <= 32'h366fbf63;
    11'b00101011011: data <= 32'h3635ad81;
    11'b00101011100: data <= 32'hb9ba4031;
    11'b00101011101: data <= 32'hbe7140b8;
    11'b00101011110: data <= 32'hbc4e3b3f;
    11'b00101011111: data <= 32'ha2bcb1f3;
    11'b00101100000: data <= 32'hace0abe3;
    11'b00101100001: data <= 32'hbb17335d;
    11'b00101100010: data <= 32'hb707196f;
    11'b00101100011: data <= 32'h3e772122;
    11'b00101100100: data <= 32'h420139cf;
    11'b00101100101: data <= 32'h3fbe3ca4;
    11'b00101100110: data <= 32'hb45c375c;
    11'b00101100111: data <= 32'hbc67b7ec;
    11'b00101101000: data <= 32'hb3ceb7c9;
    11'b00101101001: data <= 32'h37d0af55;
    11'b00101101010: data <= 32'h31b4bb03;
    11'b00101101011: data <= 32'hb141c0cb;
    11'b00101101100: data <= 32'h33a9c0f8;
    11'b00101101101: data <= 32'h3857b651;
    11'b00101101110: data <= 32'haf743ece;
    11'b00101101111: data <= 32'hbc143e4b;
    11'b00101110000: data <= 32'hbc79a90f;
    11'b00101110001: data <= 32'hbaebb9e4;
    11'b00101110010: data <= 32'hbd202af2;
    11'b00101110011: data <= 32'hbf333997;
    11'b00101110100: data <= 32'hbac63403;
    11'b00101110101: data <= 32'h3d7db22e;
    11'b00101110110: data <= 32'h410436f0;
    11'b00101110111: data <= 32'h3d0b3d81;
    11'b00101111000: data <= 32'hb8fe3da9;
    11'b00101111001: data <= 32'hba233a7a;
    11'b00101111010: data <= 32'h3863380e;
    11'b00101111011: data <= 32'h3c8433c2;
    11'b00101111100: data <= 32'h34f9bb33;
    11'b00101111101: data <= 32'hb461c0a8;
    11'b00101111110: data <= 32'h37c3c06e;
    11'b00101111111: data <= 32'h3dc2b4fa;
    11'b00110000000: data <= 32'h3c6a3cbb;
    11'b00110000001: data <= 32'hb0503870;
    11'b00110000010: data <= 32'hbba3bbbc;
    11'b00110000011: data <= 32'hbce9bc5f;
    11'b00110000100: data <= 32'hbead3021;
    11'b00110000101: data <= 32'hbfd738dc;
    11'b00110000110: data <= 32'hbc1bb688;
    11'b00110000111: data <= 32'h3a12bcb9;
    11'b00110001000: data <= 32'h3dc1b348;
    11'b00110001001: data <= 32'h33973dee;
    11'b00110001010: data <= 32'hbc364043;
    11'b00110001011: data <= 32'hb8c73e64;
    11'b00110001100: data <= 32'h3a113c08;
    11'b00110001101: data <= 32'h3ae138b7;
    11'b00110001110: data <= 32'hb57cb51c;
    11'b00110001111: data <= 32'hb97dbd95;
    11'b00110010000: data <= 32'h3aa0bd3f;
    11'b00110010001: data <= 32'h40e02582;
    11'b00110010010: data <= 32'h405b3a9b;
    11'b00110010011: data <= 32'h386da372;
    11'b00110010100: data <= 32'hb8d9bc99;
    11'b00110010101: data <= 32'hbaaeba7b;
    11'b00110010110: data <= 32'hbc1d3569;
    11'b00110010111: data <= 32'hbd5d3104;
    11'b00110011000: data <= 32'hbb61be1a;
    11'b00110011001: data <= 32'h3168c0c5;
    11'b00110011010: data <= 32'h385fbb8b;
    11'b00110011011: data <= 32'hb5673d33;
    11'b00110011100: data <= 32'hbc584028;
    11'b00110011101: data <= 32'hb7fe3d72;
    11'b00110011110: data <= 32'h35eb39f8;
    11'b00110011111: data <= 32'hb12b3a03;
    11'b00110100000: data <= 32'hbdf437b1;
    11'b00110100001: data <= 32'hbd32b489;
    11'b00110100010: data <= 32'h3b4cb7f2;
    11'b00110100011: data <= 32'h41a0332c;
    11'b00110100100: data <= 32'h40cb39b1;
    11'b00110100101: data <= 32'h39133119;
    11'b00110100110: data <= 32'hb405b6aa;
    11'b00110100111: data <= 32'h2c1d2e75;
    11'b00110101000: data <= 32'h31023a11;
    11'b00110101001: data <= 32'hb782b264;
    11'b00110101010: data <= 32'hb9e0c09c;
    11'b00110101011: data <= 32'haedcc20e;
    11'b00110101100: data <= 32'h3655bd2b;
    11'b00110101101: data <= 32'h950f3b28;
    11'b00110101110: data <= 32'hb8143d0d;
    11'b00110101111: data <= 32'hb4e9348d;
    11'b00110110000: data <= 32'hb215a4c5;
    11'b00110110001: data <= 32'hbcdb39d1;
    11'b00110110010: data <= 32'hc0da3c23;
    11'b00110110011: data <= 32'hbf323402;
    11'b00110110100: data <= 32'h38dbb6d3;
    11'b00110110101: data <= 32'h408ea7ac;
    11'b00110110110: data <= 32'h3e77399b;
    11'b00110110111: data <= 32'h2e833a71;
    11'b00110111000: data <= 32'haa6239bf;
    11'b00110111001: data <= 32'h3b5e3c88;
    11'b00110111010: data <= 32'h3c403d07;
    11'b00110111011: data <= 32'hab47af35;
    11'b00110111100: data <= 32'hba39c05c;
    11'b00110111101: data <= 32'hac78c15c;
    11'b00110111110: data <= 32'h3bccbc47;
    11'b00110111111: data <= 32'h3c1f37d4;
    11'b00111000000: data <= 32'h36ba3224;
    11'b00111000001: data <= 32'h2921bb1c;
    11'b00111000010: data <= 32'hb652b942;
    11'b00111000011: data <= 32'hbe2039ac;
    11'b00111000100: data <= 32'hc1143c81;
    11'b00111000101: data <= 32'hbf8fadb5;
    11'b00111000110: data <= 32'h2cf5bcd3;
    11'b00111000111: data <= 32'h3ca4b9da;
    11'b00111001000: data <= 32'h35de38c2;
    11'b00111001001: data <= 32'hb8d83d48;
    11'b00111001010: data <= 32'h1e8a3db1;
    11'b00111001011: data <= 32'h3d293e7d;
    11'b00111001100: data <= 32'h3c703e4a;
    11'b00111001101: data <= 32'hb7bd36bf;
    11'b00111001110: data <= 32'hbcddbccf;
    11'b00111001111: data <= 32'h2a00be4a;
    11'b00111010000: data <= 32'h3ef4b786;
    11'b00111010001: data <= 32'h40033427;
    11'b00111010010: data <= 32'h3c81b81d;
    11'b00111010011: data <= 32'h36a8bd89;
    11'b00111010100: data <= 32'h9cfab8f7;
    11'b00111010101: data <= 32'hbac53b61;
    11'b00111010110: data <= 32'hbefd3b3c;
    11'b00111010111: data <= 32'hbe2bbb96;
    11'b00111011000: data <= 32'hb614c098;
    11'b00111011001: data <= 32'h30cabdf4;
    11'b00111011010: data <= 32'hb8213544;
    11'b00111011011: data <= 32'hbb3d3ce4;
    11'b00111011100: data <= 32'h2d483c8e;
    11'b00111011101: data <= 32'h3c7f3ce5;
    11'b00111011110: data <= 32'h35d23e1c;
    11'b00111011111: data <= 32'hbdff3c62;
    11'b00111100000: data <= 32'hbf8b2264;
    11'b00111100001: data <= 32'h1498b74e;
    11'b00111100010: data <= 32'h400d247a;
    11'b00111100011: data <= 32'h405a3243;
    11'b00111100100: data <= 32'h3c72b86b;
    11'b00111100101: data <= 32'h38e6bb89;
    11'b00111100110: data <= 32'h3a4e3089;
    11'b00111100111: data <= 32'h36dc3d9f;
    11'b00111101000: data <= 32'hb8b439b6;
    11'b00111101001: data <= 32'hbc3bbe69;
    11'b00111101010: data <= 32'hb8a0c1c6;
    11'b00111101011: data <= 32'hb25fbf22;
    11'b00111101100: data <= 32'hb7c52710;
    11'b00111101101: data <= 32'hb80637c8;
    11'b00111101110: data <= 32'h3555a4cf;
    11'b00111101111: data <= 32'h3a0d322a;
    11'b00111110000: data <= 32'hb83d3cd4;
    11'b00111110001: data <= 32'hc0c33e33;
    11'b00111110010: data <= 32'hc0bd39d4;
    11'b00111110011: data <= 32'hb41cac55;
    11'b00111110100: data <= 32'h3e23a80f;
    11'b00111110101: data <= 32'h3d483089;
    11'b00111110110: data <= 32'h3574af69;
    11'b00111110111: data <= 32'h38431cf1;
    11'b00111111000: data <= 32'h3e233c73;
    11'b00111111001: data <= 32'h3e013fb3;
    11'b00111111010: data <= 32'h30dd3a78;
    11'b00111111011: data <= 32'hbae9bdf4;
    11'b00111111100: data <= 32'hb879c0f2;
    11'b00111111101: data <= 32'h3132bd6d;
    11'b00111111110: data <= 32'h3544afea;
    11'b00111111111: data <= 32'h35adb797;
    11'b01000000000: data <= 32'h39d6bd63;
    11'b01000000001: data <= 32'h38e2ba38;
    11'b01000000010: data <= 32'hba9a3b64;
    11'b01000000011: data <= 32'hc0e13e87;
    11'b01000000100: data <= 32'hc09938db;
    11'b01000000101: data <= 32'hb88eb8d3;
    11'b01000000110: data <= 32'h3826b91f;
    11'b01000000111: data <= 32'hacbca7ca;
    11'b01000001000: data <= 32'hb99134bb;
    11'b01000001001: data <= 32'h34dc393d;
    11'b01000001010: data <= 32'h3f783e3d;
    11'b01000001011: data <= 32'h3f0e4040;
    11'b01000001100: data <= 32'h9c2d3caf;
    11'b01000001101: data <= 32'hbcb9b8c6;
    11'b01000001110: data <= 32'hb818bced;
    11'b01000001111: data <= 32'h3a4bb6fd;
    11'b01000010000: data <= 32'h3ce1ab5a;
    11'b01000010001: data <= 32'h3c1dbc7f;
    11'b01000010010: data <= 32'h3c2bc01b;
    11'b01000010011: data <= 32'h3b0cbc24;
    11'b01000010100: data <= 32'hb2b13bde;
    11'b01000010101: data <= 32'hbe1f3de2;
    11'b01000010110: data <= 32'hbe9aad9a;
    11'b01000010111: data <= 32'hb9d8be4e;
    11'b01000011000: data <= 32'hb6c0bd78;
    11'b01000011001: data <= 32'hbcaab46f;
    11'b01000011010: data <= 32'hbd423439;
    11'b01000011011: data <= 32'h322036b4;
    11'b01000011100: data <= 32'h3efd3c42;
    11'b01000011101: data <= 32'h3ccd3f40;
    11'b01000011110: data <= 32'hbafc3e40;
    11'b01000011111: data <= 32'hbf433852;
    11'b01000100000: data <= 32'hb8972dc6;
    11'b01000100001: data <= 32'h3c5b3642;
    11'b01000100010: data <= 32'h3da62e83;
    11'b01000100011: data <= 32'h3b81bcc3;
    11'b01000100100: data <= 32'h3c0dbf3c;
    11'b01000100101: data <= 32'h3dabb73a;
    11'b01000100110: data <= 32'h3be33dad;
    11'b01000100111: data <= 32'hb1823d49;
    11'b01000101000: data <= 32'hba80b9b5;
    11'b01000101001: data <= 32'hb965c056;
    11'b01000101010: data <= 32'hba3cbe6e;
    11'b01000101011: data <= 32'hbd64b672;
    11'b01000101100: data <= 32'hbc81b40e;
    11'b01000101101: data <= 32'h35f9b94d;
    11'b01000101110: data <= 32'h3dbdb0e7;
    11'b01000101111: data <= 32'h35f33c8c;
    11'b01000110000: data <= 32'hbeef3ef5;
    11'b01000110001: data <= 32'hc0873cfc;
    11'b01000110010: data <= 32'hb9a539a1;
    11'b01000110011: data <= 32'h3a3238c1;
    11'b01000110100: data <= 32'h390030b5;
    11'b01000110101: data <= 32'h9431ba85;
    11'b01000110110: data <= 32'h38babbaf;
    11'b01000110111: data <= 32'h3f81379e;
    11'b01000111000: data <= 32'h40113fac;
    11'b01000111001: data <= 32'h3a6a3d58;
    11'b01000111010: data <= 32'hb53eb9dc;
    11'b01000111011: data <= 32'hb827bf3f;
    11'b01000111100: data <= 32'hb79ebc24;
    11'b01000111101: data <= 32'hb94bb38e;
    11'b01000111110: data <= 32'hb570bb73;
    11'b01000111111: data <= 32'h3a10bfd3;
    11'b01001000000: data <= 32'h3d01bd73;
    11'b01001000001: data <= 32'ha403383d;
    11'b01001000010: data <= 32'hbf5f3e95;
    11'b01001000011: data <= 32'hc0263cb2;
    11'b01001000100: data <= 32'hb9e03538;
    11'b01001000101: data <= 32'h26d22dfb;
    11'b01001000110: data <= 32'hb9d9a0f5;
    11'b01001000111: data <= 32'hbd1db66b;
    11'b01001001000: data <= 32'h2322b421;
    11'b01001001001: data <= 32'h3fff3bba;
    11'b01001001010: data <= 32'h40aa4010;
    11'b01001001011: data <= 32'h3aa43dd4;
    11'b01001001100: data <= 32'hb7ecad91;
    11'b01001001101: data <= 32'hb709b8e5;
    11'b01001001110: data <= 32'h30052fbe;
    11'b01001001111: data <= 32'h33be3224;
    11'b01001010000: data <= 32'h35dcbd62;
    11'b01001010001: data <= 32'h3c0ec161;
    11'b01001010010: data <= 32'h3d4fbf52;
    11'b01001010011: data <= 32'h361a3655;
    11'b01001010100: data <= 32'hbbd33db4;
    11'b01001010101: data <= 32'hbcd03821;
    11'b01001010110: data <= 32'hb841b8fd;
    11'b01001010111: data <= 32'hb94cb932;
    11'b01001011000: data <= 32'hbf61b33e;
    11'b01001011001: data <= 32'hc042b49a;
    11'b01001011010: data <= 32'hb564b4e5;
    11'b01001011011: data <= 32'h3f273829;
    11'b01001011100: data <= 32'h3f403e13;
    11'b01001011101: data <= 32'h25193dfb;
    11'b01001011110: data <= 32'hbc7b3a53;
    11'b01001011111: data <= 32'hb7cd39d0;
    11'b01001100000: data <= 32'h383a3cd0;
    11'b01001100001: data <= 32'h38b7390f;
    11'b01001100010: data <= 32'h354cbd27;
    11'b01001100011: data <= 32'h3a8bc0fc;
    11'b01001100100: data <= 32'h3e24bd5b;
    11'b01001100101: data <= 32'h3d453a53;
    11'b01001100110: data <= 32'h36413d10;
    11'b01001100111: data <= 32'hae1eb18d;
    11'b01001101000: data <= 32'hb104bd58;
    11'b01001101001: data <= 32'hbaebbb96;
    11'b01001101010: data <= 32'hc027b311;
    11'b01001101011: data <= 32'hc025b81a;
    11'b01001101100: data <= 32'hb37dbc8d;
    11'b01001101101: data <= 32'h3dd7b998;
    11'b01001101110: data <= 32'h3b98388e;
    11'b01001101111: data <= 32'hbb733d4d;
    11'b01001110000: data <= 32'hbe843d40;
    11'b01001110001: data <= 32'hb82f3d94;
    11'b01001110010: data <= 32'h37713e4f;
    11'b01001110011: data <= 32'h28ac3a6b;
    11'b01001110100: data <= 32'hb8ccbb10;
    11'b01001110101: data <= 32'h302ebe87;
    11'b01001110110: data <= 32'h3e88b5a7;
    11'b01001110111: data <= 32'h40513d60;
    11'b01001111000: data <= 32'h3daf3cdd;
    11'b01001111001: data <= 32'h38cdb674;
    11'b01001111010: data <= 32'h3195bcc9;
    11'b01001111011: data <= 32'hb812b656;
    11'b01001111100: data <= 32'hbd98321d;
    11'b01001111101: data <= 32'hbd0ebaa6;
    11'b01001111110: data <= 32'h3225c06c;
    11'b01001111111: data <= 32'h3cf1bfdc;
    11'b01010000000: data <= 32'h3639b486;
    11'b01010000001: data <= 32'hbcf43c05;
    11'b01010000010: data <= 32'hbde43ca4;
    11'b01010000011: data <= 32'hb5573c2c;
    11'b01010000100: data <= 32'h2c0f3c62;
    11'b01010000101: data <= 32'hbc603904;
    11'b01010000110: data <= 32'hbfbab71b;
    11'b01010000111: data <= 32'hb9bcba57;
    11'b01010001000: data <= 32'h3df13513;
    11'b01010001001: data <= 32'h40b33e08;
    11'b01010001010: data <= 32'h3df73c9b;
    11'b01010001011: data <= 32'h37fdad4b;
    11'b01010001100: data <= 32'h3456b31e;
    11'b01010001101: data <= 32'h2f2b3a7c;
    11'b01010001110: data <= 32'hb6433b3c;
    11'b01010001111: data <= 32'hb65fbb86;
    11'b01010010000: data <= 32'h381cc1a0;
    11'b01010010001: data <= 32'h3ca7c0fa;
    11'b01010010010: data <= 32'h37cdb842;
    11'b01010010011: data <= 32'hb8ca39c9;
    11'b01010010100: data <= 32'hb87d37a5;
    11'b01010010101: data <= 32'h310e2537;
    11'b01010010110: data <= 32'hb4c23318;
    11'b01010010111: data <= 32'hc01d3565;
    11'b01010011000: data <= 32'hc1b5b300;
    11'b01010011001: data <= 32'hbcecb894;
    11'b01010011010: data <= 32'h3ca72e22;
    11'b01010011011: data <= 32'h3f2a3bc7;
    11'b01010011100: data <= 32'h39143b45;
    11'b01010011101: data <= 32'hb32a3743;
    11'b01010011110: data <= 32'h30eb3b9d;
    11'b01010011111: data <= 32'h38c43fe8;
    11'b01010100000: data <= 32'h32273e36;
    11'b01010100001: data <= 32'hb2c3b9c8;
    11'b01010100010: data <= 32'h351ac11e;
    11'b01010100011: data <= 32'h3c71bfe9;
    11'b01010100100: data <= 32'h3c52ad27;
    11'b01010100101: data <= 32'h38c038ef;
    11'b01010100110: data <= 32'h391eb45b;
    11'b01010100111: data <= 32'h3a3fbb2d;
    11'b01010101000: data <= 32'hb4b3b4af;
    11'b01010101001: data <= 32'hc06f350d;
    11'b01010101010: data <= 32'hc19bb2d0;
    11'b01010101011: data <= 32'hbc77bc45;
    11'b01010101100: data <= 32'h3ae5bb7e;
    11'b01010101101: data <= 32'h3b06ac7b;
    11'b01010101110: data <= 32'hb7e03760;
    11'b01010101111: data <= 32'hbb7e39d6;
    11'b01010110000: data <= 32'h2c6d3e24;
    11'b01010110001: data <= 32'h39d640c6;
    11'b01010110010: data <= 32'ha9083f0f;
    11'b01010110011: data <= 32'hbb8eb4f2;
    11'b01010110100: data <= 32'hb739be9d;
    11'b01010110101: data <= 32'h3b53babe;
    11'b01010110110: data <= 32'h3e92394b;
    11'b01010110111: data <= 32'h3e1b390b;
    11'b01010111000: data <= 32'h3d9cb956;
    11'b01010111001: data <= 32'h3cd8bc3d;
    11'b01010111010: data <= 32'h2f1e2ab0;
    11'b01010111011: data <= 32'hbdfc3a57;
    11'b01010111100: data <= 32'hbf81b39a;
    11'b01010111101: data <= 32'hb834bf5c;
    11'b01010111110: data <= 32'h39abc02e;
    11'b01010111111: data <= 32'h31c8bc0e;
    11'b01011000000: data <= 32'hbc57a330;
    11'b01011000001: data <= 32'hbbfa37b5;
    11'b01011000010: data <= 32'h34cb3c8c;
    11'b01011000011: data <= 32'h38e23f4c;
    11'b01011000100: data <= 32'hbadc3dd5;
    11'b01011000101: data <= 32'hc04e2bca;
    11'b01011000110: data <= 32'hbda1b99a;
    11'b01011000111: data <= 32'h38822e0c;
    11'b01011001000: data <= 32'h3ec43c34;
    11'b01011001001: data <= 32'h3e2e386b;
    11'b01011001010: data <= 32'h3d08b8e2;
    11'b01011001011: data <= 32'h3ce3b674;
    11'b01011001100: data <= 32'h396d3c7e;
    11'b01011001101: data <= 32'hb64a3e7e;
    11'b01011001110: data <= 32'hba1caec7;
    11'b01011001111: data <= 32'h26e7c084;
    11'b01011010000: data <= 32'h3933c11e;
    11'b01011010001: data <= 32'h28c7bd0b;
    11'b01011010010: data <= 32'hba1cb43e;
    11'b01011010011: data <= 32'hb388b189;
    11'b01011010100: data <= 32'h3b432834;
    11'b01011010101: data <= 32'h382139d3;
    11'b01011010110: data <= 32'hbe6c3b85;
    11'b01011010111: data <= 32'hc20733ee;
    11'b01011011000: data <= 32'hbfd4b434;
    11'b01011011001: data <= 32'h32db3224;
    11'b01011011010: data <= 32'h3c81397a;
    11'b01011011011: data <= 32'h38ef3281;
    11'b01011011100: data <= 32'h3585b5ad;
    11'b01011011101: data <= 32'h3b203840;
    11'b01011011110: data <= 32'h3c6d4073;
    11'b01011011111: data <= 32'h361f40b0;
    11'b01011100000: data <= 32'hb42b3246;
    11'b01011100001: data <= 32'h2657bfd9;
    11'b01011100010: data <= 32'h3819bfed;
    11'b01011100011: data <= 32'h3583b93f;
    11'b01011100100: data <= 32'h3165b1f3;
    11'b01011100101: data <= 32'h3b2bbae7;
    11'b01011100110: data <= 32'h3e89bc37;
    11'b01011100111: data <= 32'h3941ae25;
    11'b01011101000: data <= 32'hbebf39a1;
    11'b01011101001: data <= 32'hc1cf34f5;
    11'b01011101010: data <= 32'hbeeeb7a6;
    11'b01011101011: data <= 32'h2bb8b87d;
    11'b01011101100: data <= 32'h3442b46d;
    11'b01011101101: data <= 32'hb94bb5e8;
    11'b01011101110: data <= 32'hb953b433;
    11'b01011101111: data <= 32'h389a3c01;
    11'b01011110000: data <= 32'h3d11412d;
    11'b01011110001: data <= 32'h36b340fb;
    11'b01011110010: data <= 32'hb9973812;
    11'b01011110011: data <= 32'hb929bc60;
    11'b01011110100: data <= 32'h31e1b9af;
    11'b01011110101: data <= 32'h397d35e4;
    11'b01011110110: data <= 32'h3ba82c39;
    11'b01011110111: data <= 32'h3e7dbd08;
    11'b01011111000: data <= 32'h4019bde1;
    11'b01011111001: data <= 32'h3c0eab75;
    11'b01011111010: data <= 32'hbbdc3c38;
    11'b01011111011: data <= 32'hbf6e369f;
    11'b01011111100: data <= 32'hbb0dbc03;
    11'b01011111101: data <= 32'h3090be2c;
    11'b01011111110: data <= 32'hb69fbcc3;
    11'b01011111111: data <= 32'hbdf9bb06;
    11'b01100000000: data <= 32'hbc2db827;
    11'b01100000001: data <= 32'h393a38c8;
    11'b01100000010: data <= 32'h3d0b3fb0;
    11'b01100000011: data <= 32'hb06e3fd3;
    11'b01100000100: data <= 32'hbed63941;
    11'b01100000101: data <= 32'hbe49b167;
    11'b01100000110: data <= 32'hb3c93741;
    11'b01100000111: data <= 32'h395d3c56;
    11'b01100001000: data <= 32'h3b8d315f;
    11'b01100001001: data <= 32'h3d95bd2e;
    11'b01100001010: data <= 32'h3f81bc52;
    11'b01100001011: data <= 32'h3d8a3a52;
    11'b01100001100: data <= 32'h2da73f64;
    11'b01100001101: data <= 32'hb8413934;
    11'b01100001110: data <= 32'h1ab3bd3b;
    11'b01100001111: data <= 32'h34a5bfce;
    11'b01100010000: data <= 32'hb905bd83;
    11'b01100010001: data <= 32'hbdc4bbfb;
    11'b01100010010: data <= 32'hb839bc11;
    11'b01100010011: data <= 32'h3cd6b7a4;
    11'b01100010100: data <= 32'h3d283909;
    11'b01100010101: data <= 32'hb9dc3c6f;
    11'b01100010110: data <= 32'hc0f938ef;
    11'b01100010111: data <= 32'hc0293512;
    11'b01100011000: data <= 32'hb8203a95;
    11'b01100011001: data <= 32'h32dd3be9;
    11'b01100011010: data <= 32'h2882aedf;
    11'b01100011011: data <= 32'h34e8bcae;
    11'b01100011100: data <= 32'h3cecb54c;
    11'b01100011101: data <= 32'h3e4e3f26;
    11'b01100011110: data <= 32'h3b234117;
    11'b01100011111: data <= 32'h33cb3b6b;
    11'b01100100000: data <= 32'h34cabc48;
    11'b01100100001: data <= 32'h3415bd86;
    11'b01100100010: data <= 32'hb72fb8f6;
    11'b01100100011: data <= 32'hb9c4b90e;
    11'b01100100100: data <= 32'h379ebde5;
    11'b01100100101: data <= 32'h3fb3be4f;
    11'b01100100110: data <= 32'h3dcfb76a;
    11'b01100100111: data <= 32'hba973866;
    11'b01100101000: data <= 32'hc0bd3856;
    11'b01100101001: data <= 32'hbeeb330c;
    11'b01100101010: data <= 32'hb6c034da;
    11'b01100101011: data <= 32'hb6e131cf;
    11'b01100101100: data <= 32'hbcfeb964;
    11'b01100101101: data <= 32'hbbbbbc8e;
    11'b01100101110: data <= 32'h38992eb3;
    11'b01100101111: data <= 32'h3e444043;
    11'b01100110000: data <= 32'h3c1f4131;
    11'b01100110001: data <= 32'h2b543c27;
    11'b01100110010: data <= 32'hb1ecb641;
    11'b01100110011: data <= 32'habb1aed6;
    11'b01100110100: data <= 32'hb2693940;
    11'b01100110101: data <= 32'ha043a813;
    11'b01100110110: data <= 32'h3cafbeb1;
    11'b01100110111: data <= 32'h408dc028;
    11'b01100111000: data <= 32'h3ea3b98a;
    11'b01100111001: data <= 32'hb4653970;
    11'b01100111010: data <= 32'hbd4638e9;
    11'b01100111011: data <= 32'hb922b233;
    11'b01100111100: data <= 32'h1deab884;
    11'b01100111101: data <= 32'hbb30b97f;
    11'b01100111110: data <= 32'hc04dbc99;
    11'b01100111111: data <= 32'hbe7fbd34;
    11'b01101000000: data <= 32'h3655b1cb;
    11'b01101000001: data <= 32'h3e003dd9;
    11'b01101000010: data <= 32'h38be3f65;
    11'b01101000011: data <= 32'hba713ad9;
    11'b01101000100: data <= 32'hbc2f3514;
    11'b01101000101: data <= 32'hb7a43c7a;
    11'b01101000110: data <= 32'hb18e3ea6;
    11'b01101000111: data <= 32'h2b4135c6;
    11'b01101001000: data <= 32'h3b8dbe79;
    11'b01101001001: data <= 32'h3fb0bf3b;
    11'b01101001010: data <= 32'h3ee8a54e;
    11'b01101001011: data <= 32'h38a93d87;
    11'b01101001100: data <= 32'h2c023ad2;
    11'b01101001101: data <= 32'h3854b7eb;
    11'b01101001110: data <= 32'h3797bc0b;
    11'b01101001111: data <= 32'hbbedbafe;
    11'b01101010000: data <= 32'hc06fbc81;
    11'b01101010001: data <= 32'hbd40be24;
    11'b01101010010: data <= 32'h3aa5bc39;
    11'b01101010011: data <= 32'h3e202fbb;
    11'b01101010100: data <= 32'h28ca399c;
    11'b01101010101: data <= 32'hbe54378e;
    11'b01101010110: data <= 32'hbe37393c;
    11'b01101010111: data <= 32'hb92b3e69;
    11'b01101011000: data <= 32'hb6a33f35;
    11'b01101011001: data <= 32'hb96133c7;
    11'b01101011010: data <= 32'hb1ebbdf1;
    11'b01101011011: data <= 32'h3be5bc7e;
    11'b01101011100: data <= 32'h3e403b89;
    11'b01101011101: data <= 32'h3cdc4025;
    11'b01101011110: data <= 32'h3b973c3f;
    11'b01101011111: data <= 32'h3c68b6ba;
    11'b01101100000: data <= 32'h391bb8bf;
    11'b01101100001: data <= 32'hba4dad81;
    11'b01101100010: data <= 32'hbe52b7e0;
    11'b01101100011: data <= 32'hb605be8f;
    11'b01101100100: data <= 32'h3e1fbfe1;
    11'b01101100101: data <= 32'h3ea0bc51;
    11'b01101100110: data <= 32'hb16ab0cc;
    11'b01101100111: data <= 32'hbe5d30ef;
    11'b01101101000: data <= 32'hbcba3812;
    11'b01101101001: data <= 32'hb5093cbb;
    11'b01101101010: data <= 32'hb9ce3c63;
    11'b01101101011: data <= 32'hbf11b4a8;
    11'b01101101100: data <= 32'hbe3dbdc4;
    11'b01101101101: data <= 32'h24cfb8ee;
    11'b01101101110: data <= 32'h3d133d89;
    11'b01101101111: data <= 32'h3d1c403a;
    11'b01101110000: data <= 32'h3aff3bc7;
    11'b01101110001: data <= 32'h3a14a9c3;
    11'b01101110010: data <= 32'h361b37f1;
    11'b01101110011: data <= 32'hb84d3d25;
    11'b01101110100: data <= 32'hbaad36e4;
    11'b01101110101: data <= 32'h363ebe18;
    11'b01101110110: data <= 32'h3f8ac0bc;
    11'b01101110111: data <= 32'h3ed0bdb7;
    11'b01101111000: data <= 32'h2f2ab289;
    11'b01101111001: data <= 32'hb9b83025;
    11'b01101111010: data <= 32'h9e172e20;
    11'b01101111011: data <= 32'h36f83514;
    11'b01101111100: data <= 32'hbade31ef;
    11'b01101111101: data <= 32'hc117ba3f;
    11'b01101111110: data <= 32'hc0b1bdf0;
    11'b01101111111: data <= 32'hb62eb963;
    11'b01110000000: data <= 32'h3c403b07;
    11'b01110000001: data <= 32'h3aa43d2a;
    11'b01110000010: data <= 32'h299337a3;
    11'b01110000011: data <= 32'haf13351e;
    11'b01110000100: data <= 32'haa973e57;
    11'b01110000101: data <= 32'hb6e940db;
    11'b01110000110: data <= 32'hb8aa3c59;
    11'b01110000111: data <= 32'h3510bd21;
    11'b01110001000: data <= 32'h3de6c024;
    11'b01110001001: data <= 32'h3decba82;
    11'b01110001010: data <= 32'h39093784;
    11'b01110001011: data <= 32'h382c35fd;
    11'b01110001100: data <= 32'h3d47b40f;
    11'b01110001101: data <= 32'h3cceb461;
    11'b01110001110: data <= 32'hb9c7b086;
    11'b01110001111: data <= 32'hc122b9cb;
    11'b01110010000: data <= 32'hc039bdd9;
    11'b01110010001: data <= 32'ha55dbce3;
    11'b01110010010: data <= 32'h3c50b500;
    11'b01110010011: data <= 32'h33e00cc1;
    11'b01110010100: data <= 32'hbab8b35a;
    11'b01110010101: data <= 32'hb9f03642;
    11'b01110010110: data <= 32'hb2bf4004;
    11'b01110010111: data <= 32'hb7514156;
    11'b01110011000: data <= 32'hbc0a3c56;
    11'b01110011001: data <= 32'hb945bc6b;
    11'b01110011010: data <= 32'h3670bd78;
    11'b01110011011: data <= 32'h3bd53314;
    11'b01110011100: data <= 32'h3bba3d0e;
    11'b01110011101: data <= 32'h3d5638be;
    11'b01110011110: data <= 32'h4003b5a5;
    11'b01110011111: data <= 32'h3e1eb021;
    11'b01110100000: data <= 32'hb6ff37db;
    11'b01110100001: data <= 32'hbfa627c3;
    11'b01110100010: data <= 32'hbc8bbceb;
    11'b01110100011: data <= 32'h3a0fbf48;
    11'b01110100100: data <= 32'h3ce4bdb5;
    11'b01110100101: data <= 32'hae26bbff;
    11'b01110100110: data <= 32'hbc5cba1b;
    11'b01110100111: data <= 32'hb8352fcf;
    11'b01110101000: data <= 32'h33023e47;
    11'b01110101001: data <= 32'hb7223fd3;
    11'b01110101010: data <= 32'hbf1f3803;
    11'b01110101011: data <= 32'hbfbfbc53;
    11'b01110101100: data <= 32'hb9d9ba0c;
    11'b01110101101: data <= 32'h36c33aff;
    11'b01110101110: data <= 32'h3ae23dd7;
    11'b01110101111: data <= 32'h3cf136e3;
    11'b01110110000: data <= 32'h3ec3b464;
    11'b01110110001: data <= 32'h3d0f3920;
    11'b01110110010: data <= 32'hb2683f08;
    11'b01110110011: data <= 32'hbc5b3c81;
    11'b01110110100: data <= 32'hb1f9ba81;
    11'b01110110101: data <= 32'h3d10c005;
    11'b01110110110: data <= 32'h3ce6befb;
    11'b01110110111: data <= 32'had2dbc78;
    11'b01110111000: data <= 32'hb82ebaa2;
    11'b01110111001: data <= 32'h384db4c7;
    11'b01110111010: data <= 32'h3c923929;
    11'b01110111011: data <= 32'hb4143b23;
    11'b01110111100: data <= 32'hc0a2b05a;
    11'b01110111101: data <= 32'hc15ebc6d;
    11'b01110111110: data <= 32'hbcf2b8a6;
    11'b01110111111: data <= 32'h2f9f3951;
    11'b01111000000: data <= 32'h36013a12;
    11'b01111000001: data <= 32'h35c0b351;
    11'b01111000010: data <= 32'h399eb3ce;
    11'b01111000011: data <= 32'h39933ddc;
    11'b01111000100: data <= 32'hae5241b6;
    11'b01111000101: data <= 32'hb91e3faa;
    11'b01111000110: data <= 32'h2550b6b7;
    11'b01111000111: data <= 32'h3beabe8d;
    11'b01111001000: data <= 32'h3adabc5f;
    11'b01111001001: data <= 32'h2e90b5d1;
    11'b01111001010: data <= 32'h36f3b799;
    11'b01111001011: data <= 32'h3f44b90d;
    11'b01111001100: data <= 32'h4024af12;
    11'b01111001101: data <= 32'h2d7534d1;
    11'b01111001110: data <= 32'hc073b354;
    11'b01111001111: data <= 32'hc0d7bbb9;
    11'b01111010000: data <= 32'hbaa6ba73;
    11'b01111010001: data <= 32'h32a7b396;
    11'b01111010010: data <= 32'hb22bb7ae;
    11'b01111010011: data <= 32'hb948bc7b;
    11'b01111010100: data <= 32'hb18cb6be;
    11'b01111010101: data <= 32'h36043ef7;
    11'b01111010110: data <= 32'ha8ce4224;
    11'b01111010111: data <= 32'hba1b3fab;
    11'b01111011000: data <= 32'hb947b452;
    11'b01111011001: data <= 32'ha4f5bb80;
    11'b01111011010: data <= 32'h310b2b34;
    11'b01111011011: data <= 32'h30ef3934;
    11'b01111011100: data <= 32'h3c47adb9;
    11'b01111011101: data <= 32'h40f8ba48;
    11'b01111011110: data <= 32'h40e5b3c3;
    11'b01111011111: data <= 32'h364c3918;
    11'b01111100000: data <= 32'hbe383721;
    11'b01111100001: data <= 32'hbd62b84c;
    11'b01111100010: data <= 32'h3076bc61;
    11'b01111100011: data <= 32'h3820bc97;
    11'b01111100100: data <= 32'hb885bde1;
    11'b01111100101: data <= 32'hbca3bf00;
    11'b01111100110: data <= 32'hb404ba27;
    11'b01111100111: data <= 32'h39a33d0c;
    11'b01111101000: data <= 32'h30f5408f;
    11'b01111101001: data <= 32'hbcd93cb3;
    11'b01111101010: data <= 32'hbedab656;
    11'b01111101011: data <= 32'hbc96b500;
    11'b01111101100: data <= 32'hb84f3b79;
    11'b01111101101: data <= 32'had7d3c8c;
    11'b01111101110: data <= 32'h3b3db020;
    11'b01111101111: data <= 32'h4039baeb;
    11'b01111110000: data <= 32'h40213296;
    11'b01111110001: data <= 32'h380a3ea5;
    11'b01111110010: data <= 32'hb9cf3e21;
    11'b01111110011: data <= 32'hb2382ab8;
    11'b01111110100: data <= 32'h3b76bc64;
    11'b01111110101: data <= 32'h3949bd7d;
    11'b01111110110: data <= 32'hb971be33;
    11'b01111110111: data <= 32'hbb3fbefe;
    11'b01111111000: data <= 32'h3873bc67;
    11'b01111111001: data <= 32'h3e703554;
    11'b01111111010: data <= 32'h38513c23;
    11'b01111111011: data <= 32'hbe143431;
    11'b01111111100: data <= 32'hc0aeb8a7;
    11'b01111111101: data <= 32'hbe89a861;
    11'b01111111110: data <= 32'hbaa33c1c;
    11'b01111111111: data <= 32'hb83b39a1;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    