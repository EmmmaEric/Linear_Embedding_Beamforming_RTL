
module memory_rom_11(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbc9b3c60;
    11'b00000000001: data <= 32'hb8a238ca;
    11'b00000000010: data <= 32'h3a26b91e;
    11'b00000000011: data <= 32'h3f45b76f;
    11'b00000000100: data <= 32'h3ce63ced;
    11'b00000000101: data <= 32'hb4a740b4;
    11'b00000000110: data <= 32'hb9383ea8;
    11'b00000000111: data <= 32'h3817341a;
    11'b00000001000: data <= 32'h3d07b819;
    11'b00000001001: data <= 32'h35debadc;
    11'b00000001010: data <= 32'hb952bdaf;
    11'b00000001011: data <= 32'h2c3cbe8f;
    11'b00000001100: data <= 32'h3f34b9e5;
    11'b00000001101: data <= 32'h402b3769;
    11'b00000001110: data <= 32'h34f336b2;
    11'b00000001111: data <= 32'hbe30b94f;
    11'b00000010000: data <= 32'hbf70bbc0;
    11'b00000010001: data <= 32'hbd1a2a03;
    11'b00000010010: data <= 32'hbc203938;
    11'b00000010011: data <= 32'hbb54b681;
    11'b00000010100: data <= 32'hb1c2be9b;
    11'b00000010101: data <= 32'h3926bafe;
    11'b00000010110: data <= 32'h37253df7;
    11'b00000010111: data <= 32'hb69741aa;
    11'b00000011000: data <= 32'hb7ae3fd3;
    11'b00000011001: data <= 32'h35ce36f8;
    11'b00000011010: data <= 32'h38a3a879;
    11'b00000011011: data <= 32'hb65b3019;
    11'b00000011100: data <= 32'hbaf2b3ce;
    11'b00000011101: data <= 32'h38e9bafb;
    11'b00000011110: data <= 32'h4159b991;
    11'b00000011111: data <= 32'h417d2c07;
    11'b00000100000: data <= 32'h39663202;
    11'b00000100001: data <= 32'hbc63b672;
    11'b00000100010: data <= 32'hbc17b82a;
    11'b00000100011: data <= 32'hb4492b82;
    11'b00000100100: data <= 32'hb6e5ac59;
    11'b00000100101: data <= 32'hbc59be11;
    11'b00000100110: data <= 32'hbb18c114;
    11'b00000100111: data <= 32'h253bbd2e;
    11'b00000101000: data <= 32'h350b3cee;
    11'b00000101001: data <= 32'hb3b040aa;
    11'b00000101010: data <= 32'hb8a73d19;
    11'b00000101011: data <= 32'hb6022de5;
    11'b00000101100: data <= 32'hb875361e;
    11'b00000101101: data <= 32'hbd4a3c8c;
    11'b00000101110: data <= 32'hbcd839c0;
    11'b00000101111: data <= 32'h3936b746;
    11'b00000110000: data <= 32'h4142b9cd;
    11'b00000110001: data <= 32'h40fb305f;
    11'b00000110010: data <= 32'h38ea3a42;
    11'b00000110011: data <= 32'hb7fc388b;
    11'b00000110100: data <= 32'h318b3420;
    11'b00000110101: data <= 32'h3b4532bb;
    11'b00000110110: data <= 32'h3039b6fa;
    11'b00000110111: data <= 32'hbc90bfb9;
    11'b00000111000: data <= 32'hbc0ec170;
    11'b00000111001: data <= 32'h3521bded;
    11'b00000111010: data <= 32'h3bf138a3;
    11'b00000111011: data <= 32'h34923c91;
    11'b00000111100: data <= 32'hb9652cbc;
    11'b00000111101: data <= 32'hbc2cb76f;
    11'b00000111110: data <= 32'hbd5538c2;
    11'b00000111111: data <= 32'hbf4e3e68;
    11'b00001000000: data <= 32'hbe283a9f;
    11'b00001000001: data <= 32'h2d7aba40;
    11'b00001000010: data <= 32'h3e97bc00;
    11'b00001000011: data <= 32'h3dea36d2;
    11'b00001000100: data <= 32'h32a93e9d;
    11'b00001000101: data <= 32'habc63e38;
    11'b00001000110: data <= 32'h3c0e3b46;
    11'b00001000111: data <= 32'h3dd7382b;
    11'b00001001000: data <= 32'h30bbae22;
    11'b00001001001: data <= 32'hbd00bd3a;
    11'b00001001010: data <= 32'hb95fc01a;
    11'b00001001011: data <= 32'h3cedbd52;
    11'b00001001100: data <= 32'h400cada2;
    11'b00001001101: data <= 32'h3b489a78;
    11'b00001001110: data <= 32'hb856bab3;
    11'b00001001111: data <= 32'hbc2fb9f6;
    11'b00001010000: data <= 32'hbc903945;
    11'b00001010001: data <= 32'hbe383d90;
    11'b00001010010: data <= 32'hbea82d4e;
    11'b00001010011: data <= 32'hba0bbec0;
    11'b00001010100: data <= 32'h357abdea;
    11'b00001010101: data <= 32'h36213881;
    11'b00001010110: data <= 32'hb204401e;
    11'b00001010111: data <= 32'h2d733f32;
    11'b00001011000: data <= 32'h3c5c3bdb;
    11'b00001011001: data <= 32'h3c3f3aac;
    11'b00001011010: data <= 32'hb7da3a61;
    11'b00001011011: data <= 32'hbe1ea1bd;
    11'b00001011100: data <= 32'hb487bbd1;
    11'b00001011101: data <= 32'h3ffbbc00;
    11'b00001011110: data <= 32'h4146b6f8;
    11'b00001011111: data <= 32'h3cdcb732;
    11'b00001100000: data <= 32'hb275bb02;
    11'b00001100001: data <= 32'hb471b72d;
    11'b00001100010: data <= 32'ha71039f3;
    11'b00001100011: data <= 32'hb9593ada;
    11'b00001100100: data <= 32'hbe2dbb1b;
    11'b00001100101: data <= 32'hbd8ec111;
    11'b00001100110: data <= 32'hb7c9bf87;
    11'b00001100111: data <= 32'hac4735bb;
    11'b00001101000: data <= 32'hb26e3e65;
    11'b00001101001: data <= 32'h29933c18;
    11'b00001101010: data <= 32'h3874361f;
    11'b00001101011: data <= 32'h2df03bc9;
    11'b00001101100: data <= 32'hbd7c3ee2;
    11'b00001101101: data <= 32'hbf933c95;
    11'b00001101110: data <= 32'hb3d0b338;
    11'b00001101111: data <= 32'h3fd8ba7a;
    11'b00001110000: data <= 32'h409cb669;
    11'b00001110001: data <= 32'h3b7eacab;
    11'b00001110010: data <= 32'h309cae8b;
    11'b00001110011: data <= 32'h3aa9346d;
    11'b00001110100: data <= 32'h3d553b93;
    11'b00001110101: data <= 32'h338f384a;
    11'b00001110110: data <= 32'hbd65bd25;
    11'b00001110111: data <= 32'hbe1ec14d;
    11'b00001111000: data <= 32'hb694bf94;
    11'b00001111001: data <= 32'h361cad0a;
    11'b00001111010: data <= 32'h340b37ce;
    11'b00001111011: data <= 32'h25a3b59a;
    11'b00001111100: data <= 32'ha510b822;
    11'b00001111101: data <= 32'hb9243b50;
    11'b00001111110: data <= 32'hbf55405a;
    11'b00001111111: data <= 32'hc0323dee;
    11'b00010000000: data <= 32'hb918b4ae;
    11'b00010000001: data <= 32'h3c31bbe0;
    11'b00010000010: data <= 32'h3c87b202;
    11'b00010000011: data <= 32'h3248395e;
    11'b00010000100: data <= 32'h34ca3a8a;
    11'b00010000101: data <= 32'h3e943b35;
    11'b00010000110: data <= 32'h403a3cbd;
    11'b00010000111: data <= 32'h38563a01;
    11'b00010001000: data <= 32'hbd4bb9c1;
    11'b00010001001: data <= 32'hbd08bf5d;
    11'b00010001010: data <= 32'h3583bdb8;
    11'b00010001011: data <= 32'h3d43b768;
    11'b00010001100: data <= 32'h3addb8f0;
    11'b00010001101: data <= 32'h301cbdf9;
    11'b00010001110: data <= 32'hae4ebc75;
    11'b00010001111: data <= 32'hb7e43a76;
    11'b00010010000: data <= 32'hbdc7400c;
    11'b00010010001: data <= 32'hbfc33b51;
    11'b00010010010: data <= 32'hbcd2bc48;
    11'b00010010011: data <= 32'hb2bcbdc3;
    11'b00010010100: data <= 32'hb247ac03;
    11'b00010010101: data <= 32'hb8563c6a;
    11'b00010010110: data <= 32'h33b73c5a;
    11'b00010010111: data <= 32'h3f103b14;
    11'b00010011000: data <= 32'h3fa63d0a;
    11'b00010011001: data <= 32'h2c293d94;
    11'b00010011010: data <= 32'hbe453834;
    11'b00010011011: data <= 32'hbb42b84f;
    11'b00010011100: data <= 32'h3c60b9ed;
    11'b00010011101: data <= 32'h3fc2b89c;
    11'b00010011110: data <= 32'h3c68bc61;
    11'b00010011111: data <= 32'h347fbefe;
    11'b00010100000: data <= 32'h3744bc12;
    11'b00010100001: data <= 32'h388e3ab4;
    11'b00010100010: data <= 32'hb57e3e2c;
    11'b00010100011: data <= 32'hbdd59ea4;
    11'b00010100100: data <= 32'hbe54bfa1;
    11'b00010100101: data <= 32'hbc3bbf39;
    11'b00010100110: data <= 32'hbb0eb02b;
    11'b00010100111: data <= 32'hba5e3a91;
    11'b00010101000: data <= 32'h2f7135c7;
    11'b00010101001: data <= 32'h3d2e2ddb;
    11'b00010101010: data <= 32'h3c1b3c31;
    11'b00010101011: data <= 32'hba4c401a;
    11'b00010101100: data <= 32'hbfa53ec2;
    11'b00010101101: data <= 32'hba38376e;
    11'b00010101110: data <= 32'h3ccbb445;
    11'b00010101111: data <= 32'h3e9cb6c4;
    11'b00010110000: data <= 32'h393dba44;
    11'b00010110001: data <= 32'h34cfbc5d;
    11'b00010110010: data <= 32'h3d32b58f;
    11'b00010110011: data <= 32'h3fb73c20;
    11'b00010110100: data <= 32'h3a963cb1;
    11'b00010110101: data <= 32'hbb89b80f;
    11'b00010110110: data <= 32'hbe45c023;
    11'b00010110111: data <= 32'hbc2cbeba;
    11'b00010111000: data <= 32'hb8aab467;
    11'b00010111001: data <= 32'hb6eea8bc;
    11'b00010111010: data <= 32'h2d68bc06;
    11'b00010111011: data <= 32'h39a1bc4a;
    11'b00010111100: data <= 32'h332d3923;
    11'b00010111101: data <= 32'hbd2a40a2;
    11'b00010111110: data <= 32'hc0074029;
    11'b00010111111: data <= 32'hbb5a38a5;
    11'b00011000000: data <= 32'h3829b4eb;
    11'b00011000001: data <= 32'h37d7b1f6;
    11'b00011000010: data <= 32'hb588aa98;
    11'b00011000011: data <= 32'h2e14b081;
    11'b00011000100: data <= 32'h3f983508;
    11'b00011000101: data <= 32'h41853ccf;
    11'b00011000110: data <= 32'h3d5f3cba;
    11'b00011000111: data <= 32'hb9e1b0de;
    11'b00011001000: data <= 32'hbcfebd1c;
    11'b00011001001: data <= 32'hb519bbc3;
    11'b00011001010: data <= 32'h3580b4bd;
    11'b00011001011: data <= 32'h324abb52;
    11'b00011001100: data <= 32'h30e1c065;
    11'b00011001101: data <= 32'h3772bfa7;
    11'b00011001110: data <= 32'h31f134eb;
    11'b00011001111: data <= 32'hbb74402d;
    11'b00011010000: data <= 32'hbe893e39;
    11'b00011010001: data <= 32'hbc89b0e9;
    11'b00011010010: data <= 32'hb809ba21;
    11'b00011010011: data <= 32'hbb16a94b;
    11'b00011010100: data <= 32'hbd6837f8;
    11'b00011010101: data <= 32'hb38734a8;
    11'b00011010110: data <= 32'h3fa73572;
    11'b00011010111: data <= 32'h41383c5a;
    11'b00011011000: data <= 32'h3b973dfa;
    11'b00011011001: data <= 32'hbb9b3adb;
    11'b00011011010: data <= 32'hbb122c5e;
    11'b00011011011: data <= 32'h38161d61;
    11'b00011011100: data <= 32'h3c67ae62;
    11'b00011011101: data <= 32'h37debd09;
    11'b00011011110: data <= 32'h30fbc107;
    11'b00011011111: data <= 32'h39c1bfc3;
    11'b00011100000: data <= 32'h3c113450;
    11'b00011100001: data <= 32'h32853e5c;
    11'b00011100010: data <= 32'hbadf38ac;
    11'b00011100011: data <= 32'hbcb1bc61;
    11'b00011100100: data <= 32'hbcc6bcbf;
    11'b00011100101: data <= 32'hbe931a57;
    11'b00011100110: data <= 32'hbf1a379e;
    11'b00011100111: data <= 32'hb792b2d8;
    11'b00011101000: data <= 32'h3da7b794;
    11'b00011101001: data <= 32'h3eca38bc;
    11'b00011101010: data <= 32'h25d43f30;
    11'b00011101011: data <= 32'hbd643f5f;
    11'b00011101100: data <= 32'hb9643c9b;
    11'b00011101101: data <= 32'h3ab6398a;
    11'b00011101110: data <= 32'h3c1832f0;
    11'b00011101111: data <= 32'h2955bb35;
    11'b00011110000: data <= 32'hadb6bf6c;
    11'b00011110001: data <= 32'h3cd7bcee;
    11'b00011110010: data <= 32'h405e380f;
    11'b00011110011: data <= 32'h3dd23ca8;
    11'b00011110100: data <= 32'hadcfaebb;
    11'b00011110101: data <= 32'hbb8ebdd1;
    11'b00011110110: data <= 32'hbc73bc50;
    11'b00011110111: data <= 32'hbd782e06;
    11'b00011111000: data <= 32'hbdaca915;
    11'b00011111001: data <= 32'hb7b6bd88;
    11'b00011111010: data <= 32'h3a45bee4;
    11'b00011111011: data <= 32'h39ebae0a;
    11'b00011111100: data <= 32'hb9543f38;
    11'b00011111101: data <= 32'hbdf1404a;
    11'b00011111110: data <= 32'hb8e63d41;
    11'b00011111111: data <= 32'h37bf39aa;
    11'b00100000000: data <= 32'h2c01376b;
    11'b00100000001: data <= 32'hbc28b074;
    11'b00100000010: data <= 32'hb8bbba40;
    11'b00100000011: data <= 32'h3e13b66e;
    11'b00100000100: data <= 32'h41d039da;
    11'b00100000101: data <= 32'h40153c05;
    11'b00100000110: data <= 32'h3336aaad;
    11'b00100000111: data <= 32'hb892baef;
    11'b00100001000: data <= 32'hb5b3b4c4;
    11'b00100001001: data <= 32'hb59235fd;
    11'b00100001010: data <= 32'hb927b8d5;
    11'b00100001011: data <= 32'hb596c0e7;
    11'b00100001100: data <= 32'h369cc14d;
    11'b00100001101: data <= 32'h36c8b8b8;
    11'b00100001110: data <= 32'hb8213de6;
    11'b00100001111: data <= 32'hbc3a3e52;
    11'b00100010000: data <= 32'hb8443826;
    11'b00100010001: data <= 32'hb2d83072;
    11'b00100010010: data <= 32'hbcb6385b;
    11'b00100010011: data <= 32'hc04c3819;
    11'b00100010100: data <= 32'hbc85ae4f;
    11'b00100010101: data <= 32'h3d8ab131;
    11'b00100010110: data <= 32'h416938c3;
    11'b00100010111: data <= 32'h3e793c2b;
    11'b00100011000: data <= 32'hab893902;
    11'b00100011001: data <= 32'hb41b3555;
    11'b00100011010: data <= 32'h386e3a5a;
    11'b00100011011: data <= 32'h390f3a8f;
    11'b00100011100: data <= 32'hb052ba0e;
    11'b00100011101: data <= 32'hb56fc16a;
    11'b00100011110: data <= 32'h36b3c15c;
    11'b00100011111: data <= 32'h3b69b8dc;
    11'b00100100000: data <= 32'h375f3c01;
    11'b00100100001: data <= 32'hb1373854;
    11'b00100100010: data <= 32'hb4acb8f2;
    11'b00100100011: data <= 32'hb965b7d5;
    11'b00100100100: data <= 32'hbf7a3876;
    11'b00100100101: data <= 32'hc13939a6;
    11'b00100100110: data <= 32'hbd9bb48a;
    11'b00100100111: data <= 32'h3b05ba6c;
    11'b00100101000: data <= 32'h3ef0a174;
    11'b00100101001: data <= 32'h38323c31;
    11'b00100101010: data <= 32'hb9343d69;
    11'b00100101011: data <= 32'hae193d5f;
    11'b00100101100: data <= 32'h3c453e39;
    11'b00100101101: data <= 32'h3ae63ce9;
    11'b00100101110: data <= 32'hb659b5a8;
    11'b00100101111: data <= 32'hb965bff9;
    11'b00100110000: data <= 32'h38e0bf59;
    11'b00100110001: data <= 32'h3f40b257;
    11'b00100110010: data <= 32'h3e84390f;
    11'b00100110011: data <= 32'h39afb4ed;
    11'b00100110100: data <= 32'h2d72bd16;
    11'b00100110101: data <= 32'hb80fb8aa;
    11'b00100110110: data <= 32'hbe2b39b4;
    11'b00100110111: data <= 32'hc05037b5;
    11'b00100111000: data <= 32'hbd16bca1;
    11'b00100111001: data <= 32'h34d9bfd4;
    11'b00100111010: data <= 32'h3919ba96;
    11'b00100111011: data <= 32'hb71f3adb;
    11'b00100111100: data <= 32'hbc033e1d;
    11'b00100111101: data <= 32'h19a03dd5;
    11'b00100111110: data <= 32'h3be73e13;
    11'b00100111111: data <= 32'h328d3d86;
    11'b00101000000: data <= 32'hbd7a35d4;
    11'b00101000001: data <= 32'hbd40ba65;
    11'b00101000010: data <= 32'h3972b9f1;
    11'b00101000011: data <= 32'h40bd33ff;
    11'b00101000100: data <= 32'h4058376e;
    11'b00101000101: data <= 32'h3c14b818;
    11'b00101000110: data <= 32'h36b7bbf3;
    11'b00101000111: data <= 32'h33452ca9;
    11'b00101001000: data <= 32'hb6b83c84;
    11'b00101001001: data <= 32'hbc9231c6;
    11'b00101001010: data <= 32'hbb50c010;
    11'b00101001011: data <= 32'haabbc1af;
    11'b00101001100: data <= 32'h2d64bd6d;
    11'b00101001101: data <= 32'hb8e2380d;
    11'b00101001110: data <= 32'hb9c43ba3;
    11'b00101001111: data <= 32'h32a33898;
    11'b00101010000: data <= 32'h388b39ef;
    11'b00101010001: data <= 32'hba8c3cff;
    11'b00101010010: data <= 32'hc0e03bdd;
    11'b00101010011: data <= 32'hbfb62e66;
    11'b00101010100: data <= 32'h3785b1e0;
    11'b00101010101: data <= 32'h40423494;
    11'b00101010110: data <= 32'h3eb03652;
    11'b00101010111: data <= 32'h388baf9f;
    11'b00101011000: data <= 32'h3861a81c;
    11'b00101011001: data <= 32'h3c643c7b;
    11'b00101011010: data <= 32'h3a0e3ebd;
    11'b00101011011: data <= 32'hb50d30fa;
    11'b00101011100: data <= 32'hb9a6c06f;
    11'b00101011101: data <= 32'hb00ac19f;
    11'b00101011110: data <= 32'h34d3bd01;
    11'b00101011111: data <= 32'h2edd31d4;
    11'b00101100000: data <= 32'h2f98aa59;
    11'b00101100001: data <= 32'h38a9b9ed;
    11'b00101100010: data <= 32'h347cb252;
    11'b00101100011: data <= 32'hbda53c2d;
    11'b00101100100: data <= 32'hc1b63ce9;
    11'b00101100101: data <= 32'hc0413230;
    11'b00101100110: data <= 32'h2c3db85b;
    11'b00101100111: data <= 32'h3cb8b3da;
    11'b00101101000: data <= 32'h36aa3414;
    11'b00101101001: data <= 32'hb51d365e;
    11'b00101101010: data <= 32'h37b33ad4;
    11'b00101101011: data <= 32'h3e8d3f6a;
    11'b00101101100: data <= 32'h3d054025;
    11'b00101101101: data <= 32'hb476380c;
    11'b00101101110: data <= 32'hbb85be0a;
    11'b00101101111: data <= 32'had05bf4c;
    11'b00101110000: data <= 32'h3b9bb88d;
    11'b00101110001: data <= 32'h3c8128fd;
    11'b00101110010: data <= 32'h3bd0bb43;
    11'b00101110011: data <= 32'h3beebe9d;
    11'b00101110100: data <= 32'h372bb8d8;
    11'b00101110101: data <= 32'hbc4c3c46;
    11'b00101110110: data <= 32'hc08f3c88;
    11'b00101110111: data <= 32'hbf08b6ce;
    11'b00101111000: data <= 32'hb4b8be18;
    11'b00101111001: data <= 32'h2d5dbc2f;
    11'b00101111010: data <= 32'hba6ca175;
    11'b00101111011: data <= 32'hbc003829;
    11'b00101111100: data <= 32'h36b23b86;
    11'b00101111101: data <= 32'h3ead3ee5;
    11'b00101111110: data <= 32'h3ae8400f;
    11'b00101111111: data <= 32'hbc333c23;
    11'b00110000000: data <= 32'hbe3eb521;
    11'b00110000001: data <= 32'haf52b7d7;
    11'b00110000010: data <= 32'h3da132e8;
    11'b00110000011: data <= 32'h3e7b2b6d;
    11'b00110000100: data <= 32'h3ce3bcd0;
    11'b00110000101: data <= 32'h3cbbbe98;
    11'b00110000110: data <= 32'h3c1db1ad;
    11'b00110000111: data <= 32'h296f3dcf;
    11'b00110001000: data <= 32'hbc2b3bab;
    11'b00110001001: data <= 32'hbc40bca3;
    11'b00110001010: data <= 32'hb715c0ae;
    11'b00110001011: data <= 32'hb859be2a;
    11'b00110001100: data <= 32'hbcffb468;
    11'b00110001101: data <= 32'hbbcb2b4a;
    11'b00110001110: data <= 32'h388e2b85;
    11'b00110001111: data <= 32'h3d8a39f6;
    11'b00110010000: data <= 32'h21a03e4d;
    11'b00110010001: data <= 32'hc0113dbd;
    11'b00110010010: data <= 32'hc0513916;
    11'b00110010011: data <= 32'hb4b135b4;
    11'b00110010100: data <= 32'h3ceb3852;
    11'b00110010101: data <= 32'h3c772c86;
    11'b00110010110: data <= 32'h38c5bb95;
    11'b00110010111: data <= 32'h3c0fbb15;
    11'b00110011000: data <= 32'h3eba3a1a;
    11'b00110011001: data <= 32'h3d0e4003;
    11'b00110011010: data <= 32'h2cce3b97;
    11'b00110011011: data <= 32'hb84ebd75;
    11'b00110011100: data <= 32'hb66cc098;
    11'b00110011101: data <= 32'hb751bd2d;
    11'b00110011110: data <= 32'hba0bb57e;
    11'b00110011111: data <= 32'hb449b9f5;
    11'b00110100000: data <= 32'h3b9bbd2b;
    11'b00110100001: data <= 32'h3c9cb7b0;
    11'b00110100010: data <= 32'hb87a3c20;
    11'b00110100011: data <= 32'hc0dd3e21;
    11'b00110100100: data <= 32'hc0803ace;
    11'b00110100101: data <= 32'hb7cb33cb;
    11'b00110100110: data <= 32'h37563193;
    11'b00110100111: data <= 32'hb176ac7b;
    11'b00110101000: data <= 32'hb88ab824;
    11'b00110101001: data <= 32'h38cdab82;
    11'b00110101010: data <= 32'h40183de5;
    11'b00110101011: data <= 32'h3f7c40a6;
    11'b00110101100: data <= 32'h361b3c90;
    11'b00110101101: data <= 32'hb88aba70;
    11'b00110101110: data <= 32'hb565bd21;
    11'b00110101111: data <= 32'h2d4fb5a2;
    11'b00110110000: data <= 32'h315eb07d;
    11'b00110110001: data <= 32'h3878bda9;
    11'b00110110010: data <= 32'h3d4ac09b;
    11'b00110110011: data <= 32'h3cdbbcb5;
    11'b00110110100: data <= 32'hb56e3a7e;
    11'b00110110101: data <= 32'hbf573d94;
    11'b00110110110: data <= 32'hbe9635a3;
    11'b00110110111: data <= 32'hb821b8d6;
    11'b00110111000: data <= 32'hb71bb8a0;
    11'b00110111001: data <= 32'hbdefb539;
    11'b00110111010: data <= 32'hbe35b575;
    11'b00110111011: data <= 32'h341e2f1e;
    11'b00110111100: data <= 32'h40043d51;
    11'b00110111101: data <= 32'h3e6b4029;
    11'b00110111110: data <= 32'hb33e3d74;
    11'b00110111111: data <= 32'hbc763230;
    11'b00111000000: data <= 32'hb60f3078;
    11'b00111000001: data <= 32'h386439fb;
    11'b00111000010: data <= 32'h39b03218;
    11'b00111000011: data <= 32'h3a63be71;
    11'b00111000100: data <= 32'h3d6bc0da;
    11'b00111000101: data <= 32'h3e1bbb8f;
    11'b00111000110: data <= 32'h38c53c5d;
    11'b00111000111: data <= 32'hb8203ce9;
    11'b00111001000: data <= 32'hb911b5ad;
    11'b00111001001: data <= 32'hb542bdbf;
    11'b00111001010: data <= 32'hbb94bc4b;
    11'b00111001011: data <= 32'hc01fb79a;
    11'b00111001100: data <= 32'hbf07b8a8;
    11'b00111001101: data <= 32'h3443b8d7;
    11'b00111001110: data <= 32'h3ee53482;
    11'b00111001111: data <= 32'h3a743d43;
    11'b00111010000: data <= 32'hbcc33da9;
    11'b00111010001: data <= 32'hbeda3c07;
    11'b00111010010: data <= 32'hb7b23c7b;
    11'b00111010011: data <= 32'h385b3d59;
    11'b00111010100: data <= 32'h35a13631;
    11'b00111010101: data <= 32'h2f8cbd5d;
    11'b00111010110: data <= 32'h3b31bef6;
    11'b00111010111: data <= 32'h3f55ab23;
    11'b00111011000: data <= 32'h3ea53e8d;
    11'b00111011001: data <= 32'h39e63cb1;
    11'b00111011010: data <= 32'h3211b97d;
    11'b00111011011: data <= 32'hab9cbe11;
    11'b00111011100: data <= 32'hba9fba4d;
    11'b00111011101: data <= 32'hbea7b499;
    11'b00111011110: data <= 32'hbc8dbc37;
    11'b00111011111: data <= 32'h3900bf2d;
    11'b00111100000: data <= 32'h3de2bc4f;
    11'b00111100001: data <= 32'h30cd372f;
    11'b00111100010: data <= 32'hbec53cf8;
    11'b00111100011: data <= 32'hbf223ca9;
    11'b00111100100: data <= 32'hb7543c7e;
    11'b00111100101: data <= 32'h2cd33c67;
    11'b00111100110: data <= 32'hba3334b1;
    11'b00111100111: data <= 32'hbcb2bb3c;
    11'b00111101000: data <= 32'h30c1baec;
    11'b00111101001: data <= 32'h3f9739e4;
    11'b00111101010: data <= 32'h40613fcd;
    11'b00111101011: data <= 32'h3cb43cc2;
    11'b00111101100: data <= 32'h3561b657;
    11'b00111101101: data <= 32'h2d9db93f;
    11'b00111101110: data <= 32'hb494345b;
    11'b00111101111: data <= 32'hb9cf3407;
    11'b00111110000: data <= 32'hb412bd9b;
    11'b00111110001: data <= 32'h3c07c16b;
    11'b00111110010: data <= 32'h3d98bfae;
    11'b00111110011: data <= 32'h305d1f97;
    11'b00111110100: data <= 32'hbcf93bd5;
    11'b00111110101: data <= 32'hbc4e394a;
    11'b00111110110: data <= 32'hb12d34af;
    11'b00111110111: data <= 32'hb7f4352a;
    11'b00111111000: data <= 32'hbfec2577;
    11'b00111111001: data <= 32'hc0a2b911;
    11'b00111111010: data <= 32'hb756b7f7;
    11'b00111111011: data <= 32'h3ebe39e3;
    11'b00111111100: data <= 32'h3fa03e83;
    11'b00111111101: data <= 32'h38ed3c6f;
    11'b00111111110: data <= 32'hb25d3464;
    11'b00111111111: data <= 32'h28c33938;
    11'b01000000000: data <= 32'h33c23e29;
    11'b01000000001: data <= 32'ha5c53b0f;
    11'b01000000010: data <= 32'h2fe1bd8a;
    11'b01000000011: data <= 32'h3be7c19b;
    11'b01000000100: data <= 32'h3dc2bf0e;
    11'b01000000101: data <= 32'h3a0b335a;
    11'b01000000110: data <= 32'ha9943a6a;
    11'b01000000111: data <= 32'h2eebad90;
    11'b01000001000: data <= 32'h35a6b94e;
    11'b01000001001: data <= 32'hba05b4c9;
    11'b01000001010: data <= 32'hc108ae9b;
    11'b01000001011: data <= 32'hc140b924;
    11'b01000001100: data <= 32'hb86fbb53;
    11'b01000001101: data <= 32'h3d74b1f0;
    11'b01000001110: data <= 32'h3c513993;
    11'b01000001111: data <= 32'hb7043a8a;
    11'b01000010000: data <= 32'hbb433a80;
    11'b01000010001: data <= 32'hac063e56;
    11'b01000010010: data <= 32'h36dc4087;
    11'b01000010011: data <= 32'haedd3cf1;
    11'b01000010100: data <= 32'hb6c6bc2a;
    11'b01000010101: data <= 32'h3622c02f;
    11'b01000010110: data <= 32'h3d9bba8a;
    11'b01000010111: data <= 32'h3e193aeb;
    11'b01000011000: data <= 32'h3c9d3a11;
    11'b01000011001: data <= 32'h3c61b893;
    11'b01000011010: data <= 32'h3aa7bbee;
    11'b01000011011: data <= 32'hb82ab0ee;
    11'b01000011100: data <= 32'hc03332a2;
    11'b01000011101: data <= 32'hbff0ba44;
    11'b01000011110: data <= 32'hb067bf33;
    11'b01000011111: data <= 32'h3c7ebdec;
    11'b01000100000: data <= 32'h34ccb5ac;
    11'b01000100001: data <= 32'hbca63632;
    11'b01000100010: data <= 32'hbc7e3a8c;
    11'b01000100011: data <= 32'h2add3e46;
    11'b01000100100: data <= 32'h34454017;
    11'b01000100101: data <= 32'hbb703c7e;
    11'b01000100110: data <= 32'hbe91b8e6;
    11'b01000100111: data <= 32'hb881bc7a;
    11'b01000101000: data <= 32'h3cad317f;
    11'b01000101001: data <= 32'h3f763d4d;
    11'b01000101010: data <= 32'h3e4c39b0;
    11'b01000101011: data <= 32'h3d35b87b;
    11'b01000101100: data <= 32'h3c0ab6da;
    11'b01000101101: data <= 32'h27a73a93;
    11'b01000101110: data <= 32'hbc573b8b;
    11'b01000101111: data <= 32'hbb75ba78;
    11'b01000110000: data <= 32'h3641c0fe;
    11'b01000110001: data <= 32'h3c10c09c;
    11'b01000110010: data <= 32'h28f0bb32;
    11'b01000110011: data <= 32'hbc022891;
    11'b01000110100: data <= 32'hb81a3477;
    11'b01000110101: data <= 32'h384b3970;
    11'b01000110110: data <= 32'h27203c86;
    11'b01000110111: data <= 32'hbf9339b7;
    11'b01000111000: data <= 32'hc188b53f;
    11'b01000111001: data <= 32'hbd3fb848;
    11'b01000111010: data <= 32'h3a81373b;
    11'b01000111011: data <= 32'h3e0d3c77;
    11'b01000111100: data <= 32'h3bc23763;
    11'b01000111101: data <= 32'h395db326;
    11'b01000111110: data <= 32'h3ac338fe;
    11'b01000111111: data <= 32'h38764024;
    11'b01001000000: data <= 32'hb23c3efd;
    11'b01001000001: data <= 32'hb48bb8c4;
    11'b01001000010: data <= 32'h3808c0f9;
    11'b01001000011: data <= 32'h3b52c03c;
    11'b01001000100: data <= 32'h354db901;
    11'b01001000101: data <= 32'hac7dac07;
    11'b01001000110: data <= 32'h3931b775;
    11'b01001000111: data <= 32'h3cffb6f9;
    11'b01001001000: data <= 32'h22583412;
    11'b01001001001: data <= 32'hc099370d;
    11'b01001001010: data <= 32'hc21cb349;
    11'b01001001011: data <= 32'hbd9eb923;
    11'b01001001100: data <= 32'h3830b22f;
    11'b01001001101: data <= 32'h396f3300;
    11'b01001001110: data <= 32'hb30da95b;
    11'b01001001111: data <= 32'hb45c2903;
    11'b01001010000: data <= 32'h38b13d9a;
    11'b01001010001: data <= 32'h3a934194;
    11'b01001010010: data <= 32'h2125404b;
    11'b01001010011: data <= 32'hb860b381;
    11'b01001010100: data <= 32'haa23bf05;
    11'b01001010101: data <= 32'h3951bc38;
    11'b01001010110: data <= 32'h3a6632eb;
    11'b01001010111: data <= 32'h3b972a8e;
    11'b01001011000: data <= 32'h3e93bc03;
    11'b01001011001: data <= 32'h3f4cbc1f;
    11'b01001011010: data <= 32'h35092f1a;
    11'b01001011011: data <= 32'hbf5c3965;
    11'b01001011100: data <= 32'hc0a4b167;
    11'b01001011101: data <= 32'hba85bcd9;
    11'b01001011110: data <= 32'h36debd28;
    11'b01001011111: data <= 32'hb057bacb;
    11'b01001100000: data <= 32'hbcc2b8eb;
    11'b01001100001: data <= 32'hba3aad00;
    11'b01001100010: data <= 32'h38ce3d4b;
    11'b01001100011: data <= 32'h3ab24101;
    11'b01001100100: data <= 32'hb7e73f9e;
    11'b01001100101: data <= 32'hbe312c9f;
    11'b01001100110: data <= 32'hbc0bba09;
    11'b01001100111: data <= 32'h340c311e;
    11'b01001101000: data <= 32'h3bbc3bba;
    11'b01001101001: data <= 32'h3d28301f;
    11'b01001101010: data <= 32'h3f3ebc92;
    11'b01001101011: data <= 32'h3fb3ba42;
    11'b01001101100: data <= 32'h3a373ad3;
    11'b01001101101: data <= 32'hba693dac;
    11'b01001101110: data <= 32'hbc401f7e;
    11'b01001101111: data <= 32'h9b7dbec5;
    11'b01001110000: data <= 32'h3771c006;
    11'b01001110001: data <= 32'hb82fbd86;
    11'b01001110010: data <= 32'hbd5abb90;
    11'b01001110011: data <= 32'hb6b1b895;
    11'b01001110100: data <= 32'h3c4d3685;
    11'b01001110101: data <= 32'h3a793da1;
    11'b01001110110: data <= 32'hbcd93cea;
    11'b01001110111: data <= 32'hc11a326e;
    11'b01001111000: data <= 32'hbf14ac45;
    11'b01001111001: data <= 32'hb07b39f1;
    11'b01001111010: data <= 32'h38df3c19;
    11'b01001111011: data <= 32'h3933adbe;
    11'b01001111100: data <= 32'h3c1bbc10;
    11'b01001111101: data <= 32'h3e1518d2;
    11'b01001111110: data <= 32'h3c983fdc;
    11'b01001111111: data <= 32'h31874080;
    11'b01010000000: data <= 32'hafa934f1;
    11'b01010000001: data <= 32'h365abe84;
    11'b01010000010: data <= 32'h36c2bf20;
    11'b01010000011: data <= 32'hb6e8bbe7;
    11'b01010000100: data <= 32'hb984bac3;
    11'b01010000101: data <= 32'h38b6bcb3;
    11'b01010000110: data <= 32'h3f4fba37;
    11'b01010000111: data <= 32'h3b6733e5;
    11'b01010001000: data <= 32'hbe113937;
    11'b01010001001: data <= 32'hc19332d1;
    11'b01010001010: data <= 32'hbf1d2278;
    11'b01010001011: data <= 32'hb47d3651;
    11'b01010001100: data <= 32'haec134dd;
    11'b01010001101: data <= 32'hb8cdb912;
    11'b01010001110: data <= 32'hb1d7bb5a;
    11'b01010001111: data <= 32'h3ba1391d;
    11'b01010010000: data <= 32'h3d30413f;
    11'b01010010001: data <= 32'h385c4134;
    11'b01010010010: data <= 32'hacc2389b;
    11'b01010010011: data <= 32'h2a32bbd9;
    11'b01010010100: data <= 32'h3083b94d;
    11'b01010010101: data <= 32'hb0da2e55;
    11'b01010010110: data <= 32'h30fcb6de;
    11'b01010010111: data <= 32'h3e10be50;
    11'b01010011000: data <= 32'h40c8be14;
    11'b01010011001: data <= 32'h3cc2b2cb;
    11'b01010011010: data <= 32'hbc6c3937;
    11'b01010011011: data <= 32'hbfff3484;
    11'b01010011100: data <= 32'hbbc3b5b2;
    11'b01010011101: data <= 32'hadd3b7f3;
    11'b01010011110: data <= 32'hba3db97b;
    11'b01010011111: data <= 32'hbecfbce8;
    11'b01010100000: data <= 32'hbc08bc37;
    11'b01010100001: data <= 32'h39a43894;
    11'b01010100010: data <= 32'h3d2e4092;
    11'b01010100011: data <= 32'h33d04059;
    11'b01010100100: data <= 32'hbabe3905;
    11'b01010100101: data <= 32'hba8daf81;
    11'b01010100110: data <= 32'hb5013965;
    11'b01010100111: data <= 32'haae13cad;
    11'b01010101000: data <= 32'h377aac22;
    11'b01010101001: data <= 32'h3e8ebeaf;
    11'b01010101010: data <= 32'h40b1bde1;
    11'b01010101011: data <= 32'h3dbf3461;
    11'b01010101100: data <= 32'hb2223d1a;
    11'b01010101101: data <= 32'hb9073815;
    11'b01010101110: data <= 32'h310eb9cd;
    11'b01010101111: data <= 32'h33fcbc9e;
    11'b01010110000: data <= 32'hbc61bcb8;
    11'b01010110001: data <= 32'hc016bdd7;
    11'b01010110010: data <= 32'hbb68bd88;
    11'b01010110011: data <= 32'h3c20b39e;
    11'b01010110100: data <= 32'h3d433c5a;
    11'b01010110101: data <= 32'hb54f3cc5;
    11'b01010110110: data <= 32'hbefd3717;
    11'b01010110111: data <= 32'hbe2b37a6;
    11'b01010111000: data <= 32'hb93c3dc5;
    11'b01010111001: data <= 32'hb4d33e1d;
    11'b01010111010: data <= 32'hadc4ae83;
    11'b01010111011: data <= 32'h3a23be53;
    11'b01010111100: data <= 32'h3ea4bac9;
    11'b01010111101: data <= 32'h3dfe3d04;
    11'b01010111110: data <= 32'h39684023;
    11'b01010111111: data <= 32'h37ec3a65;
    11'b01011000000: data <= 32'h3b0bb9bb;
    11'b01011000001: data <= 32'h36c6bbce;
    11'b01011000010: data <= 32'hbc17b9b5;
    11'b01011000011: data <= 32'hbe49bc73;
    11'b01011000100: data <= 32'had1ebec6;
    11'b01011000101: data <= 32'h3ef0bd3d;
    11'b01011000110: data <= 32'h3dccb3e0;
    11'b01011000111: data <= 32'hb923346f;
    11'b01011001000: data <= 32'hc004327f;
    11'b01011001001: data <= 32'hbdf8386e;
    11'b01011001010: data <= 32'hb8b93d23;
    11'b01011001011: data <= 32'hba0d3c00;
    11'b01011001100: data <= 32'hbcebb8a5;
    11'b01011001101: data <= 32'hb8dbbe16;
    11'b01011001110: data <= 32'h39f7b3f1;
    11'b01011001111: data <= 32'h3d753fa4;
    11'b01011010000: data <= 32'h3c1540c1;
    11'b01011010001: data <= 32'h39ea3b43;
    11'b01011010010: data <= 32'h3a15b497;
    11'b01011010011: data <= 32'h33762949;
    11'b01011010100: data <= 32'hba533835;
    11'b01011010101: data <= 32'hba65b5a3;
    11'b01011010110: data <= 32'h3a8fbf2e;
    11'b01011010111: data <= 32'h408ac002;
    11'b01011011000: data <= 32'h3e69bb49;
    11'b01011011001: data <= 32'hb67821eb;
    11'b01011011010: data <= 32'hbd3a30ab;
    11'b01011011011: data <= 32'hb8603375;
    11'b01011011100: data <= 32'hac9937f9;
    11'b01011011101: data <= 32'hbc7f2c2b;
    11'b01011011110: data <= 32'hc089bca0;
    11'b01011011111: data <= 32'hbe91be5d;
    11'b01011100000: data <= 32'h3250b1f9;
    11'b01011100001: data <= 32'h3cc83e98;
    11'b01011100010: data <= 32'h3a113f55;
    11'b01011100011: data <= 32'h2eaa3941;
    11'b01011100100: data <= 32'ha52a3471;
    11'b01011100101: data <= 32'hb2923d3a;
    11'b01011100110: data <= 32'hb9563f3b;
    11'b01011100111: data <= 32'hb6773573;
    11'b01011101000: data <= 32'h3c06bebb;
    11'b01011101001: data <= 32'h4044bfe8;
    11'b01011101010: data <= 32'h3e54b8a6;
    11'b01011101011: data <= 32'h334c3815;
    11'b01011101100: data <= 32'ha0c13590;
    11'b01011101101: data <= 32'h3a58b034;
    11'b01011101110: data <= 32'h38f2b26a;
    11'b01011101111: data <= 32'hbcceb7a5;
    11'b01011110000: data <= 32'hc13bbd4e;
    11'b01011110001: data <= 32'hbef3bec9;
    11'b01011110010: data <= 32'h35b9b9ed;
    11'b01011110011: data <= 32'h3cac3833;
    11'b01011110100: data <= 32'h32953929;
    11'b01011110101: data <= 32'hba692f1e;
    11'b01011110110: data <= 32'hba3238e0;
    11'b01011110111: data <= 32'hb8134024;
    11'b01011111000: data <= 32'hb9ec40bb;
    11'b01011111001: data <= 32'hb9e73819;
    11'b01011111010: data <= 32'h32b5be0e;
    11'b01011111011: data <= 32'h3d07bd8b;
    11'b01011111100: data <= 32'h3d2235d8;
    11'b01011111101: data <= 32'h3a873d3f;
    11'b01011111110: data <= 32'h3c6738f2;
    11'b01011111111: data <= 32'h3ef0b3f7;
    11'b01100000000: data <= 32'h3c2db2ac;
    11'b01100000001: data <= 32'hbc0fada3;
    11'b01100000010: data <= 32'hc05bba80;
    11'b01100000011: data <= 32'hbba9bea6;
    11'b01100000100: data <= 32'h3c2bbe1b;
    11'b01100000101: data <= 32'h3d2bba4d;
    11'b01100000110: data <= 32'hb211b80e;
    11'b01100000111: data <= 32'hbcd9b6c6;
    11'b01100001000: data <= 32'hba673849;
    11'b01100001001: data <= 32'hb4f43fc8;
    11'b01100001010: data <= 32'hbb0c3fbf;
    11'b01100001011: data <= 32'hbe622d69;
    11'b01100001100: data <= 32'hbc8abdc7;
    11'b01100001101: data <= 32'h2e1cb9df;
    11'b01100001110: data <= 32'h3a8e3c8c;
    11'b01100001111: data <= 32'h3bcf3ec7;
    11'b01100010000: data <= 32'h3d8038fe;
    11'b01100010001: data <= 32'h3effae22;
    11'b01100010010: data <= 32'h3b933856;
    11'b01100010011: data <= 32'hba1a3c75;
    11'b01100010100: data <= 32'hbd843232;
    11'b01100010101: data <= 32'h2668bda4;
    11'b01100010110: data <= 32'h3e96c002;
    11'b01100010111: data <= 32'h3d7fbdec;
    11'b01100011000: data <= 32'hb1fcbb8e;
    11'b01100011001: data <= 32'hba0eb8fa;
    11'b01100011010: data <= 32'h2e813195;
    11'b01100011011: data <= 32'h37193c9d;
    11'b01100011100: data <= 32'hbb173b9f;
    11'b01100011101: data <= 32'hc0cbb868;
    11'b01100011110: data <= 32'hc063bde0;
    11'b01100011111: data <= 32'hb945b7a6;
    11'b01100100000: data <= 32'h374f3c66;
    11'b01100100001: data <= 32'h39263cce;
    11'b01100100010: data <= 32'h3a003109;
    11'b01100100011: data <= 32'h3ba92f1d;
    11'b01100100100: data <= 32'h37773e3c;
    11'b01100100101: data <= 32'hb8ee40d6;
    11'b01100100110: data <= 32'hbaa13c7c;
    11'b01100100111: data <= 32'h36a3bc37;
    11'b01100101000: data <= 32'h3e4cbf80;
    11'b01100101001: data <= 32'h3ca9bcb0;
    11'b01100101010: data <= 32'h2e9db79d;
    11'b01100101011: data <= 32'h349cb687;
    11'b01100101100: data <= 32'h3dd8b27a;
    11'b01100101101: data <= 32'h3d8e355f;
    11'b01100101110: data <= 32'hb96b334f;
    11'b01100101111: data <= 32'hc138ba62;
    11'b01100110000: data <= 32'hc0a4bdaf;
    11'b01100110001: data <= 32'hb896b9b6;
    11'b01100110010: data <= 32'h366a3347;
    11'b01100110011: data <= 32'h2ceb0d89;
    11'b01100110100: data <= 32'hb3c0b93e;
    11'b01100110101: data <= 32'h2a3b3002;
    11'b01100110110: data <= 32'h2cdc4053;
    11'b01100110111: data <= 32'hb8954208;
    11'b01100111000: data <= 32'hbaff3da5;
    11'b01100111001: data <= 32'hb043ba7a;
    11'b01100111010: data <= 32'h398fbd07;
    11'b01100111011: data <= 32'h38cab144;
    11'b01100111100: data <= 32'h35a23731;
    11'b01100111101: data <= 32'h3cdfaa71;
    11'b01100111110: data <= 32'h40e7b672;
    11'b01100111111: data <= 32'h3feb2cc3;
    11'b01101000000: data <= 32'hb5d83602;
    11'b01101000001: data <= 32'hc040b4cb;
    11'b01101000010: data <= 32'hbe01bc85;
    11'b01101000011: data <= 32'h3268bc99;
    11'b01101000100: data <= 32'h38d1bb1d;
    11'b01101000101: data <= 32'hb603bcd7;
    11'b01101000110: data <= 32'hbaf9bd97;
    11'b01101000111: data <= 32'hb2c2affc;
    11'b01101001000: data <= 32'h339e3fe1;
    11'b01101001001: data <= 32'hb7b34123;
    11'b01101001010: data <= 32'hbd8a3b7c;
    11'b01101001011: data <= 32'hbd13ba5f;
    11'b01101001100: data <= 32'hb83ab882;
    11'b01101001101: data <= 32'haeff3a5c;
    11'b01101001110: data <= 32'h349b3c37;
    11'b01101001111: data <= 32'h3d9f2332;
    11'b01101010000: data <= 32'h40f2b732;
    11'b01101010001: data <= 32'h3f8537d7;
    11'b01101010010: data <= 32'hb0773d70;
    11'b01101010011: data <= 32'hbd2c3a1d;
    11'b01101010100: data <= 32'hb5bbb8e2;
    11'b01101010101: data <= 32'h3c0dbd73;
    11'b01101010110: data <= 32'h3a13bde5;
    11'b01101010111: data <= 32'hb851beb8;
    11'b01101011000: data <= 32'hb9ddbe98;
    11'b01101011001: data <= 32'h3772b7fc;
    11'b01101011010: data <= 32'h3c263c93;
    11'b01101011011: data <= 32'hb2ad3dce;
    11'b01101011100: data <= 32'hbf8f2f14;
    11'b01101011101: data <= 32'hc067bb46;
    11'b01101011110: data <= 32'hbd5ab182;
    11'b01101011111: data <= 32'hb8a43c36;
    11'b01101100000: data <= 32'haeb53a57;
    11'b01101100001: data <= 32'h39edb7af;
    11'b01101100010: data <= 32'h3e50b823;
    11'b01101100011: data <= 32'h3cf33cc5;
    11'b01101100100: data <= 32'had65410b;
    11'b01101100101: data <= 32'hb9123f0f;
    11'b01101100110: data <= 32'h34e8adf8;
    11'b01101100111: data <= 32'h3cb6bc7c;
    11'b01101101000: data <= 32'h385fbc77;
    11'b01101101001: data <= 32'hb815bc90;
    11'b01101101010: data <= 32'ha16bbd3d;
    11'b01101101011: data <= 32'h3eaeba56;
    11'b01101101100: data <= 32'h402233ad;
    11'b01101101101: data <= 32'h32923792;
    11'b01101101110: data <= 32'hbfc7b613;
    11'b01101101111: data <= 32'hc088bb11;
    11'b01101110000: data <= 32'hbcddb15d;
    11'b01101110001: data <= 32'hb87c380c;
    11'b01101110010: data <= 32'hb8e0b3be;
    11'b01101110011: data <= 32'hb529bd88;
    11'b01101110100: data <= 32'h3705b9ef;
    11'b01101110101: data <= 32'h38d13e62;
    11'b01101110110: data <= 32'hadc64217;
    11'b01101110111: data <= 32'hb770401b;
    11'b01101111000: data <= 32'h2d53302e;
    11'b01101111001: data <= 32'h37b2b844;
    11'b01101111010: data <= 32'haed7a9ff;
    11'b01101111011: data <= 32'hb82fa26b;
    11'b01101111100: data <= 32'h397eb9ba;
    11'b01101111101: data <= 32'h4129bb5e;
    11'b01101111110: data <= 32'h4161b2ab;
    11'b01101111111: data <= 32'h386e34ce;
    11'b01110000000: data <= 32'hbdccad55;
    11'b01110000001: data <= 32'hbd8db82b;
    11'b01110000010: data <= 32'hb452b549;
    11'b01110000011: data <= 32'hb095b5a1;
    11'b01110000100: data <= 32'hbbd5bd77;
    11'b01110000101: data <= 32'hbc73c061;
    11'b01110000110: data <= 32'hb042bc56;
    11'b01110000111: data <= 32'h38563d69;
    11'b01110001000: data <= 32'h2a354115;
    11'b01110001001: data <= 32'hb9a03dc2;
    11'b01110001010: data <= 32'hba2fa954;
    11'b01110001011: data <= 32'hb9292cff;
    11'b01110001100: data <= 32'hbb403c35;
    11'b01110001101: data <= 32'hb9dd3b25;
    11'b01110001110: data <= 32'h3a46b698;
    11'b01110001111: data <= 32'h4118bbe2;
    11'b01110010000: data <= 32'h40fcaafa;
    11'b01110010001: data <= 32'h39133bea;
    11'b01110010010: data <= 32'hb9813af1;
    11'b01110010011: data <= 32'hafba2ecf;
    11'b01110010100: data <= 32'h3aa4b5a4;
    11'b01110010101: data <= 32'h343dba78;
    11'b01110010110: data <= 32'hbc87bf24;
    11'b01110010111: data <= 32'hbce0c0c6;
    11'b01110011000: data <= 32'h3398bd73;
    11'b01110011001: data <= 32'h3cd438a0;
    11'b01110011010: data <= 32'h36e33d40;
    11'b01110011011: data <= 32'hbbdc357f;
    11'b01110011100: data <= 32'hbe2cb68c;
    11'b01110011101: data <= 32'hbda136f6;
    11'b01110011110: data <= 32'hbd7b3e27;
    11'b01110011111: data <= 32'hbc583b91;
    11'b01110100000: data <= 32'h30a9b9fd;
    11'b01110100001: data <= 32'h3e38bc9c;
    11'b01110100010: data <= 32'h3e693672;
    11'b01110100011: data <= 32'h370c3fd5;
    11'b01110100100: data <= 32'had1c3f48;
    11'b01110100101: data <= 32'h3a0e3947;
    11'b01110100110: data <= 32'h3d45add6;
    11'b01110100111: data <= 32'h338cb727;
    11'b01110101000: data <= 32'hbcbdbca7;
    11'b01110101001: data <= 32'hba02bf59;
    11'b01110101010: data <= 32'h3ce5bdb3;
    11'b01110101011: data <= 32'h405eb43e;
    11'b01110101100: data <= 32'h3b53305c;
    11'b01110101101: data <= 32'hbbb1b79c;
    11'b01110101110: data <= 32'hbe48b8c1;
    11'b01110101111: data <= 32'hbcdf37fd;
    11'b01110110000: data <= 32'hbcbc3cff;
    11'b01110110001: data <= 32'hbd9130db;
    11'b01110110010: data <= 32'hbadabe5b;
    11'b01110110011: data <= 32'h336cbde4;
    11'b01110110100: data <= 32'h391a3977;
    11'b01110110101: data <= 32'h325b40d4;
    11'b01110110110: data <= 32'h2ff0401c;
    11'b01110110111: data <= 32'h3a553a22;
    11'b01110111000: data <= 32'h3b113578;
    11'b01110111001: data <= 32'hb5693890;
    11'b01110111010: data <= 32'hbd3a303b;
    11'b01110111011: data <= 32'hb2e1bb5f;
    11'b01110111100: data <= 32'h4014bd33;
    11'b01110111101: data <= 32'h4189b9c8;
    11'b01110111110: data <= 32'h3ccbb4ac;
    11'b01110111111: data <= 32'hb893b778;
    11'b01111000000: data <= 32'hb9d2b562;
    11'b01111000001: data <= 32'hafd73733;
    11'b01111000010: data <= 32'hb76a38aa;
    11'b01111000011: data <= 32'hbe02bad1;
    11'b01111000100: data <= 32'hbe8bc0bc;
    11'b01111000101: data <= 32'hb8b8bf32;
    11'b01111000110: data <= 32'h344137e3;
    11'b01111000111: data <= 32'h32693fb5;
    11'b01111001000: data <= 32'ha0283d3f;
    11'b01111001001: data <= 32'h30d43523;
    11'b01111001010: data <= 32'hae2f39a1;
    11'b01111001011: data <= 32'hbc783e95;
    11'b01111001100: data <= 32'hbe2d3d1f;
    11'b01111001101: data <= 32'haf5cb492;
    11'b01111001110: data <= 32'h4002bcc5;
    11'b01111001111: data <= 32'h40edb945;
    11'b01111010000: data <= 32'h3c2d3137;
    11'b01111010001: data <= 32'ha8de34f0;
    11'b01111010010: data <= 32'h3817344c;
    11'b01111010011: data <= 32'h3cd937e0;
    11'b01111010100: data <= 32'h34a13179;
    11'b01111010101: data <= 32'hbdcfbd03;
    11'b01111010110: data <= 32'hbf3ec0f8;
    11'b01111010111: data <= 32'hb776bf8e;
    11'b01111011000: data <= 32'h39c9ad5e;
    11'b01111011001: data <= 32'h385e39cc;
    11'b01111011010: data <= 32'hb254a0d3;
    11'b01111011011: data <= 32'hb83fb655;
    11'b01111011100: data <= 32'hba963aad;
    11'b01111011101: data <= 32'hbe1e405d;
    11'b01111011110: data <= 32'hbf0d3e5c;
    11'b01111011111: data <= 32'hb8bfb619;
    11'b01111100000: data <= 32'h3c24bd32;
    11'b01111100001: data <= 32'h3d74b4dc;
    11'b01111100010: data <= 32'h380b3c06;
    11'b01111100011: data <= 32'h35483cd2;
    11'b01111100100: data <= 32'h3db33a5c;
    11'b01111100101: data <= 32'h3fdd3962;
    11'b01111100110: data <= 32'h384636a4;
    11'b01111100111: data <= 32'hbda9b935;
    11'b01111101000: data <= 32'hbdcabeff;
    11'b01111101001: data <= 32'h35d4be7f;
    11'b01111101010: data <= 32'h3e7bb978;
    11'b01111101011: data <= 32'h3c14b7a7;
    11'b01111101100: data <= 32'hb29cbc69;
    11'b01111101101: data <= 32'hb90bbb18;
    11'b01111101110: data <= 32'hb9303a36;
    11'b01111101111: data <= 32'hbcc03ff9;
    11'b01111110000: data <= 32'hbf183bd2;
    11'b01111110001: data <= 32'hbd6fbc74;
    11'b01111110010: data <= 32'hb4e2be74;
    11'b01111110011: data <= 32'h2faba867;
    11'b01111110100: data <= 32'hac8c3df8;
    11'b01111110101: data <= 32'h36123dcc;
    11'b01111110110: data <= 32'h3e363a41;
    11'b01111110111: data <= 32'h3ef53ad8;
    11'b01111111000: data <= 32'h2e6a3cdb;
    11'b01111111001: data <= 32'hbe1c393d;
    11'b01111111010: data <= 32'hbba1b875;
    11'b01111111011: data <= 32'h3caebc94;
    11'b01111111100: data <= 32'h4069bba9;
    11'b01111111101: data <= 32'h3cdebbf1;
    11'b01111111110: data <= 32'ha48fbd50;
    11'b01111111111: data <= 32'h254eba75;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    