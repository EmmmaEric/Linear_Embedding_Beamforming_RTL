
module memory_rom_34(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbd93ba03;
    11'b00000000001: data <= 32'hba75b600;
    11'b00000000010: data <= 32'h3a7437ac;
    11'b00000000011: data <= 32'h3c3e3e2d;
    11'b00000000100: data <= 32'hb98b3e54;
    11'b00000000101: data <= 32'hc097382f;
    11'b00000000110: data <= 32'hbf5aad75;
    11'b00000000111: data <= 32'hb0583845;
    11'b00000001000: data <= 32'h3b023c21;
    11'b00000001001: data <= 32'h3b742fe9;
    11'b00000001010: data <= 32'h3c75bc46;
    11'b00000001011: data <= 32'h3e42b831;
    11'b00000001100: data <= 32'h3d3b3d9d;
    11'b00000001101: data <= 32'h34534049;
    11'b00000001110: data <= 32'hb4c1381d;
    11'b00000001111: data <= 32'h2efdbe80;
    11'b00000010000: data <= 32'h3547c02e;
    11'b00000010001: data <= 32'hb6babce7;
    11'b00000010010: data <= 32'hbba8ba1d;
    11'b00000010011: data <= 32'h27dbbbef;
    11'b00000010100: data <= 32'h3de7b9d8;
    11'b00000010101: data <= 32'h3c6134a4;
    11'b00000010110: data <= 32'hbcb83b36;
    11'b00000010111: data <= 32'hc1983859;
    11'b00000011000: data <= 32'hc02331a0;
    11'b00000011001: data <= 32'hb5843780;
    11'b00000011010: data <= 32'h3347386c;
    11'b00000011011: data <= 32'hb387b4bc;
    11'b00000011100: data <= 32'hacf4bb42;
    11'b00000011101: data <= 32'h3be2334a;
    11'b00000011110: data <= 32'h3e1a4080;
    11'b00000011111: data <= 32'h3ae2414e;
    11'b00000100000: data <= 32'h2b123a4b;
    11'b00000100001: data <= 32'h24f1bc85;
    11'b00000100010: data <= 32'h3154bcaa;
    11'b00000100011: data <= 32'hb023b419;
    11'b00000100100: data <= 32'hae32b65c;
    11'b00000100101: data <= 32'h3c21bdf0;
    11'b00000100110: data <= 32'h4037bebb;
    11'b00000100111: data <= 32'h3d35b73e;
    11'b00000101000: data <= 32'hbbe2396b;
    11'b00000101001: data <= 32'hc0903860;
    11'b00000101010: data <= 32'hbdcaafd3;
    11'b00000101011: data <= 32'hb352b539;
    11'b00000101100: data <= 32'hb80ab64e;
    11'b00000101101: data <= 32'hbdeebaf0;
    11'b00000101110: data <= 32'hbc79bb80;
    11'b00000101111: data <= 32'h38a23666;
    11'b00000110000: data <= 32'h3e23406b;
    11'b00000110001: data <= 32'h39c940df;
    11'b00000110010: data <= 32'hb81c3b30;
    11'b00000110011: data <= 32'hb9b1b477;
    11'b00000110100: data <= 32'hb29332b8;
    11'b00000110101: data <= 32'h2d953b6b;
    11'b00000110110: data <= 32'h36e529df;
    11'b00000110111: data <= 32'h3dabbea0;
    11'b00000111000: data <= 32'h407bbf7c;
    11'b00000111001: data <= 32'h3e3eb3ca;
    11'b00000111010: data <= 32'hb17e3c70;
    11'b00000111011: data <= 32'hbbf03973;
    11'b00000111100: data <= 32'hb523b89c;
    11'b00000111101: data <= 32'h2f76bc89;
    11'b00000111110: data <= 32'hbb7fbc49;
    11'b00000111111: data <= 32'hc02fbcd1;
    11'b00001000000: data <= 32'hbd61bcd4;
    11'b00001000001: data <= 32'h399db32a;
    11'b00001000010: data <= 32'h3dfa3ccb;
    11'b00001000011: data <= 32'h30913e36;
    11'b00001000100: data <= 32'hbddc3a15;
    11'b00001000101: data <= 32'hbe1336e3;
    11'b00001000110: data <= 32'hb8883ce0;
    11'b00001000111: data <= 32'ha7a93e47;
    11'b00001001000: data <= 32'h300b31d9;
    11'b00001001001: data <= 32'h3a63be46;
    11'b00001001010: data <= 32'h3ed1bd67;
    11'b00001001011: data <= 32'h3eb8394b;
    11'b00001001100: data <= 32'h3a253f8a;
    11'b00001001101: data <= 32'h34b43b64;
    11'b00001001110: data <= 32'h38dbb9e8;
    11'b00001001111: data <= 32'h366abcf3;
    11'b00001010000: data <= 32'hbb7fbb05;
    11'b00001010001: data <= 32'hbf49bc05;
    11'b00001010010: data <= 32'hb981be27;
    11'b00001010011: data <= 32'h3d35bd28;
    11'b00001010100: data <= 32'h3e34b22c;
    11'b00001010101: data <= 32'hb5403848;
    11'b00001010110: data <= 32'hbff037d7;
    11'b00001010111: data <= 32'hbedc3920;
    11'b00001011000: data <= 32'hb8dc3d4e;
    11'b00001011001: data <= 32'hb6ec3d37;
    11'b00001011010: data <= 32'hbb3db08f;
    11'b00001011011: data <= 32'hb829bdc0;
    11'b00001011100: data <= 32'h3a4bb936;
    11'b00001011101: data <= 32'h3e553dfd;
    11'b00001011110: data <= 32'h3d2240be;
    11'b00001011111: data <= 32'h3a993c4b;
    11'b00001100000: data <= 32'h3a22b71a;
    11'b00001100001: data <= 32'h35dab6ea;
    11'b00001100010: data <= 32'hb96a3293;
    11'b00001100011: data <= 32'hbc2eb4fd;
    11'b00001100100: data <= 32'h3461bed2;
    11'b00001100101: data <= 32'h3fabc04b;
    11'b00001100110: data <= 32'h3eb6bc78;
    11'b00001100111: data <= 32'hb49526a8;
    11'b00001101000: data <= 32'hbe463532;
    11'b00001101001: data <= 32'hbbf735d3;
    11'b00001101010: data <= 32'hb2033925;
    11'b00001101011: data <= 32'hbac036de;
    11'b00001101100: data <= 32'hc018b996;
    11'b00001101101: data <= 32'hbef9bdb6;
    11'b00001101110: data <= 32'h2c2eb5f4;
    11'b00001101111: data <= 32'h3d863e2a;
    11'b00001110000: data <= 32'h3c994026;
    11'b00001110001: data <= 32'h36403b4f;
    11'b00001110010: data <= 32'h309f2e89;
    11'b00001110011: data <= 32'h24b53aae;
    11'b00001110100: data <= 32'hb7373e48;
    11'b00001110101: data <= 32'hb7453783;
    11'b00001110110: data <= 32'h39d1be84;
    11'b00001110111: data <= 32'h3ffac0a4;
    11'b00001111000: data <= 32'h3ed1bc3f;
    11'b00001111001: data <= 32'h33e334f0;
    11'b00001111010: data <= 32'hb6373699;
    11'b00001111011: data <= 32'h34efad11;
    11'b00001111100: data <= 32'h3812b1fc;
    11'b00001111101: data <= 32'hbbfdb4c6;
    11'b00001111110: data <= 32'hc13fbc04;
    11'b00001111111: data <= 32'hc048be0c;
    11'b00010000000: data <= 32'h9cfdb9fa;
    11'b00010000001: data <= 32'h3d0d3917;
    11'b00010000010: data <= 32'h38b63c18;
    11'b00010000011: data <= 32'hb85f36bd;
    11'b00010000100: data <= 32'hb983381f;
    11'b00010000101: data <= 32'hb5473f31;
    11'b00010000110: data <= 32'hb6e240cd;
    11'b00010000111: data <= 32'hb85e3abe;
    11'b00010001000: data <= 32'h32ccbdb4;
    11'b00010001001: data <= 32'h3d3dbf45;
    11'b00010001010: data <= 32'h3debb27f;
    11'b00010001011: data <= 32'h3b0b3c54;
    11'b00010001100: data <= 32'h3abf3936;
    11'b00010001101: data <= 32'h3dc3b561;
    11'b00010001110: data <= 32'h3c49b76a;
    11'b00010001111: data <= 32'hbac1b294;
    11'b00010010000: data <= 32'hc0bbb977;
    11'b00010010001: data <= 32'hbe3ebe17;
    11'b00010010010: data <= 32'h387abe08;
    11'b00010010011: data <= 32'h3d41b98b;
    11'b00010010100: data <= 32'h2b56b2ba;
    11'b00010010101: data <= 32'hbccdb14a;
    11'b00010010110: data <= 32'hbbd93844;
    11'b00010010111: data <= 32'hb47b3fa8;
    11'b00010011000: data <= 32'hb863407d;
    11'b00010011001: data <= 32'hbd2438bd;
    11'b00010011010: data <= 32'hbc25bd1c;
    11'b00010011011: data <= 32'h3187bc55;
    11'b00010011100: data <= 32'h3c2839dd;
    11'b00010011101: data <= 32'h3cad3ea0;
    11'b00010011110: data <= 32'h3d8139eb;
    11'b00010011111: data <= 32'h3ef9b48c;
    11'b00010100000: data <= 32'h3ca22c74;
    11'b00010100001: data <= 32'hb85f3a69;
    11'b00010100010: data <= 32'hbe4a3316;
    11'b00010100011: data <= 32'hb840bd52;
    11'b00010100100: data <= 32'h3d02c039;
    11'b00010100101: data <= 32'h3d9fbe73;
    11'b00010100110: data <= 32'hae8abb29;
    11'b00010100111: data <= 32'hbc22b809;
    11'b00010101000: data <= 32'hb5813211;
    11'b00010101001: data <= 32'h35573ce8;
    11'b00010101010: data <= 32'hb8d03d58;
    11'b00010101011: data <= 32'hc050a5f1;
    11'b00010101100: data <= 32'hc080bd01;
    11'b00010101101: data <= 32'hba06b922;
    11'b00010101110: data <= 32'h38e03c00;
    11'b00010101111: data <= 32'h3b773dcb;
    11'b00010110000: data <= 32'h3b93368d;
    11'b00010110001: data <= 32'h3c82ad48;
    11'b00010110010: data <= 32'h3a3a3c3e;
    11'b00010110011: data <= 32'hb50c404d;
    11'b00010110100: data <= 32'hbad63cea;
    11'b00010110101: data <= 32'h2fcdbbda;
    11'b00010110110: data <= 32'h3db6c04a;
    11'b00010110111: data <= 32'h3d2bbe45;
    11'b00010111000: data <= 32'h2ef8b94b;
    11'b00010111001: data <= 32'hb018b6c5;
    11'b00010111010: data <= 32'h3b84b425;
    11'b00010111011: data <= 32'h3d1434d2;
    11'b00010111100: data <= 32'hb72b36f5;
    11'b00010111101: data <= 32'hc11fb6f7;
    11'b00010111110: data <= 32'hc153bcea;
    11'b00010111111: data <= 32'hbb53b9c9;
    11'b00011000000: data <= 32'h370235dc;
    11'b00011000001: data <= 32'h35a736d3;
    11'b00011000010: data <= 32'hab8ab537;
    11'b00011000011: data <= 32'h30cb99a4;
    11'b00011000100: data <= 32'h35253f4f;
    11'b00011000101: data <= 32'hb31c4200;
    11'b00011000110: data <= 32'hb97f3ef2;
    11'b00011000111: data <= 32'hb01fb961;
    11'b00011001000: data <= 32'h3a4abe69;
    11'b00011001001: data <= 32'h3aa7b949;
    11'b00011001010: data <= 32'h36553313;
    11'b00011001011: data <= 32'h3b1cad67;
    11'b00011001100: data <= 32'h4032b87d;
    11'b00011001101: data <= 32'h4004b263;
    11'b00011001110: data <= 32'hb053345d;
    11'b00011001111: data <= 32'hc079b1ac;
    11'b00011010000: data <= 32'hc019bc19;
    11'b00011010001: data <= 32'hb47dbc8a;
    11'b00011010010: data <= 32'h388bb9de;
    11'b00011010011: data <= 32'hb29cbab2;
    11'b00011010100: data <= 32'hbb3dbc80;
    11'b00011010101: data <= 32'hb625b22e;
    11'b00011010110: data <= 32'h349c3f68;
    11'b00011010111: data <= 32'hb0f541a9;
    11'b00011011000: data <= 32'hbc583dd7;
    11'b00011011001: data <= 32'hbc8cb897;
    11'b00011011010: data <= 32'hb60abac4;
    11'b00011011011: data <= 32'h30cb3704;
    11'b00011011100: data <= 32'h36e63c16;
    11'b00011011101: data <= 32'h3d392ea5;
    11'b00011011110: data <= 32'h40d0b94a;
    11'b00011011111: data <= 32'h403c2244;
    11'b00011100000: data <= 32'h30e43c20;
    11'b00011100001: data <= 32'hbdae39f3;
    11'b00011100010: data <= 32'hbb10b89f;
    11'b00011100011: data <= 32'h38f4bdcc;
    11'b00011100100: data <= 32'h3a29be0f;
    11'b00011100101: data <= 32'hb7c8be32;
    11'b00011100110: data <= 32'hbc25be2a;
    11'b00011100111: data <= 32'h8813b897;
    11'b00011101000: data <= 32'h3b363c86;
    11'b00011101001: data <= 32'h29f33f3f;
    11'b00011101010: data <= 32'hbe943949;
    11'b00011101011: data <= 32'hc062b94a;
    11'b00011101100: data <= 32'hbd64b4f8;
    11'b00011101101: data <= 32'hb68d3bdc;
    11'b00011101110: data <= 32'h2ec63c48;
    11'b00011101111: data <= 32'h3aa7b28a;
    11'b00011110000: data <= 32'h3ed5b99e;
    11'b00011110001: data <= 32'h3e5b396e;
    11'b00011110010: data <= 32'h346a4069;
    11'b00011110011: data <= 32'hb90a3f39;
    11'b00011110100: data <= 32'h26a8aaa3;
    11'b00011110101: data <= 32'h3c38bd5e;
    11'b00011110110: data <= 32'h39a0bda3;
    11'b00011110111: data <= 32'hb7f9bd0d;
    11'b00011111000: data <= 32'hb753bd6d;
    11'b00011111001: data <= 32'h3c61bb79;
    11'b00011111010: data <= 32'h3f9730c8;
    11'b00011111011: data <= 32'h369e3968;
    11'b00011111100: data <= 32'hbf72a270;
    11'b00011111101: data <= 32'hc10db9b0;
    11'b00011111110: data <= 32'hbdf4b232;
    11'b00011111111: data <= 32'hb8403962;
    11'b00100000000: data <= 32'hb6ad3405;
    11'b00100000001: data <= 32'hb321bbf9;
    11'b00100000010: data <= 32'h382cbae2;
    11'b00100000011: data <= 32'h3b033ce1;
    11'b00100000100: data <= 32'h346341ee;
    11'b00100000101: data <= 32'hb4a740a5;
    11'b00100000110: data <= 32'h2e1f343c;
    11'b00100000111: data <= 32'h3910ba83;
    11'b00100001000: data <= 32'h3259b746;
    11'b00100001001: data <= 32'hb767b266;
    11'b00100001010: data <= 32'h34dfba3b;
    11'b00100001011: data <= 32'h404dbc82;
    11'b00100001100: data <= 32'h4158b7ef;
    11'b00100001101: data <= 32'h3a523271;
    11'b00100001110: data <= 32'hbe081ef6;
    11'b00100001111: data <= 32'hbf75b7bd;
    11'b00100010000: data <= 32'hb9a3b5a1;
    11'b00100010001: data <= 32'hb21eb0c9;
    11'b00100010010: data <= 32'hbaeebb2e;
    11'b00100010011: data <= 32'hbcc3bf6e;
    11'b00100010100: data <= 32'hb505bcab;
    11'b00100010101: data <= 32'h38b13cae;
    11'b00100010110: data <= 32'h355f417b;
    11'b00100010111: data <= 32'hb71e3fb9;
    11'b00100011000: data <= 32'hb8f23225;
    11'b00100011001: data <= 32'hb66ab107;
    11'b00100011010: data <= 32'hb87f39ff;
    11'b00100011011: data <= 32'hb8ba3b1c;
    11'b00100011100: data <= 32'h38dab522;
    11'b00100011101: data <= 32'h40cfbcc3;
    11'b00100011110: data <= 32'h416ab81a;
    11'b00100011111: data <= 32'h3ba1393a;
    11'b00100100000: data <= 32'hba273a38;
    11'b00100100001: data <= 32'hb8d22a09;
    11'b00100100010: data <= 32'h3778b771;
    11'b00100100011: data <= 32'h3490ba39;
    11'b00100100100: data <= 32'hbc56be38;
    11'b00100100101: data <= 32'hbe1fc07b;
    11'b00100100110: data <= 32'hb3d3bdea;
    11'b00100100111: data <= 32'h3c193804;
    11'b00100101000: data <= 32'h38e83e8a;
    11'b00100101001: data <= 32'hba393b0e;
    11'b00100101010: data <= 32'hbdf1b14f;
    11'b00100101011: data <= 32'hbd4034c6;
    11'b00100101100: data <= 32'hbc873df1;
    11'b00100101101: data <= 32'hbb3e3d08;
    11'b00100101110: data <= 32'h30ddb6da;
    11'b00100101111: data <= 32'h3e84bd29;
    11'b00100110000: data <= 32'h3fd4ad59;
    11'b00100110001: data <= 32'h3a923e73;
    11'b00100110010: data <= 32'hac6a3f18;
    11'b00100110011: data <= 32'h37ba38f4;
    11'b00100110100: data <= 32'h3ce9b4f4;
    11'b00100110101: data <= 32'h3721b93f;
    11'b00100110110: data <= 32'hbc86bccf;
    11'b00100110111: data <= 32'hbcc5bf7f;
    11'b00100111000: data <= 32'h38e4be71;
    11'b00100111001: data <= 32'h3fc5b638;
    11'b00100111010: data <= 32'h3c353564;
    11'b00100111011: data <= 32'hbb29afa3;
    11'b00100111100: data <= 32'hbf12b77b;
    11'b00100111101: data <= 32'hbd9836cb;
    11'b00100111110: data <= 32'hbc793da8;
    11'b00100111111: data <= 32'hbcf73998;
    11'b00101000000: data <= 32'hba8ebc80;
    11'b00101000001: data <= 32'h34b5be22;
    11'b00101000010: data <= 32'h3b5e3514;
    11'b00101000011: data <= 32'h38624092;
    11'b00101000100: data <= 32'h340f407d;
    11'b00101000101: data <= 32'h3a4c3acb;
    11'b00101000110: data <= 32'h3c5b2d3f;
    11'b00101000111: data <= 32'h2ba23370;
    11'b00101001000: data <= 32'hbcbd9ef3;
    11'b00101001001: data <= 32'hb8d1bbe8;
    11'b00101001010: data <= 32'h3e36be17;
    11'b00101001011: data <= 32'h415cbbf5;
    11'b00101001100: data <= 32'h3d8eb5e0;
    11'b00101001101: data <= 32'hb8fdb682;
    11'b00101001110: data <= 32'hbc99b63d;
    11'b00101001111: data <= 32'hb7f63597;
    11'b00101010000: data <= 32'hb7ee3a4d;
    11'b00101010001: data <= 32'hbda8b4ee;
    11'b00101010010: data <= 32'hbeedbfd0;
    11'b00101010011: data <= 32'hba1bbf61;
    11'b00101010100: data <= 32'h34d934bf;
    11'b00101010101: data <= 32'h36cb4029;
    11'b00101010110: data <= 32'h315c3f04;
    11'b00101010111: data <= 32'h349c383c;
    11'b00101011000: data <= 32'h333537b4;
    11'b00101011001: data <= 32'hb9553d80;
    11'b00101011010: data <= 32'hbd6a3d2d;
    11'b00101011011: data <= 32'hb51eb201;
    11'b00101011100: data <= 32'h3f37bd78;
    11'b00101011101: data <= 32'h4145bc3b;
    11'b00101011110: data <= 32'h3d65b091;
    11'b00101011111: data <= 32'haf2e312c;
    11'b00101100000: data <= 32'h2ac32e0b;
    11'b00101100001: data <= 32'h3b0434dc;
    11'b00101100010: data <= 32'h3548332e;
    11'b00101100011: data <= 32'hbd8bbb89;
    11'b00101100100: data <= 32'hc031c090;
    11'b00101100101: data <= 32'hbb70c000;
    11'b00101100110: data <= 32'h380bb1d1;
    11'b00101100111: data <= 32'h390e3c1d;
    11'b00101101000: data <= 32'had51381b;
    11'b00101101001: data <= 32'hb798b198;
    11'b00101101010: data <= 32'hb9203964;
    11'b00101101011: data <= 32'hbcd0403b;
    11'b00101101100: data <= 32'hbe433fa0;
    11'b00101101101: data <= 32'hb905a69f;
    11'b00101101110: data <= 32'h3c4cbd76;
    11'b00101101111: data <= 32'h3ed9b9b4;
    11'b00101110000: data <= 32'h3b10396e;
    11'b00101110001: data <= 32'h351b3c58;
    11'b00101110010: data <= 32'h3c863930;
    11'b00101110011: data <= 32'h3f8c3686;
    11'b00101110100: data <= 32'h3a5433dd;
    11'b00101110101: data <= 32'hbd30b906;
    11'b00101110110: data <= 32'hbf57bf10;
    11'b00101110111: data <= 32'hb39ebf4e;
    11'b00101111000: data <= 32'h3d49ba77;
    11'b00101111001: data <= 32'h3c3bb411;
    11'b00101111010: data <= 32'hb2abb9ef;
    11'b00101111011: data <= 32'hba7dba73;
    11'b00101111100: data <= 32'hba0a390a;
    11'b00101111101: data <= 32'hbc49403a;
    11'b00101111110: data <= 32'hbe893e24;
    11'b00101111111: data <= 32'hbd66b8b6;
    11'b00110000000: data <= 32'hb3a5be5c;
    11'b00110000001: data <= 32'h36c2b563;
    11'b00110000010: data <= 32'h341d3d74;
    11'b00110000011: data <= 32'h370c3e4c;
    11'b00110000100: data <= 32'h3df93a59;
    11'b00110000101: data <= 32'h3fd638a4;
    11'b00110000110: data <= 32'h389a3b4a;
    11'b00110000111: data <= 32'hbd453857;
    11'b00110001000: data <= 32'hbd2ab915;
    11'b00110001001: data <= 32'h396bbd7e;
    11'b00110001010: data <= 32'h4020bcbf;
    11'b00110001011: data <= 32'h3d5bbc06;
    11'b00110001100: data <= 32'haebbbd0f;
    11'b00110001101: data <= 32'hb61ebb86;
    11'b00110001110: data <= 32'h2f8e37fd;
    11'b00110001111: data <= 32'hb3213e31;
    11'b00110010000: data <= 32'hbdc838b3;
    11'b00110010001: data <= 32'hc009bd9f;
    11'b00110010010: data <= 32'hbd57bf7b;
    11'b00110010011: data <= 32'hb741b39a;
    11'b00110010100: data <= 32'hafd63d41;
    11'b00110010101: data <= 32'h34493c73;
    11'b00110010110: data <= 32'h3c41345f;
    11'b00110010111: data <= 32'h3cc13918;
    11'b00110011000: data <= 32'haf853f39;
    11'b00110011001: data <= 32'hbde43f7f;
    11'b00110011010: data <= 32'hbb783707;
    11'b00110011011: data <= 32'h3c33bb5d;
    11'b00110011100: data <= 32'h4019bc84;
    11'b00110011101: data <= 32'h3c84bad9;
    11'b00110011110: data <= 32'h2df3ba9c;
    11'b00110011111: data <= 32'h38a1b828;
    11'b00110100000: data <= 32'h3e113726;
    11'b00110100001: data <= 32'h3b153b93;
    11'b00110100010: data <= 32'hbc59b04e;
    11'b00110100011: data <= 32'hc075bf13;
    11'b00110100100: data <= 32'hbe4dbf91;
    11'b00110100101: data <= 32'hb6b0b709;
    11'b00110100110: data <= 32'ha4c337d2;
    11'b00110100111: data <= 32'h1decb0b4;
    11'b00110101000: data <= 32'h34bcb9b6;
    11'b00110101001: data <= 32'h344a37a5;
    11'b00110101010: data <= 32'hb98740bb;
    11'b00110101011: data <= 32'hbe5a411e;
    11'b00110101100: data <= 32'hbc073a6f;
    11'b00110101101: data <= 32'h383fba25;
    11'b00110101110: data <= 32'h3c76ba0c;
    11'b00110101111: data <= 32'h363eaadc;
    11'b00110110000: data <= 32'h313e2f87;
    11'b00110110001: data <= 32'h3dd62c47;
    11'b00110110010: data <= 32'h413337d4;
    11'b00110110011: data <= 32'h3e553a3a;
    11'b00110110100: data <= 32'hba66a2a6;
    11'b00110110101: data <= 32'hbfa9bd05;
    11'b00110110110: data <= 32'hbb5ebdda;
    11'b00110110111: data <= 32'h3614b9ab;
    11'b00110111000: data <= 32'h36c8b8b0;
    11'b00110111001: data <= 32'hb0f3bde9;
    11'b00110111010: data <= 32'hb1f8be73;
    11'b00110111011: data <= 32'ha47a3219;
    11'b00110111100: data <= 32'hb8a04091;
    11'b00110111101: data <= 32'hbdbc407a;
    11'b00110111110: data <= 32'hbd8c34ca;
    11'b00110111111: data <= 32'hb88ebbe1;
    11'b00111000000: data <= 32'hb3f4b5be;
    11'b00111000001: data <= 32'hb83739e7;
    11'b00111000010: data <= 32'h14f73a06;
    11'b00111000011: data <= 32'h3ede33dc;
    11'b00111000100: data <= 32'h417a37a2;
    11'b00111000101: data <= 32'h3ddf3c82;
    11'b00111000110: data <= 32'hba393b8d;
    11'b00111000111: data <= 32'hbd6aab3b;
    11'b00111001000: data <= 32'h2c66b9a4;
    11'b00111001001: data <= 32'h3cf9ba2a;
    11'b00111001010: data <= 32'h3a00bcd9;
    11'b00111001011: data <= 32'hb248c029;
    11'b00111001100: data <= 32'ha92fbf93;
    11'b00111001101: data <= 32'h392ba646;
    11'b00111001110: data <= 32'h35353ec8;
    11'b00111001111: data <= 32'hbb853cfb;
    11'b00111010000: data <= 32'hbeddb8e4;
    11'b00111010001: data <= 32'hbe15bd41;
    11'b00111010010: data <= 32'hbce1b0d1;
    11'b00111010011: data <= 32'hbc683b7b;
    11'b00111010100: data <= 32'hb4d637e7;
    11'b00111010101: data <= 32'h3d04b4fa;
    11'b00111010110: data <= 32'h3fcc33c6;
    11'b00111010111: data <= 32'h39b43eb3;
    11'b00111011000: data <= 32'hbbd4403b;
    11'b00111011001: data <= 32'hbb533c7f;
    11'b00111011010: data <= 32'h393ca24b;
    11'b00111011011: data <= 32'h3db3b841;
    11'b00111011100: data <= 32'h3833bc0d;
    11'b00111011101: data <= 32'hb43abe9c;
    11'b00111011110: data <= 32'h389fbdcd;
    11'b00111011111: data <= 32'h3f80a9af;
    11'b00111100000: data <= 32'h3e2d3c26;
    11'b00111100001: data <= 32'hb4e43575;
    11'b00111100010: data <= 32'hbecbbca6;
    11'b00111100011: data <= 32'hbec7bd5e;
    11'b00111100100: data <= 32'hbce4af86;
    11'b00111100101: data <= 32'hbc193709;
    11'b00111100110: data <= 32'hb876b8b7;
    11'b00111100111: data <= 32'h3717bda1;
    11'b00111101000: data <= 32'h3b05b2e3;
    11'b00111101001: data <= 32'ha8ba3fe1;
    11'b00111101010: data <= 32'hbc7e416f;
    11'b00111101011: data <= 32'hba4e3e38;
    11'b00111101100: data <= 32'h372a3313;
    11'b00111101101: data <= 32'h3960b01d;
    11'b00111101110: data <= 32'hb50ab193;
    11'b00111101111: data <= 32'hb807b8b8;
    11'b00111110000: data <= 32'h3caab9a5;
    11'b00111110001: data <= 32'h41ba29ca;
    11'b00111110010: data <= 32'h40aa399f;
    11'b00111110011: data <= 32'h2f7d3171;
    11'b00111110100: data <= 32'hbd3fbab4;
    11'b00111110101: data <= 32'hbc02baa3;
    11'b00111110110: data <= 32'hb56faced;
    11'b00111110111: data <= 32'hb73bb538;
    11'b00111111000: data <= 32'hb94ebf42;
    11'b00111111001: data <= 32'hb185c0d6;
    11'b00111111010: data <= 32'h3525b983;
    11'b00111111011: data <= 32'hafd33f12;
    11'b00111111100: data <= 32'hbb4740b5;
    11'b00111111101: data <= 32'hbaf63bfd;
    11'b00111111110: data <= 32'hb559ada6;
    11'b00111111111: data <= 32'hb89f3304;
    11'b01000000000: data <= 32'hbd7539ca;
    11'b01000000001: data <= 32'hbb3034a9;
    11'b01000000010: data <= 32'h3d0db528;
    11'b01000000011: data <= 32'h41e71bb7;
    11'b01000000100: data <= 32'h40683a35;
    11'b01000000101: data <= 32'h2de63a71;
    11'b01000000110: data <= 32'hba403382;
    11'b01000000111: data <= 32'h2cd92c72;
    11'b01000001000: data <= 32'h39f3302e;
    11'b01000001001: data <= 32'h2d12ba08;
    11'b01000001010: data <= 32'hb9a3c0bc;
    11'b01000001011: data <= 32'hb45fc173;
    11'b01000001100: data <= 32'h3954bb46;
    11'b01000001101: data <= 32'h391d3cbd;
    11'b01000001110: data <= 32'hb4723d22;
    11'b01000001111: data <= 32'hbb3daeb7;
    11'b01000010000: data <= 32'hbc37b8e9;
    11'b01000010001: data <= 32'hbdfc367c;
    11'b01000010010: data <= 32'hc0023c8d;
    11'b01000010011: data <= 32'hbd0e3581;
    11'b01000010100: data <= 32'h3a30b9c1;
    11'b01000010101: data <= 32'h4031b5a7;
    11'b01000010110: data <= 32'h3d243c12;
    11'b01000010111: data <= 32'hb4a13ee2;
    11'b01000011000: data <= 32'hb6113d6e;
    11'b01000011001: data <= 32'h3ad13aeb;
    11'b01000011010: data <= 32'h3ce937d4;
    11'b01000011011: data <= 32'h2809b7df;
    11'b01000011100: data <= 32'hbafbbf86;
    11'b01000011101: data <= 32'h295ac050;
    11'b01000011110: data <= 32'h3e7bba32;
    11'b01000011111: data <= 32'h3f2c3889;
    11'b01000100000: data <= 32'h37cd32c2;
    11'b01000100001: data <= 32'hb9b6bb96;
    11'b01000100010: data <= 32'hbc83bab3;
    11'b01000100011: data <= 32'hbdce3816;
    11'b01000100100: data <= 32'hbf633b7b;
    11'b01000100101: data <= 32'hbd9cb73e;
    11'b01000100110: data <= 32'h95c9bef4;
    11'b01000100111: data <= 32'h3b01bbae;
    11'b01000101000: data <= 32'h34133c60;
    11'b01000101001: data <= 32'hb923405f;
    11'b01000101010: data <= 32'hb29c3eff;
    11'b01000101011: data <= 32'h3b623c44;
    11'b01000101100: data <= 32'h3a2b3a9c;
    11'b01000101101: data <= 32'hb9bb3531;
    11'b01000101110: data <= 32'hbd10b983;
    11'b01000101111: data <= 32'h3613bc99;
    11'b01000110000: data <= 32'h40e2b782;
    11'b01000110001: data <= 32'h411932d7;
    11'b01000110010: data <= 32'h3b6db315;
    11'b01000110011: data <= 32'hb55ebb70;
    11'b01000110100: data <= 32'hb6f9b6ff;
    11'b01000110101: data <= 32'hb752399c;
    11'b01000110110: data <= 32'hbc28370c;
    11'b01000110111: data <= 32'hbd2fbdf3;
    11'b01000111000: data <= 32'hb8eac173;
    11'b01000111001: data <= 32'h2ccfbdfd;
    11'b01000111010: data <= 32'hb0a73ac3;
    11'b01000111011: data <= 32'hb88a3f2f;
    11'b01000111100: data <= 32'hb0e43c67;
    11'b01000111101: data <= 32'h36cd387e;
    11'b01000111110: data <= 32'hb4453bd7;
    11'b01000111111: data <= 32'hbef73cd4;
    11'b01001000000: data <= 32'hbf0d36b0;
    11'b01001000001: data <= 32'h3606b722;
    11'b01001000010: data <= 32'h40f4b57e;
    11'b01001000011: data <= 32'h40b1318c;
    11'b01001000100: data <= 32'h3a042ff0;
    11'b01001000101: data <= 32'h2813adcc;
    11'b01001000110: data <= 32'h38fe36f0;
    11'b01001000111: data <= 32'h3aab3c2a;
    11'b01001001000: data <= 32'hb20e311e;
    11'b01001001001: data <= 32'hbc95bfd9;
    11'b01001001010: data <= 32'hba6ac1f4;
    11'b01001001011: data <= 32'h302bbe76;
    11'b01001001100: data <= 32'h35c13624;
    11'b01001001101: data <= 32'h259839e5;
    11'b01001001110: data <= 32'ha884b22b;
    11'b01001001111: data <= 32'haee6b461;
    11'b01001010000: data <= 32'hbc573ba9;
    11'b01001010001: data <= 32'hc0b33ebb;
    11'b01001010010: data <= 32'hc0293a0b;
    11'b01001010011: data <= 32'ha8d7b882;
    11'b01001010100: data <= 32'h3e7db913;
    11'b01001010101: data <= 32'h3d07341c;
    11'b01001010110: data <= 32'h2d133a8e;
    11'b01001010111: data <= 32'h330f3b48;
    11'b01001011000: data <= 32'h3dc53cde;
    11'b01001011001: data <= 32'h3e623da0;
    11'b01001011010: data <= 32'h2c083656;
    11'b01001011011: data <= 32'hbcdebddc;
    11'b01001011100: data <= 32'hb91cc085;
    11'b01001011101: data <= 32'h3abbbcdf;
    11'b01001011110: data <= 32'h3d77a6e2;
    11'b01001011111: data <= 32'h3a4db5d5;
    11'b01001100000: data <= 32'h32cbbd3b;
    11'b01001100001: data <= 32'hb107ba84;
    11'b01001100010: data <= 32'hbc123b7e;
    11'b01001100011: data <= 32'hc0263e78;
    11'b01001100100: data <= 32'hbffc32fa;
    11'b01001100101: data <= 32'hb8fabda4;
    11'b01001100110: data <= 32'h3613bcf8;
    11'b01001100111: data <= 32'ha8f7339a;
    11'b01001101000: data <= 32'hb8d83cd9;
    11'b01001101001: data <= 32'h33a23d0f;
    11'b01001101010: data <= 32'h3e8a3d58;
    11'b01001101011: data <= 32'h3da53e48;
    11'b01001101100: data <= 32'hb7c53c33;
    11'b01001101101: data <= 32'hbe6ab418;
    11'b01001101110: data <= 32'hb6c7bc01;
    11'b01001101111: data <= 32'h3e31b897;
    11'b01001110000: data <= 32'h4025b272;
    11'b01001110001: data <= 32'h3cb5bb39;
    11'b01001110010: data <= 32'h3794be4b;
    11'b01001110011: data <= 32'h3690b926;
    11'b01001110100: data <= 32'ha0573c69;
    11'b01001110101: data <= 32'hbc243d0b;
    11'b01001110110: data <= 32'hbe3ab957;
    11'b01001110111: data <= 32'hbc29c0a9;
    11'b01001111000: data <= 32'hb817bf06;
    11'b01001111001: data <= 32'hb9df2a48;
    11'b01001111010: data <= 32'hba573b3d;
    11'b01001111011: data <= 32'h33cd38cd;
    11'b01001111100: data <= 32'h3d213901;
    11'b01001111101: data <= 32'h38683da5;
    11'b01001111110: data <= 32'hbdb53eed;
    11'b01001111111: data <= 32'hc0323b6e;
    11'b01010000000: data <= 32'hb6ac1e29;
    11'b01010000001: data <= 32'h3e7fb0e5;
    11'b01010000010: data <= 32'h3f66b139;
    11'b01010000011: data <= 32'h3aa2b9a1;
    11'b01010000100: data <= 32'h387fbb85;
    11'b01010000101: data <= 32'h3d1c2fce;
    11'b01010000110: data <= 32'h3d663dd2;
    11'b01010000111: data <= 32'h2fad3c0f;
    11'b01010001000: data <= 32'hbc55bc94;
    11'b01010001001: data <= 32'hbc77c120;
    11'b01010001010: data <= 32'hb8cabef5;
    11'b01010001011: data <= 32'hb768b1a7;
    11'b01010001100: data <= 32'hb567253f;
    11'b01010001101: data <= 32'h3605ba07;
    11'b01010001110: data <= 32'h3a8fb814;
    11'b01010001111: data <= 32'hb3783c32;
    11'b01010010000: data <= 32'hc0084023;
    11'b01010010001: data <= 32'hc0a43d9a;
    11'b01010010010: data <= 32'hb92730c6;
    11'b01010010011: data <= 32'h3b5ab45b;
    11'b01010010100: data <= 32'h39a7ad74;
    11'b01010010101: data <= 32'hb02faedf;
    11'b01010010110: data <= 32'h3680a069;
    11'b01010010111: data <= 32'h3fbf3b12;
    11'b01010011000: data <= 32'h407a3f0e;
    11'b01010011001: data <= 32'h39423c75;
    11'b01010011010: data <= 32'hbb8aba2a;
    11'b01010011011: data <= 32'hbb83bf34;
    11'b01010011100: data <= 32'h9de0bc4e;
    11'b01010011101: data <= 32'h3706b402;
    11'b01010011110: data <= 32'h3659bb4d;
    11'b01010011111: data <= 32'h38cfbff7;
    11'b01010100000: data <= 32'h397ebd6d;
    11'b01010100001: data <= 32'hb42d3a36;
    11'b01010100010: data <= 32'hbed43fd9;
    11'b01010100011: data <= 32'hc0013bf1;
    11'b01010100100: data <= 32'hbb4bb876;
    11'b01010100101: data <= 32'hb0ebbaa4;
    11'b01010100110: data <= 32'hb9a9aebf;
    11'b01010100111: data <= 32'hbc8d3524;
    11'b01010101000: data <= 32'h30673699;
    11'b01010101001: data <= 32'h401f3bdb;
    11'b01010101010: data <= 32'h40613ef0;
    11'b01010101011: data <= 32'h348a3dee;
    11'b01010101100: data <= 32'hbd01345f;
    11'b01010101101: data <= 32'hb9e1b6da;
    11'b01010101110: data <= 32'h3992ae71;
    11'b01010101111: data <= 32'h3cb8af0d;
    11'b01010110000: data <= 32'h3a39bd71;
    11'b01010110001: data <= 32'h39b8c0cd;
    11'b01010110010: data <= 32'h3c08bd96;
    11'b01010110011: data <= 32'h38bd3aa5;
    11'b01010110100: data <= 32'hb8863e77;
    11'b01010110101: data <= 32'hbcee309c;
    11'b01010110110: data <= 32'hbbf7bded;
    11'b01010110111: data <= 32'hbb7cbd5e;
    11'b01010111000: data <= 32'hbe38b214;
    11'b01010111001: data <= 32'hbe4c32d2;
    11'b01010111010: data <= 32'ha03eaf19;
    11'b01010111011: data <= 32'h3ed831f2;
    11'b01010111100: data <= 32'h3d933d0b;
    11'b01010111101: data <= 32'hb90c3f4c;
    11'b01010111110: data <= 32'hbef93d56;
    11'b01010111111: data <= 32'hb94c39e7;
    11'b01011000000: data <= 32'h3b6838db;
    11'b01011000001: data <= 32'h3c542fd3;
    11'b01011000010: data <= 32'h35d0bc99;
    11'b01011000011: data <= 32'h3823bf6b;
    11'b01011000100: data <= 32'h3e2db989;
    11'b01011000101: data <= 32'h3f453cb1;
    11'b01011000110: data <= 32'h3a013d54;
    11'b01011000111: data <= 32'hb70cb71d;
    11'b01011001000: data <= 32'hbaaebf49;
    11'b01011001001: data <= 32'hbbf2bd1e;
    11'b01011001010: data <= 32'hbd94b156;
    11'b01011001011: data <= 32'hbce2b5c6;
    11'b01011001100: data <= 32'h2e26bd50;
    11'b01011001101: data <= 32'h3ceebc6d;
    11'b01011001110: data <= 32'h38483879;
    11'b01011001111: data <= 32'hbd3f3f8c;
    11'b01011010000: data <= 32'hbfc33f08;
    11'b01011010001: data <= 32'hb9743c0f;
    11'b01011010010: data <= 32'h38053916;
    11'b01011010011: data <= 32'h2cb6341e;
    11'b01011010100: data <= 32'hb9f7b866;
    11'b01011010101: data <= 32'h239ebb11;
    11'b01011010110: data <= 32'h3f9d308b;
    11'b01011010111: data <= 32'h41493de7;
    11'b01011011000: data <= 32'h3dc43d12;
    11'b01011011001: data <= 32'hae91b525;
    11'b01011011010: data <= 32'hb87dbcc5;
    11'b01011011011: data <= 32'hb666b7b2;
    11'b01011011100: data <= 32'hb7d12e79;
    11'b01011011101: data <= 32'hb708bbd8;
    11'b01011011110: data <= 32'h3545c0fb;
    11'b01011011111: data <= 32'h3bcdc040;
    11'b01011100000: data <= 32'h34a22977;
    11'b01011100001: data <= 32'hbc893e91;
    11'b01011100010: data <= 32'hbe083d61;
    11'b01011100011: data <= 32'hb8fb3564;
    11'b01011100100: data <= 32'hb40e2c30;
    11'b01011100101: data <= 32'hbd083341;
    11'b01011100110: data <= 32'hbfc0a838;
    11'b01011100111: data <= 32'hb84fb475;
    11'b01011101000: data <= 32'h3f6435f0;
    11'b01011101001: data <= 32'h41293d71;
    11'b01011101010: data <= 32'h3c853d58;
    11'b01011101011: data <= 32'hb61c3695;
    11'b01011101100: data <= 32'hb5b62ddf;
    11'b01011101101: data <= 32'h35cc3981;
    11'b01011101110: data <= 32'h366d3879;
    11'b01011101111: data <= 32'h2c66bcd9;
    11'b01011110000: data <= 32'h3637c1c2;
    11'b01011110001: data <= 32'h3c22c085;
    11'b01011110010: data <= 32'h3ac0253e;
    11'b01011110011: data <= 32'hadae3d17;
    11'b01011110100: data <= 32'hb85c3743;
    11'b01011110101: data <= 32'hb5ddb99e;
    11'b01011110110: data <= 32'hba50b882;
    11'b01011110111: data <= 32'hc0293165;
    11'b01011111000: data <= 32'hc1012d3e;
    11'b01011111001: data <= 32'hba7fb82a;
    11'b01011111010: data <= 32'h3dc7b517;
    11'b01011111011: data <= 32'h3f0339a7;
    11'b01011111100: data <= 32'h30423d4f;
    11'b01011111101: data <= 32'hbbcc3ccf;
    11'b01011111110: data <= 32'hb46f3ceb;
    11'b01011111111: data <= 32'h3a363e3c;
    11'b01100000000: data <= 32'h38823bc8;
    11'b01100000001: data <= 32'hb34cbb51;
    11'b01100000010: data <= 32'h282ec09f;
    11'b01100000011: data <= 32'h3ce6be08;
    11'b01100000100: data <= 32'h3f243701;
    11'b01100000101: data <= 32'h3cc73bf0;
    11'b01100000110: data <= 32'h3703b494;
    11'b01100000111: data <= 32'h26dcbd1e;
    11'b01100001000: data <= 32'hb9ccb907;
    11'b01100001001: data <= 32'hbf9f3523;
    11'b01100001010: data <= 32'hc049b14a;
    11'b01100001011: data <= 32'hb955bdcc;
    11'b01100001100: data <= 32'h3bc3be47;
    11'b01100001101: data <= 32'h3a2ab294;
    11'b01100001110: data <= 32'hba183c73;
    11'b01100001111: data <= 32'hbd3a3de0;
    11'b01100010000: data <= 32'hb2573dfe;
    11'b01100010001: data <= 32'h393c3e82;
    11'b01100010010: data <= 32'hb10a3c71;
    11'b01100010011: data <= 32'hbd24b4f1;
    11'b01100010100: data <= 32'hb97ebcf6;
    11'b01100010101: data <= 32'h3d19b7bb;
    11'b01100010110: data <= 32'h40d83b0c;
    11'b01100010111: data <= 32'h3f883ade;
    11'b01100011000: data <= 32'h3ae6b6fc;
    11'b01100011001: data <= 32'h35b7bb77;
    11'b01100011010: data <= 32'haed92ebd;
    11'b01100011011: data <= 32'hbb5f3a69;
    11'b01100011100: data <= 32'hbccdb750;
    11'b01100011101: data <= 32'hb4bdc0cc;
    11'b01100011110: data <= 32'h395dc12d;
    11'b01100011111: data <= 32'h347abad2;
    11'b01100100000: data <= 32'hbae83a07;
    11'b01100100001: data <= 32'hbba73c05;
    11'b01100100010: data <= 32'h2b853a1a;
    11'b01100100011: data <= 32'h33733b75;
    11'b01100100100: data <= 32'hbd093ba9;
    11'b01100100101: data <= 32'hc0f73358;
    11'b01100100110: data <= 32'hbda2b6b3;
    11'b01100100111: data <= 32'h3c342510;
    11'b01100101000: data <= 32'h408f3af3;
    11'b01100101001: data <= 32'h3e203a03;
    11'b01100101010: data <= 32'h3807a89a;
    11'b01100101011: data <= 32'h377a2ef4;
    11'b01100101100: data <= 32'h39563d1e;
    11'b01100101101: data <= 32'h310b3dd6;
    11'b01100101110: data <= 32'hb6d8b794;
    11'b01100101111: data <= 32'haf30c15c;
    11'b01100110000: data <= 32'h38aac167;
    11'b01100110001: data <= 32'h3816bac1;
    11'b01100110010: data <= 32'hac9e3708;
    11'b01100110011: data <= 32'h1d302e7c;
    11'b01100110100: data <= 32'h3848b707;
    11'b01100110101: data <= 32'haa482afb;
    11'b01100110110: data <= 32'hbfcf3a12;
    11'b01100110111: data <= 32'hc2163754;
    11'b01100111000: data <= 32'hbed0b5a5;
    11'b01100111001: data <= 32'h393fb676;
    11'b01100111010: data <= 32'h3db73367;
    11'b01100111011: data <= 32'h364f381e;
    11'b01100111100: data <= 32'hb50b378d;
    11'b01100111101: data <= 32'h36663c63;
    11'b01100111110: data <= 32'h3caa4054;
    11'b01100111111: data <= 32'h38dd3fc9;
    11'b01101000000: data <= 32'hb72fb04b;
    11'b01101000001: data <= 32'hb6d7c026;
    11'b01101000010: data <= 32'h3869bf56;
    11'b01101000011: data <= 32'h3c98b369;
    11'b01101000100: data <= 32'h3c2b34cf;
    11'b01101000101: data <= 32'h3c14b99f;
    11'b01101000110: data <= 32'h3c37bd24;
    11'b01101000111: data <= 32'h2efab4b1;
    11'b01101001000: data <= 32'hbee83abf;
    11'b01101001001: data <= 32'hc13136ab;
    11'b01101001010: data <= 32'hbd9bbbbd;
    11'b01101001011: data <= 32'h34e6bddf;
    11'b01101001100: data <= 32'h3653b9c0;
    11'b01101001101: data <= 32'hba043030;
    11'b01101001110: data <= 32'hbb7838c1;
    11'b01101001111: data <= 32'h362a3d34;
    11'b01101010000: data <= 32'h3ce8405a;
    11'b01101010001: data <= 32'h32843fe8;
    11'b01101010010: data <= 32'hbd3335f8;
    11'b01101010011: data <= 32'hbcbabbae;
    11'b01101010100: data <= 32'h366ab89c;
    11'b01101010101: data <= 32'h3e6337f3;
    11'b01101010110: data <= 32'h3e9a3487;
    11'b01101010111: data <= 32'h3daebc0c;
    11'b01101011000: data <= 32'h3d55bd04;
    11'b01101011001: data <= 32'h395132e7;
    11'b01101011010: data <= 32'hb99b3d63;
    11'b01101011011: data <= 32'hbdc53577;
    11'b01101011100: data <= 32'hba09bec6;
    11'b01101011101: data <= 32'h3076c0c8;
    11'b01101011110: data <= 32'hb36ebd7d;
    11'b01101011111: data <= 32'hbca9b390;
    11'b01101100000: data <= 32'hbaa030c1;
    11'b01101100001: data <= 32'h392a382f;
    11'b01101100010: data <= 32'h3c1b3d34;
    11'b01101100011: data <= 32'hb9323e45;
    11'b01101100100: data <= 32'hc0c53a2b;
    11'b01101100101: data <= 32'hbfbda582;
    11'b01101100110: data <= 32'h2f46338e;
    11'b01101100111: data <= 32'h3db43a03;
    11'b01101101000: data <= 32'h3d033255;
    11'b01101101001: data <= 32'h3b52baa4;
    11'b01101101010: data <= 32'h3ce3b7b1;
    11'b01101101011: data <= 32'h3d363d0e;
    11'b01101101100: data <= 32'h37a6401a;
    11'b01101101101: data <= 32'hb5df36ff;
    11'b01101101110: data <= 32'hb489bf9b;
    11'b01101101111: data <= 32'h2e9ac0e8;
    11'b01101110000: data <= 32'hb2bbbd06;
    11'b01101110001: data <= 32'hb947b5ff;
    11'b01101110010: data <= 32'ha242b919;
    11'b01101110011: data <= 32'h3cb7ba22;
    11'b01101110100: data <= 32'h3b2c3041;
    11'b01101110101: data <= 32'hbceb3c46;
    11'b01101110110: data <= 32'hc1ca3b5b;
    11'b01101110111: data <= 32'hc05233a9;
    11'b01101111000: data <= 32'hb1162f46;
    11'b01101111001: data <= 32'h39523490;
    11'b01101111010: data <= 32'h28c0adfa;
    11'b01101111011: data <= 32'hb19fb806;
    11'b01101111100: data <= 32'h3ad235c6;
    11'b01101111101: data <= 32'h3ecb4030;
    11'b01101111110: data <= 32'h3c6e4105;
    11'b01101111111: data <= 32'hacb839ad;
    11'b01110000000: data <= 32'hb659bd6a;
    11'b01110000001: data <= 32'h27e5be0d;
    11'b01110000010: data <= 32'h333fb656;
    11'b01110000011: data <= 32'h346bb327;
    11'b01110000100: data <= 32'h3b8bbd4d;
    11'b01110000101: data <= 32'h3ed4bf1b;
    11'b01110000110: data <= 32'h3c2cb84f;
    11'b01110000111: data <= 32'hbc1d3b5a;
    11'b01110001000: data <= 32'hc0c33b28;
    11'b01110001001: data <= 32'hbe93b14a;
    11'b01110001010: data <= 32'hb3b8b9ef;
    11'b01110001011: data <= 32'hb403b8c0;
    11'b01110001100: data <= 32'hbd0cb823;
    11'b01110001101: data <= 32'hbc7eb6c3;
    11'b01110001110: data <= 32'h389a3871;
    11'b01110001111: data <= 32'h3efe401a;
    11'b01110010000: data <= 32'h3b4f40bc;
    11'b01110010001: data <= 32'hb9833bde;
    11'b01110010010: data <= 32'hbc3db59c;
    11'b01110010011: data <= 32'hb1abaf32;
    11'b01110010100: data <= 32'h38b0394d;
    11'b01110010101: data <= 32'h3abb29a9;
    11'b01110010110: data <= 32'h3d34be64;
    11'b01110010111: data <= 32'h3f70bfd0;
    11'b01110011000: data <= 32'h3da3b4a9;
    11'b01110011001: data <= 32'hae863d38;
    11'b01110011010: data <= 32'hbc633b0e;
    11'b01110011011: data <= 32'hb961ba1f;
    11'b01110011100: data <= 32'haef2be5c;
    11'b01110011101: data <= 32'hba8fbcdb;
    11'b01110011110: data <= 32'hbf86ba75;
    11'b01110011111: data <= 32'hbd38b9d8;
    11'b01110100000: data <= 32'h397fb085;
    11'b01110100001: data <= 32'h3e6b3c3d;
    11'b01110100010: data <= 32'h32cf3e9a;
    11'b01110100011: data <= 32'hbead3c50;
    11'b01110100100: data <= 32'hbf22381b;
    11'b01110100101: data <= 32'hb6ea3b3d;
    11'b01110100110: data <= 32'h37fa3ceb;
    11'b01110100111: data <= 32'h3806308c;
    11'b01110101000: data <= 32'h3995bdd6;
    11'b01110101001: data <= 32'h3de2bd68;
    11'b01110101010: data <= 32'h3f0438f8;
    11'b01110101011: data <= 32'h3bf03fe8;
    11'b01110101100: data <= 32'h31cb3bdb;
    11'b01110101101: data <= 32'h304bbc06;
    11'b01110101110: data <= 32'h2cc8bec0;
    11'b01110101111: data <= 32'hba97bc14;
    11'b01110110000: data <= 32'hbe41b9ac;
    11'b01110110001: data <= 32'hb93fbcfd;
    11'b01110110010: data <= 32'h3cb4bd5f;
    11'b01110110011: data <= 32'h3e05b4db;
    11'b01110110100: data <= 32'hb5b13a66;
    11'b01110110101: data <= 32'hc0613bc9;
    11'b01110110110: data <= 32'hbfce3a3d;
    11'b01110110111: data <= 32'hb81f3be2;
    11'b01110111000: data <= 32'ha7363bbb;
    11'b01110111001: data <= 32'hb908ad71;
    11'b01110111010: data <= 32'hb89cbcb9;
    11'b01110111011: data <= 32'h39f8b87c;
    11'b01110111100: data <= 32'h3f7c3dc5;
    11'b01110111101: data <= 32'h3e6e40cb;
    11'b01110111110: data <= 32'h39853c73;
    11'b01110111111: data <= 32'h3435b936;
    11'b01111000000: data <= 32'h2e2cba94;
    11'b01111000001: data <= 32'hb716206d;
    11'b01111000010: data <= 32'hb9b4b2c5;
    11'b01111000011: data <= 32'h3445be95;
    11'b01111000100: data <= 32'h3ebbc0a5;
    11'b01111000101: data <= 32'h3e3bbccd;
    11'b01111000110: data <= 32'hb4e235eb;
    11'b01111000111: data <= 32'hbef93a89;
    11'b01111001000: data <= 32'hbd2536dc;
    11'b01111001001: data <= 32'hb45a33e3;
    11'b01111001010: data <= 32'hb93d30bc;
    11'b01111001011: data <= 32'hbf8db7f3;
    11'b01111001100: data <= 32'hbf06bc33;
    11'b01111001101: data <= 32'h30ecb41e;
    11'b01111001110: data <= 32'h3f003dd6;
    11'b01111001111: data <= 32'h3dd44043;
    11'b01111010000: data <= 32'h330a3c5e;
    11'b01111010001: data <= 32'hb4e02cba;
    11'b01111010010: data <= 32'hae3f3845;
    11'b01111010011: data <= 32'hac823d36;
    11'b01111010100: data <= 32'had21365d;
    11'b01111010101: data <= 32'h396abed8;
    11'b01111010110: data <= 32'h3efac110;
    11'b01111010111: data <= 32'h3eaebc7f;
    11'b01111011000: data <= 32'h35d038f4;
    11'b01111011001: data <= 32'hb80b3a34;
    11'b01111011010: data <= 32'had2fb10f;
    11'b01111011011: data <= 32'h3307b908;
    11'b01111011100: data <= 32'hbbebb81a;
    11'b01111011101: data <= 32'hc10fb9d1;
    11'b01111011110: data <= 32'hc044bc9b;
    11'b01111011111: data <= 32'h2d7cb9c6;
    11'b01111100000: data <= 32'h3e363825;
    11'b01111100001: data <= 32'h3a473cc4;
    11'b01111100010: data <= 32'hba013a94;
    11'b01111100011: data <= 32'hbc343979;
    11'b01111100100: data <= 32'hb51c3e44;
    11'b01111100101: data <= 32'h830d402f;
    11'b01111100110: data <= 32'hb2f539c4;
    11'b01111100111: data <= 32'h3028bdf4;
    11'b01111101000: data <= 32'h3c9ebfdd;
    11'b01111101001: data <= 32'h3ea2b416;
    11'b01111101010: data <= 32'h3cc53d2b;
    11'b01111101011: data <= 32'h3a423ade;
    11'b01111101100: data <= 32'h3bc3b818;
    11'b01111101101: data <= 32'h3962bb27;
    11'b01111101110: data <= 32'hbb03b611;
    11'b01111101111: data <= 32'hc081b758;
    11'b01111110000: data <= 32'hbe40bd55;
    11'b01111110001: data <= 32'h3860bea1;
    11'b01111110010: data <= 32'h3dc5baca;
    11'b01111110011: data <= 32'h307c2d23;
    11'b01111110100: data <= 32'hbda03681;
    11'b01111110101: data <= 32'hbd223a66;
    11'b01111110110: data <= 32'hb4433ec4;
    11'b01111110111: data <= 32'hb3363fc6;
    11'b01111111000: data <= 32'hbc5d3877;
    11'b01111111001: data <= 32'hbc8fbcc8;
    11'b01111111010: data <= 32'h3136bc83;
    11'b01111111011: data <= 32'h3dbc395e;
    11'b01111111100: data <= 32'h3e803f1d;
    11'b01111111101: data <= 32'h3d5b3b1b;
    11'b01111111110: data <= 32'h3d06b6b7;
    11'b01111111111: data <= 32'h3a70b45c;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    