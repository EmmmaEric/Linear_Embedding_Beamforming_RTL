
module memory_rom_45(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h38353df6;
    11'b00000000001: data <= 32'h35d03abc;
    11'b00000000010: data <= 32'hb46ebaec;
    11'b00000000011: data <= 32'h3313bf6f;
    11'b00000000100: data <= 32'h3e35b9fe;
    11'b00000000101: data <= 32'h40203c7b;
    11'b00000000110: data <= 32'h3d513d3b;
    11'b00000000111: data <= 32'h377db46c;
    11'b00000001000: data <= 32'h2998bd67;
    11'b00000001001: data <= 32'hb8c2b9dd;
    11'b00000001010: data <= 32'hbe202a57;
    11'b00000001011: data <= 32'hbe1eb90d;
    11'b00000001100: data <= 32'hac4fbf9d;
    11'b00000001101: data <= 32'h3ce3bf2e;
    11'b00000001110: data <= 32'h38bcb2e2;
    11'b00000001111: data <= 32'hbc903c7f;
    11'b00000010000: data <= 32'hbe9a3d5b;
    11'b00000010001: data <= 32'hb8393cc6;
    11'b00000010010: data <= 32'h328a3cd6;
    11'b00000010011: data <= 32'hb94c39e0;
    11'b00000010100: data <= 32'hbe56b6c1;
    11'b00000010101: data <= 32'hb93cbb9e;
    11'b00000010110: data <= 32'h3dca2dae;
    11'b00000010111: data <= 32'h40e43dcd;
    11'b00000011000: data <= 32'h3eb73d13;
    11'b00000011001: data <= 32'h38a9ae3c;
    11'b00000011010: data <= 32'h3278b891;
    11'b00000011011: data <= 32'ha3d435be;
    11'b00000011100: data <= 32'hb85139e7;
    11'b00000011101: data <= 32'hb8b9ba50;
    11'b00000011110: data <= 32'h358bc159;
    11'b00000011111: data <= 32'h3c83c125;
    11'b00000100000: data <= 32'h380cb945;
    11'b00000100001: data <= 32'hba063a89;
    11'b00000100010: data <= 32'hbb4e3a22;
    11'b00000100011: data <= 32'had8b347f;
    11'b00000100100: data <= 32'hb1a035b3;
    11'b00000100101: data <= 32'hbeeb36b9;
    11'b00000100110: data <= 32'hc164b090;
    11'b00000100111: data <= 32'hbd40b846;
    11'b00000101000: data <= 32'h3c9a304e;
    11'b00000101001: data <= 32'h40233c6b;
    11'b00000101010: data <= 32'h3c153c45;
    11'b00000101011: data <= 32'ha9183673;
    11'b00000101100: data <= 32'h2e9f38ec;
    11'b00000101101: data <= 32'h38303e7d;
    11'b00000101110: data <= 32'h32f03dde;
    11'b00000101111: data <= 32'hb141b91e;
    11'b00000110000: data <= 32'h3517c14d;
    11'b00000110001: data <= 32'h3c52c0a5;
    11'b00000110010: data <= 32'h3befb5bd;
    11'b00000110011: data <= 32'h35a13975;
    11'b00000110100: data <= 32'h349a8fc5;
    11'b00000110101: data <= 32'h3872b9f7;
    11'b00000110110: data <= 32'hb433b55f;
    11'b00000110111: data <= 32'hc043348a;
    11'b00000111000: data <= 32'hc1daadad;
    11'b00000111001: data <= 32'hbd77bad3;
    11'b00000111010: data <= 32'h3abcb9ca;
    11'b00000111011: data <= 32'h3cd43083;
    11'b00000111100: data <= 32'hafc33920;
    11'b00000111101: data <= 32'hbac63a18;
    11'b00000111110: data <= 32'ha8db3da0;
    11'b00000111111: data <= 32'h3a024092;
    11'b00001000000: data <= 32'h32d73f4a;
    11'b00001000001: data <= 32'hb952b42f;
    11'b00001000010: data <= 32'hb54abf85;
    11'b00001000011: data <= 32'h3b47bd1d;
    11'b00001000100: data <= 32'h3e62363b;
    11'b00001000101: data <= 32'h3db239a5;
    11'b00001000110: data <= 32'h3cf2b80d;
    11'b00001000111: data <= 32'h3c50bc9c;
    11'b00001001000: data <= 32'h2b13b3c5;
    11'b00001001001: data <= 32'hbe77390f;
    11'b00001001010: data <= 32'hc05caed7;
    11'b00001001011: data <= 32'hbabcbe61;
    11'b00001001100: data <= 32'h3963bfb3;
    11'b00001001101: data <= 32'h36b1bb40;
    11'b00001001110: data <= 32'hbb69303b;
    11'b00001001111: data <= 32'hbc8c392a;
    11'b00001010000: data <= 32'h2db13d0f;
    11'b00001010001: data <= 32'h39883fd5;
    11'b00001010010: data <= 32'hb7c33e7f;
    11'b00001010011: data <= 32'hbf482f9b;
    11'b00001010100: data <= 32'hbd3dbb1c;
    11'b00001010101: data <= 32'h388eb279;
    11'b00001010110: data <= 32'h3f2f3b97;
    11'b00001010111: data <= 32'h3ed9397e;
    11'b00001011000: data <= 32'h3d5eb884;
    11'b00001011001: data <= 32'h3ccab993;
    11'b00001011010: data <= 32'h38c53978;
    11'b00001011011: data <= 32'hb86f3db2;
    11'b00001011100: data <= 32'hbc1a944c;
    11'b00001011101: data <= 32'hb264c04a;
    11'b00001011110: data <= 32'h38fdc144;
    11'b00001011111: data <= 32'h2fc2bd82;
    11'b00001100000: data <= 32'hbaddb22e;
    11'b00001100001: data <= 32'hb8a22cea;
    11'b00001100010: data <= 32'h38ff34a5;
    11'b00001100011: data <= 32'h38b93b5b;
    11'b00001100100: data <= 32'hbd363c5f;
    11'b00001100101: data <= 32'hc1b4355c;
    11'b00001100110: data <= 32'hc00eb496;
    11'b00001100111: data <= 32'h323f310b;
    11'b00001101000: data <= 32'h3d863a6a;
    11'b00001101001: data <= 32'h3bf9368c;
    11'b00001101010: data <= 32'h388db593;
    11'b00001101011: data <= 32'h3b403302;
    11'b00001101100: data <= 32'h3c403f72;
    11'b00001101101: data <= 32'h35c7407c;
    11'b00001101110: data <= 32'hb4b2347a;
    11'b00001101111: data <= 32'ha159c016;
    11'b00001110000: data <= 32'h3832c0a8;
    11'b00001110001: data <= 32'h353fbbb9;
    11'b00001110010: data <= 32'ha916b18a;
    11'b00001110011: data <= 32'h3835b8fb;
    11'b00001110100: data <= 32'h3d84bafe;
    11'b00001110101: data <= 32'h3975ac2b;
    11'b00001110110: data <= 32'hbe5a39c7;
    11'b00001110111: data <= 32'hc20f368c;
    11'b00001111000: data <= 32'hc006b56d;
    11'b00001111001: data <= 32'h9cb6b666;
    11'b00001111010: data <= 32'h3892aa88;
    11'b00001111011: data <= 32'hb447b08a;
    11'b00001111100: data <= 32'hb81ab2a5;
    11'b00001111101: data <= 32'h382e3ae1;
    11'b00001111110: data <= 32'h3d2040f5;
    11'b00001111111: data <= 32'h38d94126;
    11'b00010000000: data <= 32'hb7bb38d0;
    11'b00010000001: data <= 32'hb834bd33;
    11'b00010000010: data <= 32'h336dbcb2;
    11'b00010000011: data <= 32'h397a2889;
    11'b00010000100: data <= 32'h3ad02dd4;
    11'b00010000101: data <= 32'h3dbbbc65;
    11'b00010000110: data <= 32'h3fb2be0a;
    11'b00010000111: data <= 32'h3c00b4a6;
    11'b00010001000: data <= 32'hbc4d3b4a;
    11'b00010001001: data <= 32'hc06037fe;
    11'b00010001010: data <= 32'hbd0fba89;
    11'b00010001011: data <= 32'h2b09bd93;
    11'b00010001100: data <= 32'hb199bc39;
    11'b00010001101: data <= 32'hbd23b9b9;
    11'b00010001110: data <= 32'hbc82b61a;
    11'b00010001111: data <= 32'h37683987;
    11'b00010010000: data <= 32'h3d3c4024;
    11'b00010010001: data <= 32'h31a74061;
    11'b00010010010: data <= 32'hbda03a39;
    11'b00010010011: data <= 32'hbdd2b5af;
    11'b00010010100: data <= 32'hb29a2e6c;
    11'b00010010101: data <= 32'h3a313b5d;
    11'b00010010110: data <= 32'h3c543485;
    11'b00010010111: data <= 32'h3de8bce0;
    11'b00010011000: data <= 32'h3f9fbd4a;
    11'b00010011001: data <= 32'h3d7e361f;
    11'b00010011010: data <= 32'hab533e8f;
    11'b00010011011: data <= 32'hbacf39c9;
    11'b00010011100: data <= 32'hb4cabcd8;
    11'b00010011101: data <= 32'h3391c007;
    11'b00010011110: data <= 32'hb813bdee;
    11'b00010011111: data <= 32'hbdedbba6;
    11'b00010100000: data <= 32'hbabebaa1;
    11'b00010100001: data <= 32'h3b54b3f9;
    11'b00010100010: data <= 32'h3d553af0;
    11'b00010100011: data <= 32'hb73b3d64;
    11'b00010100100: data <= 32'hc0a63a01;
    11'b00010100101: data <= 32'hc04a3433;
    11'b00010100110: data <= 32'hb86339c8;
    11'b00010100111: data <= 32'h36d63c48;
    11'b00010101000: data <= 32'h362a2f4f;
    11'b00010101001: data <= 32'h387bbc80;
    11'b00010101010: data <= 32'h3d4fb8f8;
    11'b00010101011: data <= 32'h3e623db0;
    11'b00010101100: data <= 32'h3ad940e0;
    11'b00010101101: data <= 32'h30693c14;
    11'b00010101110: data <= 32'h32b0bc7f;
    11'b00010101111: data <= 32'h3472bed5;
    11'b00010110000: data <= 32'hb6aabb9b;
    11'b00010110001: data <= 32'hbb2fb97c;
    11'b00010110010: data <= 32'h2e64bd31;
    11'b00010110011: data <= 32'h3e9dbd9a;
    11'b00010110100: data <= 32'h3dedb5de;
    11'b00010110101: data <= 32'hb99f391f;
    11'b00010110110: data <= 32'hc0f73934;
    11'b00010110111: data <= 32'hc01134eb;
    11'b00010111000: data <= 32'hb85736a6;
    11'b00010111001: data <= 32'hb1c13687;
    11'b00010111010: data <= 32'hbae7b6a8;
    11'b00010111011: data <= 32'hba14bc4b;
    11'b00010111100: data <= 32'h38c7ab62;
    11'b00010111101: data <= 32'h3e724001;
    11'b00010111110: data <= 32'h3cb64167;
    11'b00010111111: data <= 32'h32c43cbf;
    11'b00011000000: data <= 32'had4eb862;
    11'b00011000001: data <= 32'h2597b889;
    11'b00011000010: data <= 32'hb1693461;
    11'b00011000011: data <= 32'hafddacf1;
    11'b00011000100: data <= 32'h3ba4be35;
    11'b00011000101: data <= 32'h4051c030;
    11'b00011000110: data <= 32'h3ecabaea;
    11'b00011000111: data <= 32'hb5113893;
    11'b00011001000: data <= 32'hbe99396c;
    11'b00011001001: data <= 32'hbc52aa9b;
    11'b00011001010: data <= 32'hb0e1b6d5;
    11'b00011001011: data <= 32'hb991b835;
    11'b00011001100: data <= 32'hbfb2bbc9;
    11'b00011001101: data <= 32'hbe9cbccb;
    11'b00011001110: data <= 32'h33ecb08e;
    11'b00011001111: data <= 32'h3e2b3e67;
    11'b00011010000: data <= 32'h3aef4047;
    11'b00011010001: data <= 32'hb83f3c39;
    11'b00011010010: data <= 32'hbb56316a;
    11'b00011010011: data <= 32'hb6a139f1;
    11'b00011010100: data <= 32'had1f3dc5;
    11'b00011010101: data <= 32'h30c236ee;
    11'b00011010110: data <= 32'h3c01be2c;
    11'b00011010111: data <= 32'h3ffcc009;
    11'b00011011000: data <= 32'h3f33b65c;
    11'b00011011001: data <= 32'h37ca3cb2;
    11'b00011011010: data <= 32'hb4853b36;
    11'b00011011011: data <= 32'h316db680;
    11'b00011011100: data <= 32'h35edbc2f;
    11'b00011011101: data <= 32'hbafcbb9b;
    11'b00011011110: data <= 32'hc073bc6e;
    11'b00011011111: data <= 32'hbe65bdb1;
    11'b00011100000: data <= 32'h3851bb1d;
    11'b00011100001: data <= 32'h3e3b35fa;
    11'b00011100010: data <= 32'h34e23c13;
    11'b00011100011: data <= 32'hbda33964;
    11'b00011100100: data <= 32'hbe6238d8;
    11'b00011100101: data <= 32'hb97f3dd8;
    11'b00011100110: data <= 32'hb41c3f64;
    11'b00011100111: data <= 32'hb621376b;
    11'b00011101000: data <= 32'h2c57bdb1;
    11'b00011101001: data <= 32'h3ca1bd9c;
    11'b00011101010: data <= 32'h3eab388c;
    11'b00011101011: data <= 32'h3cce3fcd;
    11'b00011101100: data <= 32'h3a613ca3;
    11'b00011101101: data <= 32'h3baab6ff;
    11'b00011101110: data <= 32'h3937bafb;
    11'b00011101111: data <= 32'hb9d3b68a;
    11'b00011110000: data <= 32'hbef4b8d5;
    11'b00011110001: data <= 32'hba1bbe34;
    11'b00011110010: data <= 32'h3cf5bf56;
    11'b00011110011: data <= 32'h3ec2bb8e;
    11'b00011110100: data <= 32'ha4332185;
    11'b00011110101: data <= 32'hbeab34ae;
    11'b00011110110: data <= 32'hbded388f;
    11'b00011110111: data <= 32'hb7bb3d0c;
    11'b00011111000: data <= 32'hb8693d4f;
    11'b00011111001: data <= 32'hbdb69d4d;
    11'b00011111010: data <= 32'hbd51bd78;
    11'b00011111011: data <= 32'h2f55ba77;
    11'b00011111100: data <= 32'h3d773cdf;
    11'b00011111101: data <= 32'h3da74070;
    11'b00011111110: data <= 32'h3bdf3caa;
    11'b00011111111: data <= 32'h3ac5b057;
    11'b00100000000: data <= 32'h37db2cdf;
    11'b00100000001: data <= 32'hb7b53b14;
    11'b00100000010: data <= 32'hbbbe3515;
    11'b00100000011: data <= 32'h3034bddb;
    11'b00100000100: data <= 32'h3f06c0c8;
    11'b00100000101: data <= 32'h3f24be3c;
    11'b00100000110: data <= 32'h3062b46f;
    11'b00100000111: data <= 32'hbc0b31d5;
    11'b00100001000: data <= 32'hb7813286;
    11'b00100001001: data <= 32'h32c53740;
    11'b00100001010: data <= 32'hb9bd362d;
    11'b00100001011: data <= 32'hc0abb89b;
    11'b00100001100: data <= 32'hc0aebda6;
    11'b00100001101: data <= 32'hb7dbb9a1;
    11'b00100001110: data <= 32'h3c743bcf;
    11'b00100001111: data <= 32'h3c4f3e71;
    11'b00100010000: data <= 32'h34ce3a02;
    11'b00100010001: data <= 32'h295f337d;
    11'b00100010010: data <= 32'h2a3a3ce3;
    11'b00100010011: data <= 32'hb585405a;
    11'b00100010100: data <= 32'hb8683c76;
    11'b00100010101: data <= 32'h3524bce8;
    11'b00100010110: data <= 32'h3e43c089;
    11'b00100010111: data <= 32'h3e88bcae;
    11'b00100011000: data <= 32'h38d93414;
    11'b00100011001: data <= 32'h32073649;
    11'b00100011010: data <= 32'h3b3eb19c;
    11'b00100011011: data <= 32'h3c30b452;
    11'b00100011100: data <= 32'hb902b13a;
    11'b00100011101: data <= 32'hc122b9a1;
    11'b00100011110: data <= 32'hc0c4bdad;
    11'b00100011111: data <= 32'hb4fdbc8e;
    11'b00100100000: data <= 32'h3c57ad3b;
    11'b00100100001: data <= 32'h380335e7;
    11'b00100100010: data <= 32'hb92a2907;
    11'b00100100011: data <= 32'hb9ea35ed;
    11'b00100100100: data <= 32'hb38b3f6a;
    11'b00100100101: data <= 32'hb5924164;
    11'b00100100110: data <= 32'hba6a3d38;
    11'b00100100111: data <= 32'hb718bc1b;
    11'b00100101000: data <= 32'h38f1be8e;
    11'b00100101001: data <= 32'h3cabb16b;
    11'b00100101010: data <= 32'h3bfc3c6e;
    11'b00100101011: data <= 32'h3caa3962;
    11'b00100101100: data <= 32'h3f4eb56c;
    11'b00100101101: data <= 32'h3e24b576;
    11'b00100101110: data <= 32'hb5c232cd;
    11'b00100101111: data <= 32'hc01faf1a;
    11'b00100110000: data <= 32'hbe2bbce7;
    11'b00100110001: data <= 32'h36f1bf00;
    11'b00100110010: data <= 32'h3cf7bd25;
    11'b00100110011: data <= 32'h2d3eba4e;
    11'b00100110100: data <= 32'hbc73b8c2;
    11'b00100110101: data <= 32'hba493166;
    11'b00100110110: data <= 32'h28323e82;
    11'b00100110111: data <= 32'hb5864066;
    11'b00100111000: data <= 32'hbe0e3a9d;
    11'b00100111001: data <= 32'hbeddbbe6;
    11'b00100111010: data <= 32'hb8a9bbc9;
    11'b00100111011: data <= 32'h38963943;
    11'b00100111100: data <= 32'h3c003e1f;
    11'b00100111101: data <= 32'h3d443920;
    11'b00100111110: data <= 32'h3f17b4d7;
    11'b00100111111: data <= 32'h3da43498;
    11'b00101000000: data <= 32'haf223d80;
    11'b00101000001: data <= 32'hbcf43bc1;
    11'b00101000010: data <= 32'hb802ba8d;
    11'b00101000011: data <= 32'h3c63c01e;
    11'b00101000100: data <= 32'h3d4bbf69;
    11'b00101000101: data <= 32'h1dcabcab;
    11'b00101000110: data <= 32'hba11ba5a;
    11'b00101000111: data <= 32'h2db3b34d;
    11'b00101001000: data <= 32'h3b073a3d;
    11'b00101001001: data <= 32'hb1b33c93;
    11'b00101001010: data <= 32'hc04a2fd3;
    11'b00101001011: data <= 32'hc157bc28;
    11'b00101001100: data <= 32'hbd3db965;
    11'b00101001101: data <= 32'h31a03997;
    11'b00101001110: data <= 32'h38c33c44;
    11'b00101001111: data <= 32'h38cf2dc9;
    11'b00101010000: data <= 32'h3b1eb441;
    11'b00101010001: data <= 32'h3ad83c90;
    11'b00101010010: data <= 32'h1a484133;
    11'b00101010011: data <= 32'hb94c3fa9;
    11'b00101010100: data <= 32'haa1cb624;
    11'b00101010101: data <= 32'h3c3ebf4d;
    11'b00101010110: data <= 32'h3c3cbdbc;
    11'b00101010111: data <= 32'h30dcb8c3;
    11'b00101011000: data <= 32'h3076b80b;
    11'b00101011001: data <= 32'h3d91b8a8;
    11'b00101011010: data <= 32'h3f88ac9c;
    11'b00101011011: data <= 32'h310835a8;
    11'b00101011100: data <= 32'hc074b175;
    11'b00101011101: data <= 32'hc15dbbb7;
    11'b00101011110: data <= 32'hbc86ba72;
    11'b00101011111: data <= 32'h31d2aaff;
    11'b00101100000: data <= 32'h286aae14;
    11'b00101100001: data <= 32'hb72cba6e;
    11'b00101100010: data <= 32'haee1b695;
    11'b00101100011: data <= 32'h366a3e5a;
    11'b00101100100: data <= 32'h2a6b422f;
    11'b00101100101: data <= 32'hb917404b;
    11'b00101100110: data <= 32'hb811b156;
    11'b00101100111: data <= 32'h3297bcc2;
    11'b00101101000: data <= 32'h3685b590;
    11'b00101101001: data <= 32'h3386371e;
    11'b00101101010: data <= 32'h3b3dab70;
    11'b00101101011: data <= 32'h4093ba25;
    11'b00101101100: data <= 32'h40e9b63b;
    11'b00101101101: data <= 32'h37eb36e0;
    11'b00101101110: data <= 32'hbec134fb;
    11'b00101101111: data <= 32'hbf14b8c6;
    11'b00101110000: data <= 32'hb360bc5f;
    11'b00101110001: data <= 32'h37debc17;
    11'b00101110010: data <= 32'hb636bceb;
    11'b00101110011: data <= 32'hbc87be42;
    11'b00101110100: data <= 32'hb721b9eb;
    11'b00101110101: data <= 32'h384f3d31;
    11'b00101110110: data <= 32'h32944113;
    11'b00101110111: data <= 32'hbc173e34;
    11'b00101111000: data <= 32'hbe1bb421;
    11'b00101111001: data <= 32'hbbc3b83e;
    11'b00101111010: data <= 32'hb58f395d;
    11'b00101111011: data <= 32'h2b333c99;
    11'b00101111100: data <= 32'h3bb02b9d;
    11'b00101111101: data <= 32'h4062bad9;
    11'b00101111110: data <= 32'h4084acf6;
    11'b00101111111: data <= 32'h392c3d4b;
    11'b00110000000: data <= 32'hbaf93d70;
    11'b00110000001: data <= 32'hb87a9cb4;
    11'b00110000010: data <= 32'h399fbcb3;
    11'b00110000011: data <= 32'h39e9bddc;
    11'b00110000100: data <= 32'hb87abe56;
    11'b00110000101: data <= 32'hbc51bef7;
    11'b00110000110: data <= 32'h30d4bc56;
    11'b00110000111: data <= 32'h3d5a3731;
    11'b00110001000: data <= 32'h388b3d56;
    11'b00110001001: data <= 32'hbd9038bd;
    11'b00110001010: data <= 32'hc0a8b7c2;
    11'b00110001011: data <= 32'hbebfb13a;
    11'b00110001100: data <= 32'hba383bfa;
    11'b00110001101: data <= 32'hb5973bc7;
    11'b00110001110: data <= 32'h335eb6d0;
    11'b00110001111: data <= 32'h3cbdbc0d;
    11'b00110010000: data <= 32'h3de637d6;
    11'b00110010001: data <= 32'h38ae40bf;
    11'b00110010010: data <= 32'hb3ff409c;
    11'b00110010011: data <= 32'h3136381b;
    11'b00110010100: data <= 32'h3bb2bb13;
    11'b00110010101: data <= 32'h387fbc0b;
    11'b00110010110: data <= 32'hb8c4bb4a;
    11'b00110010111: data <= 32'hb7b0bd0c;
    11'b00110011000: data <= 32'h3d0abd19;
    11'b00110011001: data <= 32'h40b3b6e2;
    11'b00110011010: data <= 32'h3c1d34ad;
    11'b00110011011: data <= 32'hbd729bfa;
    11'b00110011100: data <= 32'hc091b835;
    11'b00110011101: data <= 32'hbdbbb031;
    11'b00110011110: data <= 32'hb9013864;
    11'b00110011111: data <= 32'hba2c25b6;
    11'b00110100000: data <= 32'hbab4bd4f;
    11'b00110100001: data <= 32'ha9c0bd45;
    11'b00110100010: data <= 32'h39b73a40;
    11'b00110100011: data <= 32'h37d44193;
    11'b00110100100: data <= 32'had6b40f9;
    11'b00110100101: data <= 32'h21463919;
    11'b00110100110: data <= 32'h356fb598;
    11'b00110100111: data <= 32'hadaf2e05;
    11'b00110101000: data <= 32'hb9903571;
    11'b00110101001: data <= 32'h2dc4b81f;
    11'b00110101010: data <= 32'h4020bd2f;
    11'b00110101011: data <= 32'h41ccbae4;
    11'b00110101100: data <= 32'h3d502bf1;
    11'b00110101101: data <= 32'hbb0c331f;
    11'b00110101110: data <= 32'hbd62b1a6;
    11'b00110101111: data <= 32'hb57eb327;
    11'b00110110000: data <= 32'ha870b220;
    11'b00110110001: data <= 32'hbc16bc02;
    11'b00110110010: data <= 32'hbe74c02e;
    11'b00110110011: data <= 32'hb979bea7;
    11'b00110110100: data <= 32'h38973804;
    11'b00110110101: data <= 32'h38cb4067;
    11'b00110110110: data <= 32'hb46d3eea;
    11'b00110110111: data <= 32'hba0934ad;
    11'b00110111000: data <= 32'hb9a8307e;
    11'b00110111001: data <= 32'hbaee3cbf;
    11'b00110111010: data <= 32'hbb8d3d5b;
    11'b00110111011: data <= 32'h2f14ae67;
    11'b00110111100: data <= 32'h3fb6bd3b;
    11'b00110111101: data <= 32'h4124b9dd;
    11'b00110111110: data <= 32'h3d0e3977;
    11'b00110111111: data <= 32'hb30a3c79;
    11'b00111000000: data <= 32'hac843729;
    11'b00111000001: data <= 32'h3b01b216;
    11'b00111000010: data <= 32'h3831b86d;
    11'b00111000011: data <= 32'hbc5abd3f;
    11'b00111000100: data <= 32'hbeeac05a;
    11'b00111000101: data <= 32'hb5fbbf5c;
    11'b00111000110: data <= 32'h3cc7b2d8;
    11'b00111000111: data <= 32'h3bec3b86;
    11'b00111001000: data <= 32'hb7f137f0;
    11'b00111001001: data <= 32'hbdbdb40e;
    11'b00111001010: data <= 32'hbd7d360f;
    11'b00111001011: data <= 32'hbcf83eaa;
    11'b00111001100: data <= 32'hbcf43dd6;
    11'b00111001101: data <= 32'hb826b612;
    11'b00111001110: data <= 32'h3af1bdec;
    11'b00111001111: data <= 32'h3e21b558;
    11'b00111010000: data <= 32'h3b163e4e;
    11'b00111010001: data <= 32'h34194001;
    11'b00111010010: data <= 32'h3a553b95;
    11'b00111010011: data <= 32'h3dc72a1c;
    11'b00111010100: data <= 32'h38abb139;
    11'b00111010101: data <= 32'hbc7ab8bd;
    11'b00111010110: data <= 32'hbd3bbde0;
    11'b00111010111: data <= 32'h3863beea;
    11'b00111011000: data <= 32'h4043bb84;
    11'b00111011001: data <= 32'h3dd9b359;
    11'b00111011010: data <= 32'hb773b6b9;
    11'b00111011011: data <= 32'hbda8b87f;
    11'b00111011100: data <= 32'hbc4e3617;
    11'b00111011101: data <= 32'hbb373d9a;
    11'b00111011110: data <= 32'hbd8f39c9;
    11'b00111011111: data <= 32'hbdbdbcc2;
    11'b00111100000: data <= 32'hb7a6bf42;
    11'b00111100001: data <= 32'h3726adde;
    11'b00111100010: data <= 32'h37e53fe8;
    11'b00111100011: data <= 32'h35ce404b;
    11'b00111100100: data <= 32'h3a923b65;
    11'b00111100101: data <= 32'h3c4035ae;
    11'b00111100110: data <= 32'h2a253a6c;
    11'b00111100111: data <= 32'hbd083a1d;
    11'b00111101000: data <= 32'hba99b66c;
    11'b00111101001: data <= 32'h3d37bdbc;
    11'b00111101010: data <= 32'h414bbd23;
    11'b00111101011: data <= 32'h3ea1b91d;
    11'b00111101100: data <= 32'hb133b768;
    11'b00111101101: data <= 32'hb8c0b5c2;
    11'b00111101110: data <= 32'h2eec3535;
    11'b00111101111: data <= 32'h9abd3a3b;
    11'b00111110000: data <= 32'hbd42b325;
    11'b00111110001: data <= 32'hc034bfb1;
    11'b00111110010: data <= 32'hbd2bc032;
    11'b00111110011: data <= 32'h20fab3d1;
    11'b00111110100: data <= 32'h36b23df0;
    11'b00111110101: data <= 32'h32403d37;
    11'b00111110110: data <= 32'h326234b6;
    11'b00111110111: data <= 32'h300a3836;
    11'b00111111000: data <= 32'hb9973f1a;
    11'b00111111001: data <= 32'hbdef3fba;
    11'b00111111010: data <= 32'hb9d33554;
    11'b00111111011: data <= 32'h3cf4bce2;
    11'b00111111100: data <= 32'h4080bca3;
    11'b00111111101: data <= 32'h3d5cb1b1;
    11'b00111111110: data <= 32'h3258349b;
    11'b00111111111: data <= 32'h38773321;
    11'b01000000000: data <= 32'h3df735e1;
    11'b01000000001: data <= 32'h3b22363d;
    11'b01000000010: data <= 32'hbc7cb8a0;
    11'b01000000011: data <= 32'hc064bfd4;
    11'b01000000100: data <= 32'hbc9cc020;
    11'b01000000101: data <= 32'h3733b982;
    11'b01000000110: data <= 32'h39f8357b;
    11'b01000000111: data <= 32'h1adead98;
    11'b01000001000: data <= 32'hb76bb8c7;
    11'b01000001001: data <= 32'hb87837a1;
    11'b01000001010: data <= 32'hbc2c406d;
    11'b01000001011: data <= 32'hbe734077;
    11'b01000001100: data <= 32'hbc7e3456;
    11'b01000001101: data <= 32'h34a9bd32;
    11'b01000001110: data <= 32'h3c40ba5a;
    11'b01000001111: data <= 32'h38ec394b;
    11'b01000010000: data <= 32'h35e33ca8;
    11'b01000010001: data <= 32'h3d7239a5;
    11'b01000010010: data <= 32'h408037d3;
    11'b01000010011: data <= 32'h3cd338b6;
    11'b01000010100: data <= 32'hbc1728be;
    11'b01000010101: data <= 32'hbf39bc79;
    11'b01000010110: data <= 32'hb504be79;
    11'b01000010111: data <= 32'h3d65bc66;
    11'b01000011000: data <= 32'h3cd3ba0b;
    11'b01000011001: data <= 32'ha8d8bcd0;
    11'b01000011010: data <= 32'hb8b4bcca;
    11'b01000011011: data <= 32'hb5ae34f7;
    11'b01000011100: data <= 32'hb8c03fdf;
    11'b01000011101: data <= 32'hbdd43e6c;
    11'b01000011110: data <= 32'hbeebb781;
    11'b01000011111: data <= 32'hbbc9be7a;
    11'b01000100000: data <= 32'hb352b81e;
    11'b01000100001: data <= 32'hae8e3ca7;
    11'b01000100010: data <= 32'h34453d8c;
    11'b01000100011: data <= 32'h3d9a38cc;
    11'b01000100100: data <= 32'h40023838;
    11'b01000100101: data <= 32'h3a373d0c;
    11'b01000100110: data <= 32'hbc8b3d3a;
    11'b01000100111: data <= 32'hbd3f30f2;
    11'b01000101000: data <= 32'h3809bbc9;
    11'b01000101001: data <= 32'h3fb9bccd;
    11'b01000101010: data <= 32'h3d61bca6;
    11'b01000101011: data <= 32'h2924bda1;
    11'b01000101100: data <= 32'ha852bc94;
    11'b01000101101: data <= 32'h39ed32ad;
    11'b01000101110: data <= 32'h38023d69;
    11'b01000101111: data <= 32'hbc16390e;
    11'b01000110000: data <= 32'hc040bd03;
    11'b01000110001: data <= 32'hbf15bf7c;
    11'b01000110010: data <= 32'hbad1b7cb;
    11'b01000110011: data <= 32'hb6043b3f;
    11'b01000110100: data <= 32'h25903910;
    11'b01000110101: data <= 32'h3a5db2be;
    11'b01000110110: data <= 32'h3c4d3577;
    11'b01000110111: data <= 32'h90833fcb;
    11'b01000111000: data <= 32'hbd6440e5;
    11'b01000111001: data <= 32'hbc503c63;
    11'b01000111010: data <= 32'h3923b81a;
    11'b01000111011: data <= 32'h3e7cbbae;
    11'b01000111100: data <= 32'h3af5b9c4;
    11'b01000111101: data <= 32'h2ba8b99b;
    11'b01000111110: data <= 32'h3aa0b87b;
    11'b01000111111: data <= 32'h402e33e8;
    11'b01001000000: data <= 32'h3e7b3aed;
    11'b01001000001: data <= 32'hb84e2ec1;
    11'b01001000010: data <= 32'hc021bd83;
    11'b01001000011: data <= 32'hbe9abed2;
    11'b01001000100: data <= 32'hb7e3b8ed;
    11'b01001000101: data <= 32'had5d2a33;
    11'b01001000110: data <= 32'hb19eb9c3;
    11'b01001000111: data <= 32'h2c5cbd58;
    11'b01001001000: data <= 32'h3405a7f4;
    11'b01001001001: data <= 32'hb7044064;
    11'b01001001010: data <= 32'hbd854187;
    11'b01001001011: data <= 32'hbcc43c9b;
    11'b01001001100: data <= 32'ha7dab814;
    11'b01001001101: data <= 32'h37a9b898;
    11'b01001001110: data <= 32'hadd9310a;
    11'b01001001111: data <= 32'haf7a347c;
    11'b01001010000: data <= 32'h3da72299;
    11'b01001010001: data <= 32'h41ba34e4;
    11'b01001010010: data <= 32'h402d3a95;
    11'b01001010011: data <= 32'hb4ef375f;
    11'b01001010100: data <= 32'hbe84b8c1;
    11'b01001010101: data <= 32'hba51bc21;
    11'b01001010110: data <= 32'h379cb95a;
    11'b01001010111: data <= 32'h3746ba7f;
    11'b01001011000: data <= 32'hb40bbf68;
    11'b01001011001: data <= 32'hb41bc040;
    11'b01001011010: data <= 32'h32d2b614;
    11'b01001011011: data <= 32'hab693f82;
    11'b01001011100: data <= 32'hbc134041;
    11'b01001011101: data <= 32'hbdc33611;
    11'b01001011110: data <= 32'hbc2dbb19;
    11'b01001011111: data <= 32'hba9fb46a;
    11'b01001100000: data <= 32'hbc1f3a92;
    11'b01001100001: data <= 32'hb73339ca;
    11'b01001100010: data <= 32'h3d65a147;
    11'b01001100011: data <= 32'h413e315e;
    11'b01001100100: data <= 32'h3eaa3c9e;
    11'b01001100101: data <= 32'hb72b3de3;
    11'b01001100110: data <= 32'hbc7c3983;
    11'b01001100111: data <= 32'h3118b088;
    11'b01001101000: data <= 32'h3d06b7e3;
    11'b01001101001: data <= 32'h3980bc57;
    11'b01001101010: data <= 32'hb511c025;
    11'b01001101011: data <= 32'ha4eac040;
    11'b01001101100: data <= 32'h3c32b7e9;
    11'b01001101101: data <= 32'h3c273cfa;
    11'b01001101110: data <= 32'hb5363c33;
    11'b01001101111: data <= 32'hbe19b8a3;
    11'b01001110000: data <= 32'hbeb9bcf5;
    11'b01001110001: data <= 32'hbdecb074;
    11'b01001110010: data <= 32'hbda03ad0;
    11'b01001110011: data <= 32'hba0c3342;
    11'b01001110100: data <= 32'h39bbba77;
    11'b01001110101: data <= 32'h3e73b45e;
    11'b01001110110: data <= 32'h39ec3e07;
    11'b01001110111: data <= 32'hba1b40db;
    11'b01001111000: data <= 32'hba763eaf;
    11'b01001111001: data <= 32'h38713784;
    11'b01001111010: data <= 32'h3ccbb068;
    11'b01001111011: data <= 32'h33bdb8ca;
    11'b01001111100: data <= 32'hb84fbd3e;
    11'b01001111101: data <= 32'h3802bdb6;
    11'b01001111110: data <= 32'h4066b5c5;
    11'b01001111111: data <= 32'h4068399e;
    11'b01010000000: data <= 32'h35a134b4;
    11'b01010000001: data <= 32'hbd2ebba0;
    11'b01010000010: data <= 32'hbdf8bc80;
    11'b01010000011: data <= 32'hbc5eaa32;
    11'b01010000100: data <= 32'hbc2e3558;
    11'b01010000101: data <= 32'hbb08bb52;
    11'b01010000110: data <= 32'haa6ebfee;
    11'b01010000111: data <= 32'h38b1bafd;
    11'b01010001000: data <= 32'h2ba43e26;
    11'b01010001001: data <= 32'hbaf5414f;
    11'b01010001010: data <= 32'hb9d63ee2;
    11'b01010001011: data <= 32'h32d73745;
    11'b01010001100: data <= 32'h346f32a3;
    11'b01010001101: data <= 32'hba1f34ff;
    11'b01010001110: data <= 32'hbbbab0fe;
    11'b01010001111: data <= 32'h3aa8b8fe;
    11'b01010010000: data <= 32'h41b9b2a3;
    11'b01010010001: data <= 32'h416037fe;
    11'b01010010010: data <= 32'h38f0354a;
    11'b01010010011: data <= 32'hbadab66c;
    11'b01010010100: data <= 32'hb8c6b6ac;
    11'b01010010101: data <= 32'h25b4312a;
    11'b01010010110: data <= 32'hb4bdb3c8;
    11'b01010010111: data <= 32'hbacabfaf;
    11'b01010011000: data <= 32'hb806c1a0;
    11'b01010011001: data <= 32'h33e5bd3f;
    11'b01010011010: data <= 32'h324b3cad;
    11'b01010011011: data <= 32'hb7e33fe7;
    11'b01010011100: data <= 32'hb9bc3aa4;
    11'b01010011101: data <= 32'hb7ecaea0;
    11'b01010011110: data <= 32'hbb1f3660;
    11'b01010011111: data <= 32'hbf113c50;
    11'b01010100000: data <= 32'hbdc3388e;
    11'b01010100001: data <= 32'h395bb64b;
    11'b01010100010: data <= 32'h4121b553;
    11'b01010100011: data <= 32'h405c38a8;
    11'b01010100100: data <= 32'h355d3c19;
    11'b01010100101: data <= 32'hb71b39d1;
    11'b01010100110: data <= 32'h36fb3866;
    11'b01010100111: data <= 32'h3c423834;
    11'b01010101000: data <= 32'h3247b5f6;
    11'b01010101001: data <= 32'hbaf9c029;
    11'b01010101010: data <= 32'hb7e3c186;
    11'b01010101011: data <= 32'h3a15bd52;
    11'b01010101100: data <= 32'h3c7b38df;
    11'b01010101101: data <= 32'h347a3a97;
    11'b01010101110: data <= 32'hb89bb5ed;
    11'b01010101111: data <= 32'hbb92b9ba;
    11'b01010110000: data <= 32'hbde63781;
    11'b01010110001: data <= 32'hc0423d3e;
    11'b01010110010: data <= 32'hbed2364d;
    11'b01010110011: data <= 32'h2d0ebbff;
    11'b01010110100: data <= 32'h3df7bac2;
    11'b01010110101: data <= 32'h3c243980;
    11'b01010110110: data <= 32'hb3723f0b;
    11'b01010110111: data <= 32'hb2e33e87;
    11'b01010111000: data <= 32'h3c0b3cbd;
    11'b01010111001: data <= 32'h3d4e3b32;
    11'b01010111010: data <= 32'ha8ec2eff;
    11'b01010111011: data <= 32'hbc96bd09;
    11'b01010111100: data <= 32'hb34bbf7e;
    11'b01010111101: data <= 32'h3ea5bbb0;
    11'b01010111110: data <= 32'h4065312c;
    11'b01010111111: data <= 32'h3c0cadcf;
    11'b01011000000: data <= 32'hb44fbc3c;
    11'b01011000001: data <= 32'hb9c3baa9;
    11'b01011000010: data <= 32'hbc1e38b9;
    11'b01011000011: data <= 32'hbe753c2f;
    11'b01011000100: data <= 32'hbe7db7ae;
    11'b01011000101: data <= 32'hb8bcc026;
    11'b01011000110: data <= 32'h3532be17;
    11'b01011000111: data <= 32'h29a638b6;
    11'b01011001000: data <= 32'hb8b93fa0;
    11'b01011001001: data <= 32'hb0433e83;
    11'b01011001010: data <= 32'h3b533c3d;
    11'b01011001011: data <= 32'h39823c53;
    11'b01011001100: data <= 32'hbb713b7b;
    11'b01011001101: data <= 32'hbea92522;
    11'b01011001110: data <= 32'hac56ba26;
    11'b01011001111: data <= 32'h406ab851;
    11'b01011010000: data <= 32'h4143a439;
    11'b01011010001: data <= 32'h3cdab4a0;
    11'b01011010010: data <= 32'h2b80ba75;
    11'b01011010011: data <= 32'h2f1ab42c;
    11'b01011010100: data <= 32'h323a3b27;
    11'b01011010101: data <= 32'hb8aa395e;
    11'b01011010110: data <= 32'hbd46bd59;
    11'b01011010111: data <= 32'hbbf6c1b6;
    11'b01011011000: data <= 32'hb390bfc4;
    11'b01011011001: data <= 32'hb0483464;
    11'b01011011010: data <= 32'hb60a3d0d;
    11'b01011011011: data <= 32'ha86c391e;
    11'b01011011100: data <= 32'h36e533e2;
    11'b01011011101: data <= 32'hb4d53c06;
    11'b01011011110: data <= 32'hbf8a3e89;
    11'b01011011111: data <= 32'hc0523b9d;
    11'b01011100000: data <= 32'hb368b2bd;
    11'b01011100001: data <= 32'h3fabb785;
    11'b01011100010: data <= 32'h40139766;
    11'b01011100011: data <= 32'h39ae3154;
    11'b01011100100: data <= 32'h333b2f87;
    11'b01011100101: data <= 32'h3c483940;
    11'b01011100110: data <= 32'h3db73d43;
    11'b01011100111: data <= 32'h33cb38c4;
    11'b01011101000: data <= 32'hbc76bde5;
    11'b01011101001: data <= 32'hbc1cc178;
    11'b01011101010: data <= 32'h2844bf1f;
    11'b01011101011: data <= 32'h3878ac9d;
    11'b01011101100: data <= 32'h355131ce;
    11'b01011101101: data <= 32'h3211b9ed;
    11'b01011101110: data <= 32'h2d38b99c;
    11'b01011101111: data <= 32'hbab03a9d;
    11'b01011110000: data <= 32'hc0633f87;
    11'b01011110001: data <= 32'hc0963c14;
    11'b01011110010: data <= 32'hb933b877;
    11'b01011110011: data <= 32'h3b38bb2d;
    11'b01011110100: data <= 32'h39cd200f;
    11'b01011110101: data <= 32'hb1ff3a16;
    11'b01011110110: data <= 32'h32133b8d;
    11'b01011110111: data <= 32'h3e8f3d05;
    11'b01011111000: data <= 32'h3fbb3e71;
    11'b01011111001: data <= 32'h34b13ba0;
    11'b01011111010: data <= 32'hbd1bb997;
    11'b01011111011: data <= 32'hbadcbec6;
    11'b01011111100: data <= 32'h3a18bc62;
    11'b01011111101: data <= 32'h3e1db3fd;
    11'b01011111110: data <= 32'h3c29b9b1;
    11'b01011111111: data <= 32'h377ebeaf;
    11'b01100000000: data <= 32'h3387bc82;
    11'b01100000001: data <= 32'hb6c43a68;
    11'b01100000010: data <= 32'hbe333ed1;
    11'b01100000011: data <= 32'hbfb33577;
    11'b01100000100: data <= 32'hbc3abdfe;
    11'b01100000101: data <= 32'hb369be36;
    11'b01100000110: data <= 32'hb80caeca;
    11'b01100000111: data <= 32'hbb053b6b;
    11'b01100001000: data <= 32'h2ddf3ba3;
    11'b01100001001: data <= 32'h3e763c1b;
    11'b01100001010: data <= 32'h3e083e2f;
    11'b01100001011: data <= 32'hb6f33e23;
    11'b01100001100: data <= 32'hbf113855;
    11'b01100001101: data <= 32'hb9f6b5aa;
    11'b01100001110: data <= 32'h3d20b533;
    11'b01100001111: data <= 32'h3fd6b2e9;
    11'b01100010000: data <= 32'h3ca8bbb9;
    11'b01100010001: data <= 32'h38ccbe97;
    11'b01100010010: data <= 32'h3ad4ba04;
    11'b01100010011: data <= 32'h3a193c40;
    11'b01100010100: data <= 32'hb4b73d98;
    11'b01100010101: data <= 32'hbd0db734;
    11'b01100010110: data <= 32'hbce3c084;
    11'b01100010111: data <= 32'hbaa7bfae;
    11'b01100011000: data <= 32'hbb6fb46c;
    11'b01100011001: data <= 32'hbb2f3751;
    11'b01100011010: data <= 32'h30071801;
    11'b01100011011: data <= 32'h3cda1f0c;
    11'b01100011100: data <= 32'h38ef3c7a;
    11'b01100011101: data <= 32'hbd643feb;
    11'b01100011110: data <= 32'hc0783dfe;
    11'b01100011111: data <= 32'hba853766;
    11'b01100100000: data <= 32'h3c7e2473;
    11'b01100100001: data <= 32'h3d94aebd;
    11'b01100100010: data <= 32'h37a9b8c6;
    11'b01100100011: data <= 32'h36fabad7;
    11'b01100100100: data <= 32'h3e3a2e81;
    11'b01100100101: data <= 32'h40043de3;
    11'b01100100110: data <= 32'h3a653d1a;
    11'b01100100111: data <= 32'hba01b96e;
    11'b01100101000: data <= 32'hbc7dc052;
    11'b01100101001: data <= 32'hb92cbe6b;
    11'b01100101010: data <= 32'hb665b52c;
    11'b01100101011: data <= 32'hb480b60c;
    11'b01100101100: data <= 32'h357fbd8a;
    11'b01100101101: data <= 32'h3adcbcd9;
    11'b01100101110: data <= 32'h279238d1;
    11'b01100101111: data <= 32'hbeb8401f;
    11'b01100110000: data <= 32'hc07e3e92;
    11'b01100110001: data <= 32'hbbca34eb;
    11'b01100110010: data <= 32'h3564b474;
    11'b01100110011: data <= 32'h2d18ad4e;
    11'b01100110100: data <= 32'hb981a752;
    11'b01100110101: data <= 32'h29a8a2cb;
    11'b01100110110: data <= 32'h3fb939c2;
    11'b01100110111: data <= 32'h412a3eba;
    11'b01100111000: data <= 32'h3c473dad;
    11'b01100111001: data <= 32'hb9e8aefb;
    11'b01100111010: data <= 32'hbb5fbc7d;
    11'b01100111011: data <= 32'h2856b94b;
    11'b01100111100: data <= 32'h3863b06e;
    11'b01100111101: data <= 32'h36fbbc3b;
    11'b01100111110: data <= 32'h3892c0c2;
    11'b01100111111: data <= 32'h3ac7bf8a;
    11'b01101000000: data <= 32'h343c35bf;
    11'b01101000001: data <= 32'hbc2f3f4c;
    11'b01101000010: data <= 32'hbe8c3c1a;
    11'b01101000011: data <= 32'hbc18b897;
    11'b01101000100: data <= 32'hb895bb6b;
    11'b01101000101: data <= 32'hbcdab179;
    11'b01101000110: data <= 32'hbe99340d;
    11'b01101000111: data <= 32'hb50830ab;
    11'b01101001000: data <= 32'h3f483816;
    11'b01101001001: data <= 32'h40743da3;
    11'b01101001010: data <= 32'h36fa3ea6;
    11'b01101001011: data <= 32'hbcc93b3c;
    11'b01101001100: data <= 32'hba5f3464;
    11'b01101001101: data <= 32'h39043669;
    11'b01101001110: data <= 32'h3c62323f;
    11'b01101001111: data <= 32'h38b8bcc8;
    11'b01101010000: data <= 32'h3841c0de;
    11'b01101010001: data <= 32'h3ca2be90;
    11'b01101010010: data <= 32'h3ce83871;
    11'b01101010011: data <= 32'h34273e09;
    11'b01101010100: data <= 32'hb964323f;
    11'b01101010101: data <= 32'hbadcbdae;
    11'b01101010110: data <= 32'hbc20bd51;
    11'b01101010111: data <= 32'hbee2b2bc;
    11'b01101011000: data <= 32'hbf5e2a87;
    11'b01101011001: data <= 32'hb62eb8c2;
    11'b01101011010: data <= 32'h3d9bb862;
    11'b01101011011: data <= 32'h3d4c3979;
    11'b01101011100: data <= 32'hb8463f05;
    11'b01101011101: data <= 32'hbecb3ec8;
    11'b01101011110: data <= 32'hba2c3cbb;
    11'b01101011111: data <= 32'h398e3ba9;
    11'b01101100000: data <= 32'h39d43756;
    11'b01101100001: data <= 32'hafcaba5f;
    11'b01101100010: data <= 32'h2d80be9d;
    11'b01101100011: data <= 32'h3e05ba1b;
    11'b01101100100: data <= 32'h40963bf5;
    11'b01101100101: data <= 32'h3dcd3d4a;
    11'b01101100110: data <= 32'h2de0b304;
    11'b01101100111: data <= 32'hb870be04;
    11'b01101101000: data <= 32'hba5cbc04;
    11'b01101101001: data <= 32'hbce99054;
    11'b01101101010: data <= 32'hbcf6b6fa;
    11'b01101101011: data <= 32'hb0dbbf2c;
    11'b01101101100: data <= 32'h3c05bf75;
    11'b01101101101: data <= 32'h38b5af86;
    11'b01101101110: data <= 32'hbc203e5a;
    11'b01101101111: data <= 32'hbee13f11;
    11'b01101110000: data <= 32'hb9a53c58;
    11'b01101110001: data <= 32'h339d39c7;
    11'b01101110010: data <= 32'hb65237da;
    11'b01101110011: data <= 32'hbd89b279;
    11'b01101110100: data <= 32'hb8e2b996;
    11'b01101110101: data <= 32'h3e5f1bd9;
    11'b01101110110: data <= 32'h41893cee;
    11'b01101110111: data <= 32'h3f313d1d;
    11'b01101111000: data <= 32'h32de29a7;
    11'b01101111001: data <= 32'hb4e5b944;
    11'b01101111010: data <= 32'haded271b;
    11'b01101111011: data <= 32'hb26437f9;
    11'b01101111100: data <= 32'hb655ba6c;
    11'b01101111101: data <= 32'h2fa0c158;
    11'b01101111110: data <= 32'h3ac4c144;
    11'b01101111111: data <= 32'h385cb82b;
    11'b01110000000: data <= 32'hb8b93d08;
    11'b01110000001: data <= 32'hbc263c7c;
    11'b01110000010: data <= 32'hb71c30fe;
    11'b01110000011: data <= 32'hb57fa5ef;
    11'b01110000100: data <= 32'hbe3e35a9;
    11'b01110000101: data <= 32'hc0ea3226;
    11'b01110000110: data <= 32'hbcb5b4a9;
    11'b01110000111: data <= 32'h3d5ea1b8;
    11'b01110001000: data <= 32'h40c03b47;
    11'b01110001001: data <= 32'h3c943ce6;
    11'b01110001010: data <= 32'hb4d739c8;
    11'b01110001011: data <= 32'hb32338d2;
    11'b01110001100: data <= 32'h38ad3cde;
    11'b01110001101: data <= 32'h38823c55;
    11'b01110001110: data <= 32'haa69ba0e;
    11'b01110001111: data <= 32'h2b4ec15a;
    11'b01110010000: data <= 32'h3b18c0cc;
    11'b01110010001: data <= 32'h3cb2b4f2;
    11'b01110010010: data <= 32'h388b3bba;
    11'b01110010011: data <= 32'h2bb23336;
    11'b01110010100: data <= 32'h205cbb01;
    11'b01110010101: data <= 32'hb89eb8e2;
    11'b01110010110: data <= 32'hc00534f7;
    11'b01110010111: data <= 32'hc163333d;
    11'b01110011000: data <= 32'hbd22b9ae;
    11'b01110011001: data <= 32'h3b58bb4c;
    11'b01110011010: data <= 32'h3dac2afc;
    11'b01110011011: data <= 32'h24a83c09;
    11'b01110011100: data <= 32'hbbd63d05;
    11'b01110011101: data <= 32'hb3253dc7;
    11'b01110011110: data <= 32'h3ad43f6a;
    11'b01110011111: data <= 32'h38043dbe;
    11'b01110100000: data <= 32'hb8beb516;
    11'b01110100001: data <= 32'hb809bf65;
    11'b01110100010: data <= 32'h3b55bd96;
    11'b01110100011: data <= 32'h3fd33493;
    11'b01110100100: data <= 32'h3ebb3a8a;
    11'b01110100101: data <= 32'h3b7eb5c1;
    11'b01110100110: data <= 32'h3754bcfe;
    11'b01110100111: data <= 32'hb42db771;
    11'b01110101000: data <= 32'hbde538e8;
    11'b01110101001: data <= 32'hc0012a6d;
    11'b01110101010: data <= 32'hbb5dbe6f;
    11'b01110101011: data <= 32'h3885c049;
    11'b01110101100: data <= 32'h384dbb0e;
    11'b01110101101: data <= 32'hba013920;
    11'b01110101110: data <= 32'hbcc33cd0;
    11'b01110101111: data <= 32'hadd03d39;
    11'b01110110000: data <= 32'h398b3e46;
    11'b01110110001: data <= 32'hb50d3d84;
    11'b01110110010: data <= 32'hbf0933a0;
    11'b01110110011: data <= 32'hbd67ba2d;
    11'b01110110100: data <= 32'h3a15b606;
    11'b01110110101: data <= 32'h408a39c9;
    11'b01110110110: data <= 32'h3ff539e3;
    11'b01110110111: data <= 32'h3c37b5f1;
    11'b01110111000: data <= 32'h3959b9ae;
    11'b01110111001: data <= 32'h36b93755;
    11'b01110111010: data <= 32'hb57e3d11;
    11'b01110111011: data <= 32'hbb6ea95e;
    11'b01110111100: data <= 32'hb724c096;
    11'b01110111101: data <= 32'h3656c1be;
    11'b01110111110: data <= 32'h33c1bd4c;
    11'b01110111111: data <= 32'hb8f434af;
    11'b01111000000: data <= 32'hb910386c;
    11'b01111000001: data <= 32'h352034a2;
    11'b01111000010: data <= 32'h367c38fc;
    11'b01111000011: data <= 32'hbd0b3c2f;
    11'b01111000100: data <= 32'hc19638f5;
    11'b01111000101: data <= 32'hbffdb06e;
    11'b01111000110: data <= 32'h36f0ad31;
    11'b01111000111: data <= 32'h3f5a3860;
    11'b01111001000: data <= 32'h3d0d3861;
    11'b01111001001: data <= 32'h35fb1c04;
    11'b01111001010: data <= 32'h389a34f3;
    11'b01111001011: data <= 32'h3c493e6f;
    11'b01111001100: data <= 32'h38fa3fdf;
    11'b01111001101: data <= 32'hb469304a;
    11'b01111001110: data <= 32'hb565c074;
    11'b01111001111: data <= 32'h353cc127;
    11'b01111010000: data <= 32'h388cbbee;
    11'b01111010001: data <= 32'h347a309a;
    11'b01111010010: data <= 32'h36b9b510;
    11'b01111010011: data <= 32'h3b5abb62;
    11'b01111010100: data <= 32'h359bb436;
    11'b01111010101: data <= 32'hbe703a7c;
    11'b01111010110: data <= 32'hc1f839df;
    11'b01111010111: data <= 32'hc00fb431;
    11'b01111011000: data <= 32'h2f24b9a5;
    11'b01111011001: data <= 32'h3b31b401;
    11'b01111011010: data <= 32'ha6823164;
    11'b01111011011: data <= 32'hb8b43510;
    11'b01111011100: data <= 32'h35ed3c17;
    11'b01111011101: data <= 32'h3d91406d;
    11'b01111011110: data <= 32'h3abd4098;
    11'b01111011111: data <= 32'hb8373829;
    11'b01111100000: data <= 32'hba8fbd9c;
    11'b01111100001: data <= 32'h3218bdb7;
    11'b01111100010: data <= 32'h3c65b032;
    11'b01111100011: data <= 32'h3cf6327e;
    11'b01111100100: data <= 32'h3d1fbb72;
    11'b01111100101: data <= 32'h3d98be40;
    11'b01111100110: data <= 32'h3956b6be;
    11'b01111100111: data <= 32'hbc3d3c08;
    11'b01111101000: data <= 32'hc05639b8;
    11'b01111101001: data <= 32'hbdb8bb1e;
    11'b01111101010: data <= 32'ha94bbf08;
    11'b01111101011: data <= 32'h1cc8bcb7;
    11'b01111101100: data <= 32'hbc32b474;
    11'b01111101101: data <= 32'hbc7432af;
    11'b01111101110: data <= 32'h35eb3ad0;
    11'b01111101111: data <= 32'h3d7c3f53;
    11'b01111110000: data <= 32'h34e54017;
    11'b01111110001: data <= 32'hbdf73b29;
    11'b01111110010: data <= 32'hbea1b522;
    11'b01111110011: data <= 32'had49b15a;
    11'b01111110100: data <= 32'h3d383907;
    11'b01111110101: data <= 32'h3df9347f;
    11'b01111110110: data <= 32'h3d4fbc3f;
    11'b01111110111: data <= 32'h3ddabd3e;
    11'b01111111000: data <= 32'h3ccb3474;
    11'b01111111001: data <= 32'h2cad3e95;
    11'b01111111010: data <= 32'hbaf23a20;
    11'b01111111011: data <= 32'hb90dbdb1;
    11'b01111111100: data <= 32'ha6f4c0d2;
    11'b01111111101: data <= 32'hb637be4f;
    11'b01111111110: data <= 32'hbcd5b84b;
    11'b01111111111: data <= 32'hba6cb557;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    