
module memory_rom_5(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbd69baab;
    11'b00000000001: data <= 32'hb9b2b671;
    11'b00000000010: data <= 32'h3a9938bf;
    11'b00000000011: data <= 32'h3b323e95;
    11'b00000000100: data <= 32'hbb363df4;
    11'b00000000101: data <= 32'hc0b434d9;
    11'b00000000110: data <= 32'hbf0bb2a6;
    11'b00000000111: data <= 32'haeae388d;
    11'b00000001000: data <= 32'h3a893c56;
    11'b00000001001: data <= 32'h3b622ff0;
    11'b00000001010: data <= 32'h3cd8bc07;
    11'b00000001011: data <= 32'h3e6ab55d;
    11'b00000001100: data <= 32'h3ca43e49;
    11'b00000001101: data <= 32'h2c834041;
    11'b00000001110: data <= 32'hb530361f;
    11'b00000001111: data <= 32'h341cbeb6;
    11'b00000010000: data <= 32'h3768c014;
    11'b00000010001: data <= 32'hb60dbcdc;
    11'b00000010010: data <= 32'hbb1fbaa9;
    11'b00000010011: data <= 32'h31abbbea;
    11'b00000010100: data <= 32'h3e3bb8ac;
    11'b00000010101: data <= 32'h3bef368f;
    11'b00000010110: data <= 32'hbd693a77;
    11'b00000010111: data <= 32'hc1b13500;
    11'b00000011000: data <= 32'hbffe2823;
    11'b00000011001: data <= 32'hb5143775;
    11'b00000011010: data <= 32'h31b73861;
    11'b00000011011: data <= 32'hb345b5cb;
    11'b00000011100: data <= 32'h2612bb31;
    11'b00000011101: data <= 32'h3c083649;
    11'b00000011110: data <= 32'h3d6440da;
    11'b00000011111: data <= 32'h39004152;
    11'b00000100000: data <= 32'ha2a0396c;
    11'b00000100001: data <= 32'h2f5fbcb0;
    11'b00000100010: data <= 32'h33c6bc74;
    11'b00000100011: data <= 32'hb01ab3a9;
    11'b00000100100: data <= 32'ha8afb713;
    11'b00000100101: data <= 32'h3cd4bdc6;
    11'b00000100110: data <= 32'h4078bdfa;
    11'b00000100111: data <= 32'h3cf4b4b8;
    11'b00000101000: data <= 32'hbc8938f6;
    11'b00000101001: data <= 32'hc0a235a0;
    11'b00000101010: data <= 32'hbd76b3cd;
    11'b00000101011: data <= 32'hb1bcb56e;
    11'b00000101100: data <= 32'hb82ab722;
    11'b00000101101: data <= 32'hbdc1bbf9;
    11'b00000101110: data <= 32'hbbeabbdc;
    11'b00000101111: data <= 32'h38f43847;
    11'b00000110000: data <= 32'h3d7640be;
    11'b00000110001: data <= 32'h37c640de;
    11'b00000110010: data <= 32'hb8dc3a34;
    11'b00000110011: data <= 32'hb961b575;
    11'b00000110100: data <= 32'hb27633c6;
    11'b00000110101: data <= 32'h27363b75;
    11'b00000110110: data <= 32'h37681662;
    11'b00000110111: data <= 32'h3e5dbe6a;
    11'b00000111000: data <= 32'h40bfbea4;
    11'b00000111001: data <= 32'h3dfeaa21;
    11'b00000111010: data <= 32'hb5303c71;
    11'b00000111011: data <= 32'hbc1f386f;
    11'b00000111100: data <= 32'hb374b924;
    11'b00000111101: data <= 32'h31d2bc82;
    11'b00000111110: data <= 32'hbb6bbc8f;
    11'b00000111111: data <= 32'hc007bd75;
    11'b00001000000: data <= 32'hbcb2bd19;
    11'b00001000001: data <= 32'h3a59ae64;
    11'b00001000010: data <= 32'h3d843d67;
    11'b00001000011: data <= 32'hab323e21;
    11'b00001000100: data <= 32'hbe3838e4;
    11'b00001000101: data <= 32'hbe0d356d;
    11'b00001000110: data <= 32'hb8ec3ce1;
    11'b00001000111: data <= 32'hb03e3e27;
    11'b00001001000: data <= 32'h30502e63;
    11'b00001001001: data <= 32'h3ba9be32;
    11'b00001001010: data <= 32'h3f46bc9e;
    11'b00001001011: data <= 32'h3e5d3afc;
    11'b00001001100: data <= 32'h38b63fbd;
    11'b00001001101: data <= 32'h33883ae8;
    11'b00001001110: data <= 32'h3969b9fb;
    11'b00001001111: data <= 32'h3727bccc;
    11'b00001010000: data <= 32'hbb86bb7c;
    11'b00001010001: data <= 32'hbef3bca1;
    11'b00001010010: data <= 32'hb7b6be5c;
    11'b00001010011: data <= 32'h3dd1bc98;
    11'b00001010100: data <= 32'h3e06a84a;
    11'b00001010101: data <= 32'hb782381c;
    11'b00001010110: data <= 32'hc0173566;
    11'b00001010111: data <= 32'hbed63859;
    11'b00001011000: data <= 32'hb9573d3c;
    11'b00001011001: data <= 32'hb8553ceb;
    11'b00001011010: data <= 32'hbb2cb4a3;
    11'b00001011011: data <= 32'hb5dbbdf0;
    11'b00001011100: data <= 32'h3b13b804;
    11'b00001011101: data <= 32'h3de43ec7;
    11'b00001011110: data <= 32'h3c5640df;
    11'b00001011111: data <= 32'h39f03c2d;
    11'b00001100000: data <= 32'h3a5eb6c9;
    11'b00001100001: data <= 32'h35aeb604;
    11'b00001100010: data <= 32'hb9e33134;
    11'b00001100011: data <= 32'hbbefb711;
    11'b00001100100: data <= 32'h37ccbeea;
    11'b00001100101: data <= 32'h4036bfeb;
    11'b00001100110: data <= 32'h3ebbbb7b;
    11'b00001100111: data <= 32'hb62127fd;
    11'b00001101000: data <= 32'hbe6532b8;
    11'b00001101001: data <= 32'hbbc134dd;
    11'b00001101010: data <= 32'hb34f3919;
    11'b00001101011: data <= 32'hbb71353e;
    11'b00001101100: data <= 32'hc009bb3a;
    11'b00001101101: data <= 32'hbe4dbe28;
    11'b00001101110: data <= 32'h318ab462;
    11'b00001101111: data <= 32'h3d223ed3;
    11'b00001110000: data <= 32'h3bb7403f;
    11'b00001110001: data <= 32'h34db3afe;
    11'b00001110010: data <= 32'h30522f4f;
    11'b00001110011: data <= 32'habcf3b16;
    11'b00001110100: data <= 32'hb8a93e1c;
    11'b00001110101: data <= 32'hb7383587;
    11'b00001110110: data <= 32'h3b5bbe94;
    11'b00001110111: data <= 32'h405dc04a;
    11'b00001111000: data <= 32'h3eddbae6;
    11'b00001111001: data <= 32'h311e35b0;
    11'b00001111010: data <= 32'hb67b35d2;
    11'b00001111011: data <= 32'h35a2ac7a;
    11'b00001111100: data <= 32'h37cdb0cc;
    11'b00001111101: data <= 32'hbc43b655;
    11'b00001111110: data <= 32'hc126bced;
    11'b00001111111: data <= 32'hbfccbe9b;
    11'b00010000000: data <= 32'h307eb968;
    11'b00010000001: data <= 32'h3cdf3a33;
    11'b00010000010: data <= 32'h374d3c2c;
    11'b00010000011: data <= 32'hb8d835ac;
    11'b00010000100: data <= 32'hb9b2380b;
    11'b00010000101: data <= 32'hb7463f54;
    11'b00010000110: data <= 32'hb8e940ad;
    11'b00010000111: data <= 32'hb8ad3988;
    11'b00010001000: data <= 32'h35f9bde7;
    11'b00010001001: data <= 32'h3de0beb1;
    11'b00010001010: data <= 32'h3ddca1cd;
    11'b00010001011: data <= 32'h3a353ca2;
    11'b00010001100: data <= 32'h3a8f394f;
    11'b00010001101: data <= 32'h3decb426;
    11'b00010001110: data <= 32'h3c29b602;
    11'b00010001111: data <= 32'hbb6ab464;
    11'b00010010000: data <= 32'hc0a7bb26;
    11'b00010010001: data <= 32'hbd6dbe99;
    11'b00010010010: data <= 32'h39f9bdb8;
    11'b00010010011: data <= 32'h3d57b87d;
    11'b00010010100: data <= 32'h9d15b296;
    11'b00010010101: data <= 32'hbcd7b3c8;
    11'b00010010110: data <= 32'hbbe0382b;
    11'b00010010111: data <= 32'hb6843fc6;
    11'b00010011000: data <= 32'hb9ef4052;
    11'b00010011001: data <= 32'hbd57364f;
    11'b00010011010: data <= 32'hbb2abd91;
    11'b00010011011: data <= 32'h34d6bbff;
    11'b00010011100: data <= 32'h3bf73b1a;
    11'b00010011101: data <= 32'h3c323eea;
    11'b00010011110: data <= 32'h3d603a34;
    11'b00010011111: data <= 32'h3f0db18e;
    11'b00010100000: data <= 32'h3c573210;
    11'b00010100001: data <= 32'hb9763a1b;
    11'b00010100010: data <= 32'hbe5029d7;
    11'b00010100011: data <= 32'hb581bdb2;
    11'b00010100100: data <= 32'h3dd3c006;
    11'b00010100101: data <= 32'h3de0bde4;
    11'b00010100110: data <= 32'haf35bb0f;
    11'b00010100111: data <= 32'hbbf7b877;
    11'b00010101000: data <= 32'hb4f732dc;
    11'b00010101001: data <= 32'h339a3d22;
    11'b00010101010: data <= 32'hba273cff;
    11'b00010101011: data <= 32'hc062b426;
    11'b00010101100: data <= 32'hc037bdb2;
    11'b00010101101: data <= 32'hb90bb8f3;
    11'b00010101110: data <= 32'h388b3c6b;
    11'b00010101111: data <= 32'h3a9f3df2;
    11'b00010110000: data <= 32'h3b6736cb;
    11'b00010110001: data <= 32'h3c8624e4;
    11'b00010110010: data <= 32'h393f3cbb;
    11'b00010110011: data <= 32'hb8294041;
    11'b00010110100: data <= 32'hbb613c4c;
    11'b00010110101: data <= 32'h344abc3a;
    11'b00010110110: data <= 32'h3e73c015;
    11'b00010110111: data <= 32'h3d69bdb4;
    11'b00010111000: data <= 32'h2efdb909;
    11'b00010111001: data <= 32'hac51b6d8;
    11'b00010111010: data <= 32'h3c05b161;
    11'b00010111011: data <= 32'h3cd436a0;
    11'b00010111100: data <= 32'hb8b235f9;
    11'b00010111101: data <= 32'hc129b965;
    11'b00010111110: data <= 32'hc106bdb0;
    11'b00010111111: data <= 32'hba37b9d7;
    11'b00011000000: data <= 32'h36ef36ea;
    11'b00011000001: data <= 32'h34cb36ba;
    11'b00011000010: data <= 32'ha8e3b5a2;
    11'b00011000011: data <= 32'h31372c6e;
    11'b00011000100: data <= 32'h31883fbd;
    11'b00011000101: data <= 32'hb78a41f2;
    11'b00011000110: data <= 32'hba683e4e;
    11'b00011000111: data <= 32'ha730ba23;
    11'b00011001000: data <= 32'h3b66be1c;
    11'b00011001001: data <= 32'h3ad2b856;
    11'b00011001010: data <= 32'h35f53427;
    11'b00011001011: data <= 32'h3b92aa06;
    11'b00011001100: data <= 32'h4059b68a;
    11'b00011001101: data <= 32'h3fd2a759;
    11'b00011001110: data <= 32'hb4673418;
    11'b00011001111: data <= 32'hc088b61c;
    11'b00011010000: data <= 32'hbf9ebcc4;
    11'b00011010001: data <= 32'hafe6bc86;
    11'b00011010010: data <= 32'h38e4b970;
    11'b00011010011: data <= 32'hb237bafa;
    11'b00011010100: data <= 32'hba98bcb8;
    11'b00011010101: data <= 32'hb557b05c;
    11'b00011010110: data <= 32'h30f73fd2;
    11'b00011010111: data <= 32'hb66c4197;
    11'b00011011000: data <= 32'hbcd63d19;
    11'b00011011001: data <= 32'hbc41b9b8;
    11'b00011011010: data <= 32'hb487baa1;
    11'b00011011011: data <= 32'h30073810;
    11'b00011011100: data <= 32'h36153c25;
    11'b00011011101: data <= 32'h3d6b30ae;
    11'b00011011110: data <= 32'h40f4b7c4;
    11'b00011011111: data <= 32'h401732e2;
    11'b00011100000: data <= 32'ha6523c38;
    11'b00011100001: data <= 32'hbdf638b6;
    11'b00011100010: data <= 32'hba24b98e;
    11'b00011100011: data <= 32'h3a2ebda8;
    11'b00011100100: data <= 32'h3ab4bdd2;
    11'b00011100101: data <= 32'hb6e4be5d;
    11'b00011100110: data <= 32'hbb40be5f;
    11'b00011100111: data <= 32'h2e57b7ef;
    11'b00011101000: data <= 32'h3a863d0b;
    11'b00011101001: data <= 32'hb1123f26;
    11'b00011101010: data <= 32'hbefa375d;
    11'b00011101011: data <= 32'hc03dbabe;
    11'b00011101100: data <= 32'hbd1ab591;
    11'b00011101101: data <= 32'hb73c3bf8;
    11'b00011101110: data <= 32'h2b0a3c26;
    11'b00011101111: data <= 32'h3b22b25d;
    11'b00011110000: data <= 32'h3f1cb866;
    11'b00011110001: data <= 32'h3df43b02;
    11'b00011110010: data <= 32'h2a27407e;
    11'b00011110011: data <= 32'hba0f3ec0;
    11'b00011110100: data <= 32'h2dddb032;
    11'b00011110101: data <= 32'h3cb0bd25;
    11'b00011110110: data <= 32'h3a01bd63;
    11'b00011110111: data <= 32'hb71ebd33;
    11'b00011111000: data <= 32'hb4f6bd86;
    11'b00011111001: data <= 32'h3cecba74;
    11'b00011111010: data <= 32'h3f70354f;
    11'b00011111011: data <= 32'h34193982;
    11'b00011111100: data <= 32'hbfb8b257;
    11'b00011111101: data <= 32'hc0e5bb29;
    11'b00011111110: data <= 32'hbda8b3fa;
    11'b00011111111: data <= 32'hb8783935;
    11'b00100000000: data <= 32'hb6eb3155;
    11'b00100000001: data <= 32'hafd5bc31;
    11'b00100000010: data <= 32'h38e6ba0d;
    11'b00100000011: data <= 32'h3a283d8f;
    11'b00100000100: data <= 32'h251e4201;
    11'b00100000101: data <= 32'hb748406d;
    11'b00100000110: data <= 32'h2f663203;
    11'b00100000111: data <= 32'h398fba2f;
    11'b00100001000: data <= 32'h3210b6a4;
    11'b00100001001: data <= 32'hb736b3d3;
    11'b00100001010: data <= 32'h3700ba40;
    11'b00100001011: data <= 32'h4098bba4;
    11'b00100001100: data <= 32'h4151b436;
    11'b00100001101: data <= 32'h3939342e;
    11'b00100001110: data <= 32'hbe48b03c;
    11'b00100001111: data <= 32'hbf28b8fe;
    11'b00100010000: data <= 32'hb903b614;
    11'b00100010001: data <= 32'hb21eb193;
    11'b00100010010: data <= 32'hbaa7bc0e;
    11'b00100010011: data <= 32'hbc24bfd0;
    11'b00100010100: data <= 32'hb1c7bc66;
    11'b00100010101: data <= 32'h38123d49;
    11'b00100010110: data <= 32'h2e7f418a;
    11'b00100010111: data <= 32'hb8d23f3f;
    11'b00100011000: data <= 32'hb8f12dc2;
    11'b00100011001: data <= 32'hb632b10f;
    11'b00100011010: data <= 32'hb90d39f4;
    11'b00100011011: data <= 32'hb9043a80;
    11'b00100011100: data <= 32'h39bbb558;
    11'b00100011101: data <= 32'h4117bc0d;
    11'b00100011110: data <= 32'h4161b431;
    11'b00100011111: data <= 32'h3a6839fb;
    11'b00100100000: data <= 32'hbae0398c;
    11'b00100100001: data <= 32'hb86fa6e8;
    11'b00100100010: data <= 32'h383eb70f;
    11'b00100100011: data <= 32'h34afba41;
    11'b00100100100: data <= 32'hbc18beb5;
    11'b00100100101: data <= 32'hbd5ac0b2;
    11'b00100100110: data <= 32'hac31bda4;
    11'b00100100111: data <= 32'h3c02394f;
    11'b00100101000: data <= 32'h37003eb3;
    11'b00100101001: data <= 32'hbb223a12;
    11'b00100101010: data <= 32'hbde5b4a4;
    11'b00100101011: data <= 32'hbd493427;
    11'b00100101100: data <= 32'hbcf13dbb;
    11'b00100101101: data <= 32'hbbb43c88;
    11'b00100101110: data <= 32'h341db7cf;
    11'b00100101111: data <= 32'h3f12bc9d;
    11'b00100110000: data <= 32'h3fb2308e;
    11'b00100110001: data <= 32'h39183ed9;
    11'b00100110010: data <= 32'hb2653eea;
    11'b00100110011: data <= 32'h37d038ca;
    11'b00100110100: data <= 32'h3d02b3d2;
    11'b00100110101: data <= 32'h36bcb924;
    11'b00100110110: data <= 32'hbc5cbd47;
    11'b00100110111: data <= 32'hbc00bfde;
    11'b00100111000: data <= 32'h3a87be0d;
    11'b00100111001: data <= 32'h3fe2b219;
    11'b00100111010: data <= 32'h3b853683;
    11'b00100111011: data <= 32'hbba7b317;
    11'b00100111100: data <= 32'hbeeeb8a5;
    11'b00100111101: data <= 32'hbd9f3627;
    11'b00100111110: data <= 32'hbce13d5e;
    11'b00100111111: data <= 32'hbd223841;
    11'b00101000000: data <= 32'hb984bcfc;
    11'b00101000001: data <= 32'h3735bdd9;
    11'b00101000010: data <= 32'h3b1d37e6;
    11'b00101000011: data <= 32'h35a240bb;
    11'b00101000100: data <= 32'h2e98406a;
    11'b00101000101: data <= 32'h3a163ac3;
    11'b00101000110: data <= 32'h3c4130e7;
    11'b00101000111: data <= 32'ha70e33a2;
    11'b00101001000: data <= 32'hbccfb018;
    11'b00101001001: data <= 32'hb725bc46;
    11'b00101001010: data <= 32'h3f03bd96;
    11'b00101001011: data <= 32'h4177ba1a;
    11'b00101001100: data <= 32'h3d40b42c;
    11'b00101001101: data <= 32'hb943b771;
    11'b00101001110: data <= 32'hbc69b738;
    11'b00101001111: data <= 32'hb7fa35ac;
    11'b00101010000: data <= 32'hb8a439df;
    11'b00101010001: data <= 32'hbdb1b7e4;
    11'b00101010010: data <= 32'hbe41c03d;
    11'b00101010011: data <= 32'hb896bf4d;
    11'b00101010100: data <= 32'h34cf36e8;
    11'b00101010101: data <= 32'h34244047;
    11'b00101010110: data <= 32'h29423ed2;
    11'b00101010111: data <= 32'h342f3818;
    11'b00101011000: data <= 32'h31403839;
    11'b00101011001: data <= 32'hba883d67;
    11'b00101011010: data <= 32'hbdbf3c98;
    11'b00101011011: data <= 32'hb2bcb47c;
    11'b00101011100: data <= 32'h3fefbcfc;
    11'b00101011101: data <= 32'h415dba9a;
    11'b00101011110: data <= 32'h3d13a50c;
    11'b00101011111: data <= 32'hb0f830c4;
    11'b00101100000: data <= 32'h2d892e9e;
    11'b00101100001: data <= 32'h3af0360f;
    11'b00101100010: data <= 32'h33f332d9;
    11'b00101100011: data <= 32'hbd86bc77;
    11'b00101100100: data <= 32'hbfa0c0ea;
    11'b00101100101: data <= 32'hb9afbffa;
    11'b00101100110: data <= 32'h3866ab15;
    11'b00101100111: data <= 32'h383e3c53;
    11'b00101101000: data <= 32'hb0b23751;
    11'b00101101001: data <= 32'hb77ab2a8;
    11'b00101101010: data <= 32'hb9ab3992;
    11'b00101101011: data <= 32'hbd8b401f;
    11'b00101101100: data <= 32'hbebc3ee7;
    11'b00101101101: data <= 32'hb858b11e;
    11'b00101101110: data <= 32'h3cf1bd2b;
    11'b00101101111: data <= 32'h3ef6b832;
    11'b00101110000: data <= 32'h3a3e3a47;
    11'b00101110001: data <= 32'h33fc3c63;
    11'b00101110010: data <= 32'h3c8c39b1;
    11'b00101110011: data <= 32'h3f653851;
    11'b00101110100: data <= 32'h39713463;
    11'b00101110101: data <= 32'hbd47ba41;
    11'b00101110110: data <= 32'hbea9bfb4;
    11'b00101110111: data <= 32'ha37abf33;
    11'b00101111000: data <= 32'h3d9eb949;
    11'b00101111001: data <= 32'h3c17b1f1;
    11'b00101111010: data <= 32'hb27dba49;
    11'b00101111011: data <= 32'hba10baa1;
    11'b00101111100: data <= 32'hba723949;
    11'b00101111101: data <= 32'hbd01401c;
    11'b00101111110: data <= 32'hbefd3d54;
    11'b00101111111: data <= 32'hbd07ba2e;
    11'b00110000000: data <= 32'hacc9be59;
    11'b00110000001: data <= 32'h371db2eb;
    11'b00110000010: data <= 32'h30a33db4;
    11'b00110000011: data <= 32'h35c93e4f;
    11'b00110000100: data <= 32'h3df03afa;
    11'b00110000101: data <= 32'h3f8e39d6;
    11'b00110000110: data <= 32'h36973b99;
    11'b00110000111: data <= 32'hbd9e3662;
    11'b00110001000: data <= 32'hbcb5ba34;
    11'b00110001001: data <= 32'h3afcbd4a;
    11'b00110001010: data <= 32'h404fbc11;
    11'b00110001011: data <= 32'h3d5bbb58;
    11'b00110001100: data <= 32'hab87bd1f;
    11'b00110001101: data <= 32'hb4c6bb58;
    11'b00110001110: data <= 32'h2dab38a6;
    11'b00110001111: data <= 32'hb6143e1d;
    11'b00110010000: data <= 32'hbe1f363e;
    11'b00110010001: data <= 32'hbf99be79;
    11'b00110010010: data <= 32'hbc9cbfad;
    11'b00110010011: data <= 32'hb6a4b18e;
    11'b00110010100: data <= 32'hb2b53d55;
    11'b00110010101: data <= 32'h33153c5b;
    11'b00110010110: data <= 32'h3c4c3558;
    11'b00110010111: data <= 32'h3c6c3a25;
    11'b00110011000: data <= 32'hb5443f4e;
    11'b00110011001: data <= 32'hbe813ee3;
    11'b00110011010: data <= 32'hbb0e34c3;
    11'b00110011011: data <= 32'h3ccebaf9;
    11'b00110011100: data <= 32'h403dbbbe;
    11'b00110011101: data <= 32'h3c7eba28;
    11'b00110011110: data <= 32'h306dba8a;
    11'b00110011111: data <= 32'h394eb70a;
    11'b00110100000: data <= 32'h3df938d1;
    11'b00110100001: data <= 32'h39ee3bea;
    11'b00110100010: data <= 32'hbca0b4c6;
    11'b00110100011: data <= 32'hc032bfe7;
    11'b00110100100: data <= 32'hbd87bfcf;
    11'b00110100101: data <= 32'hb5a3b64f;
    11'b00110100110: data <= 32'haaae37cd;
    11'b00110100111: data <= 32'h26dcb227;
    11'b00110101000: data <= 32'h35c1b96b;
    11'b00110101001: data <= 32'h327838ad;
    11'b00110101010: data <= 32'hbb5c40bb;
    11'b00110101011: data <= 32'hbf1a40c7;
    11'b00110101100: data <= 32'hbbf0391d;
    11'b00110101101: data <= 32'h392fba12;
    11'b00110101110: data <= 32'h3c9bb928;
    11'b00110101111: data <= 32'h35a89cc8;
    11'b00110110000: data <= 32'h31e83009;
    11'b00110110001: data <= 32'h3e1a31ec;
    11'b00110110010: data <= 32'h4121399d;
    11'b00110110011: data <= 32'h3db43afc;
    11'b00110110100: data <= 32'hbb1eb05f;
    11'b00110110101: data <= 32'hbf3fbdb8;
    11'b00110110110: data <= 32'hb9f2bdfd;
    11'b00110110111: data <= 32'h375eb92b;
    11'b00110111000: data <= 32'h3714b8a8;
    11'b00110111001: data <= 32'hac02be1a;
    11'b00110111010: data <= 32'habcfbe50;
    11'b00110111011: data <= 32'ha9d534cd;
    11'b00110111100: data <= 32'hba4d4094;
    11'b00110111101: data <= 32'hbe714021;
    11'b00110111110: data <= 32'hbd792ee0;
    11'b00110111111: data <= 32'hb765bc20;
    11'b00111000000: data <= 32'hb379b51b;
    11'b00111000001: data <= 32'hb8af39cf;
    11'b00111000010: data <= 32'h207a39db;
    11'b00111000011: data <= 32'h3f1c35d2;
    11'b00111000100: data <= 32'h4160399f;
    11'b00111000101: data <= 32'h3d1d3cf5;
    11'b00111000110: data <= 32'hbb5c3ac1;
    11'b00111000111: data <= 32'hbd3db24f;
    11'b00111001000: data <= 32'h3261b9a0;
    11'b00111001001: data <= 32'h3d3db976;
    11'b00111001010: data <= 32'h3a4fbcc9;
    11'b00111001011: data <= 32'hac36c03d;
    11'b00111001100: data <= 32'h2ffabf57;
    11'b00111001101: data <= 32'h393c300a;
    11'b00111001110: data <= 32'h30ea3efb;
    11'b00111001111: data <= 32'hbc503c63;
    11'b00111010000: data <= 32'hbeafba79;
    11'b00111010001: data <= 32'hbd9ebd97;
    11'b00111010010: data <= 32'hbcd2b158;
    11'b00111010011: data <= 32'hbc9c3af2;
    11'b00111010100: data <= 32'hb45836e0;
    11'b00111010101: data <= 32'h3d5cb33e;
    11'b00111010110: data <= 32'h3fa03710;
    11'b00111010111: data <= 32'h37fc3f14;
    11'b00111011000: data <= 32'hbcb14008;
    11'b00111011001: data <= 32'hbb7e3bfd;
    11'b00111011010: data <= 32'h39d01af0;
    11'b00111011011: data <= 32'h3dcdb71f;
    11'b00111011100: data <= 32'h3854bc07;
    11'b00111011101: data <= 32'hb08bbebe;
    11'b00111011110: data <= 32'h39f7bd6d;
    11'b00111011111: data <= 32'h3f993151;
    11'b00111100000: data <= 32'h3d9a3c9a;
    11'b00111100001: data <= 32'hb69f33c9;
    11'b00111100010: data <= 32'hbe8bbd54;
    11'b00111100011: data <= 32'hbe4cbdb0;
    11'b00111100100: data <= 32'hbccdb0b4;
    11'b00111100101: data <= 32'hbc2d3591;
    11'b00111100110: data <= 32'hb789b980;
    11'b00111100111: data <= 32'h38b1bd73;
    11'b00111101000: data <= 32'h3af6ab0c;
    11'b00111101001: data <= 32'hb3df4013;
    11'b00111101010: data <= 32'hbd584137;
    11'b00111101011: data <= 32'hbabc3db2;
    11'b00111101100: data <= 32'h37a632f8;
    11'b00111101101: data <= 32'h3934ad38;
    11'b00111101110: data <= 32'hb583b2c1;
    11'b00111101111: data <= 32'hb6b2b923;
    11'b00111110000: data <= 32'h3d3fb8c4;
    11'b00111110001: data <= 32'h41c334c4;
    11'b00111110010: data <= 32'h40633aef;
    11'b00111110011: data <= 32'h1fa82fd2;
    11'b00111110100: data <= 32'hbd0fbbb0;
    11'b00111110101: data <= 32'hbb3dbaf0;
    11'b00111110110: data <= 32'hb527acf9;
    11'b00111110111: data <= 32'hb70eb690;
    11'b00111111000: data <= 32'hb828bfb2;
    11'b00111111001: data <= 32'h2832c0ca;
    11'b00111111010: data <= 32'h35d3b85b;
    11'b00111111011: data <= 32'hb4b53f55;
    11'b00111111100: data <= 32'hbc62407f;
    11'b00111111101: data <= 32'hbb493ae4;
    11'b00111111110: data <= 32'hb502b003;
    11'b00111111111: data <= 32'hb90932a3;
    11'b01000000000: data <= 32'hbdba38fe;
    11'b01000000001: data <= 32'hbac0323f;
    11'b01000000010: data <= 32'h3d93b368;
    11'b01000000011: data <= 32'h41ee3410;
    11'b01000000100: data <= 32'h401b3b98;
    11'b01000000101: data <= 32'haa1d3a44;
    11'b01000000110: data <= 32'hba453102;
    11'b01000000111: data <= 32'h2fd02d6c;
    11'b01000001000: data <= 32'h39d83177;
    11'b01000001001: data <= 32'h2dc2ba8d;
    11'b01000001010: data <= 32'hb84ec0f2;
    11'b01000001011: data <= 32'ha868c163;
    11'b01000001100: data <= 32'h39feb9f4;
    11'b01000001101: data <= 32'h38233d21;
    11'b01000001110: data <= 32'hb68b3cd6;
    11'b01000001111: data <= 32'hbb3ab359;
    11'b01000010000: data <= 32'hbc12b958;
    11'b01000010001: data <= 32'hbe3935a0;
    11'b01000010010: data <= 32'hc02a3be5;
    11'b01000010011: data <= 32'hbcd33254;
    11'b01000010100: data <= 32'h3b5bb968;
    11'b01000010101: data <= 32'h403eb0b9;
    11'b01000010110: data <= 32'h3c843ca3;
    11'b01000010111: data <= 32'hb75d3ec6;
    11'b01000011000: data <= 32'hb6ec3d36;
    11'b01000011001: data <= 32'h3aba3b4b;
    11'b01000011010: data <= 32'h3ca83861;
    11'b01000011011: data <= 32'h1ca1b874;
    11'b01000011100: data <= 32'hb9d8bff4;
    11'b01000011101: data <= 32'h3454c038;
    11'b01000011110: data <= 32'h3eddb892;
    11'b01000011111: data <= 32'h3ed539bc;
    11'b01000100000: data <= 32'h367c3206;
    11'b01000100001: data <= 32'hb967bc22;
    11'b01000100010: data <= 32'hbc51baf5;
    11'b01000100011: data <= 32'hbe0a375d;
    11'b01000100100: data <= 32'hbfa63a28;
    11'b01000100101: data <= 32'hbd3eb90d;
    11'b01000100110: data <= 32'h3219befa;
    11'b01000100111: data <= 32'h3b84ba7c;
    11'b01000101000: data <= 32'h2f8c3cc4;
    11'b01000101001: data <= 32'hba824048;
    11'b01000101010: data <= 32'hb4713ec9;
    11'b01000101011: data <= 32'h3b073c75;
    11'b01000101100: data <= 32'h39463aed;
    11'b01000101101: data <= 32'hba673349;
    11'b01000101110: data <= 32'hbcb8ba8f;
    11'b01000101111: data <= 32'h388cbc69;
    11'b01000110000: data <= 32'h410cb3cb;
    11'b01000110001: data <= 32'h40f43664;
    11'b01000110010: data <= 32'h3ae9b266;
    11'b01000110011: data <= 32'hb4b2bbb4;
    11'b01000110100: data <= 32'hb662b6a1;
    11'b01000110101: data <= 32'hb8353994;
    11'b01000110110: data <= 32'hbc5e34cb;
    11'b01000110111: data <= 32'hbcaabeae;
    11'b01000111000: data <= 32'hb5fcc184;
    11'b01000111001: data <= 32'h31f5bd88;
    11'b01000111010: data <= 32'hb39e3b59;
    11'b01000111011: data <= 32'hb9933efa;
    11'b01000111100: data <= 32'hb22f3c30;
    11'b01000111101: data <= 32'h362d38bd;
    11'b01000111110: data <= 32'hb6763bd8;
    11'b01000111111: data <= 32'hbf7d3c3d;
    11'b01001000000: data <= 32'hbee833d2;
    11'b01001000001: data <= 32'h383cb6d7;
    11'b01001000010: data <= 32'h4116b05a;
    11'b01001000011: data <= 32'h4088359d;
    11'b01001000100: data <= 32'h3968310f;
    11'b01001000101: data <= 32'h29bbad46;
    11'b01001000110: data <= 32'h38f83825;
    11'b01001000111: data <= 32'h39dd3c64;
    11'b01001001000: data <= 32'hb4102b6b;
    11'b01001001001: data <= 32'hbc0ac043;
    11'b01001001010: data <= 32'hb85bc205;
    11'b01001001011: data <= 32'h3455be00;
    11'b01001001100: data <= 32'h35103785;
    11'b01001001101: data <= 32'ha95439a6;
    11'b01001001110: data <= 32'ha309b365;
    11'b01001001111: data <= 32'haf2cb3e2;
    11'b01001010000: data <= 32'hbce23b77;
    11'b01001010001: data <= 32'hc0ff3dff;
    11'b01001010010: data <= 32'hc01e3852;
    11'b01001010011: data <= 32'h2f15b8c1;
    11'b01001010100: data <= 32'h3ec3b7bd;
    11'b01001010101: data <= 32'h3cb53622;
    11'b01001010110: data <= 32'ha2c63aa4;
    11'b01001010111: data <= 32'h32693b77;
    11'b01001011000: data <= 32'h3d953d5d;
    11'b01001011001: data <= 32'h3dcd3e00;
    11'b01001011010: data <= 32'ha999350a;
    11'b01001011011: data <= 32'hbc7bbe80;
    11'b01001011100: data <= 32'hb693c091;
    11'b01001011101: data <= 32'h3bd0bc51;
    11'b01001011110: data <= 32'h3d6a2df0;
    11'b01001011111: data <= 32'h3a3fb5b4;
    11'b01001100000: data <= 32'h34a5bd3d;
    11'b01001100001: data <= 32'hb015ba12;
    11'b01001100010: data <= 32'hbc903b71;
    11'b01001100011: data <= 32'hc06e3dc0;
    11'b01001100100: data <= 32'hbfd4a319;
    11'b01001100101: data <= 32'hb726bdf1;
    11'b01001100110: data <= 32'h3799bca1;
    11'b01001100111: data <= 32'hae6434c6;
    11'b01001101000: data <= 32'hb9833cbc;
    11'b01001101001: data <= 32'h32ea3d1e;
    11'b01001101010: data <= 32'h3e493ddc;
    11'b01001101011: data <= 32'h3cec3ea7;
    11'b01001101100: data <= 32'hb92b3ba5;
    11'b01001101101: data <= 32'hbe4ab6da;
    11'b01001101110: data <= 32'hb41abc19;
    11'b01001101111: data <= 32'h3e99b6cb;
    11'b01001110000: data <= 32'h401fabed;
    11'b01001110001: data <= 32'h3cc7baee;
    11'b01001110010: data <= 32'h3896be22;
    11'b01001110011: data <= 32'h3725b844;
    11'b01001110100: data <= 32'hb0323c9e;
    11'b01001110101: data <= 32'hbca93c82;
    11'b01001110110: data <= 32'hbdf8bb10;
    11'b01001110111: data <= 32'hbaaac0d8;
    11'b01001111000: data <= 32'hb624bedb;
    11'b01001111001: data <= 32'hba122c49;
    11'b01001111010: data <= 32'hbaa93acc;
    11'b01001111011: data <= 32'h343c38d4;
    11'b01001111100: data <= 32'h3cfb39ef;
    11'b01001111101: data <= 32'h35d93de9;
    11'b01001111110: data <= 32'hbe813e6a;
    11'b01001111111: data <= 32'hc04039d0;
    11'b01010000000: data <= 32'hb4e6a93f;
    11'b01010000001: data <= 32'h3ec0a6c6;
    11'b01010000010: data <= 32'h3f4aa9d8;
    11'b01010000011: data <= 32'h3ab6b964;
    11'b01010000100: data <= 32'h392ebb03;
    11'b01010000101: data <= 32'h3d29349a;
    11'b01010000110: data <= 32'h3cd43e4e;
    11'b01010000111: data <= 32'ha48c3b86;
    11'b01010001000: data <= 32'hbc13bd4c;
    11'b01010001001: data <= 32'hbb42c14a;
    11'b01010001010: data <= 32'hb75cbece;
    11'b01010001011: data <= 32'hb743b12e;
    11'b01010001100: data <= 32'hb50fa7ec;
    11'b01010001101: data <= 32'h3783b9f6;
    11'b01010001110: data <= 32'h3ab7b660;
    11'b01010001111: data <= 32'hb6533c65;
    11'b01010010000: data <= 32'hc0713fad;
    11'b01010010001: data <= 32'hc0bc3cb2;
    11'b01010010010: data <= 32'hb8722c42;
    11'b01010010011: data <= 32'h3bbdb268;
    11'b01010010100: data <= 32'h3957a7df;
    11'b01010010101: data <= 32'hb060afde;
    11'b01010010110: data <= 32'h377b2a22;
    11'b01010010111: data <= 32'h3faf3c50;
    11'b01010011000: data <= 32'h40223fb7;
    11'b01010011001: data <= 32'h37d13c52;
    11'b01010011010: data <= 32'hbb56bb60;
    11'b01010011011: data <= 32'hba2cbf73;
    11'b01010011100: data <= 32'h2ec5bc11;
    11'b01010011101: data <= 32'h3754b2d2;
    11'b01010011110: data <= 32'h3778bb86;
    11'b01010011111: data <= 32'h3a12bfd8;
    11'b01010100000: data <= 32'h3a13bce6;
    11'b01010100001: data <= 32'hb63f3ac3;
    11'b01010100010: data <= 32'hbf933f52;
    11'b01010100011: data <= 32'hc0113a2b;
    11'b01010100100: data <= 32'hba77b952;
    11'b01010100101: data <= 32'hae09ba8a;
    11'b01010100110: data <= 32'hb9ecb006;
    11'b01010100111: data <= 32'hbc9033d9;
    11'b01010101000: data <= 32'h32663708;
    11'b01010101001: data <= 32'h40163caf;
    11'b01010101010: data <= 32'h40023f9b;
    11'b01010101011: data <= 32'h2d0e3dcb;
    11'b01010101100: data <= 32'hbd253007;
    11'b01010101101: data <= 32'hb91db7a6;
    11'b01010101110: data <= 32'h3a03a69e;
    11'b01010101111: data <= 32'h3cb7ab6d;
    11'b01010110000: data <= 32'h3ae4bd7e;
    11'b01010110001: data <= 32'h3b30c0b1;
    11'b01010110010: data <= 32'h3c69bce7;
    11'b01010110011: data <= 32'h37b13ba2;
    11'b01010110100: data <= 32'hb9d63e2a;
    11'b01010110101: data <= 32'hbcf3a8e7;
    11'b01010110110: data <= 32'hbaefbe57;
    11'b01010110111: data <= 32'hbadbbd72;
    11'b01010111000: data <= 32'hbe45b427;
    11'b01010111001: data <= 32'hbe2f2e02;
    11'b01010111010: data <= 32'h2e1daf3e;
    11'b01010111011: data <= 32'h3eec359d;
    11'b01010111100: data <= 32'h3ce63d9a;
    11'b01010111101: data <= 32'hbad23f0f;
    11'b01010111110: data <= 32'hbf503cae;
    11'b01010111111: data <= 32'hb90b3970;
    11'b01011000000: data <= 32'h3b66395b;
    11'b01011000001: data <= 32'h3c2f30e3;
    11'b01011000010: data <= 32'h36d8bcba;
    11'b01011000011: data <= 32'h397ebf32;
    11'b01011000100: data <= 32'h3e80b7ca;
    11'b01011000101: data <= 32'h3ecc3d6e;
    11'b01011000110: data <= 32'h38bd3d4f;
    11'b01011000111: data <= 32'hb6fdb891;
    11'b01011001000: data <= 32'hb9a5bf94;
    11'b01011001001: data <= 32'hbb57bd2b;
    11'b01011001010: data <= 32'hbd94b3b6;
    11'b01011001011: data <= 32'hbc9ab7cb;
    11'b01011001100: data <= 32'h3441bd5d;
    11'b01011001101: data <= 32'h3d47bbaf;
    11'b01011001110: data <= 32'h36963966;
    11'b01011001111: data <= 32'hbe123f3b;
    11'b01011010000: data <= 32'hc0123e55;
    11'b01011010001: data <= 32'hb9673b86;
    11'b01011010010: data <= 32'h37923949;
    11'b01011010011: data <= 32'h20ee3355;
    11'b01011010100: data <= 32'hb9aeb91d;
    11'b01011010101: data <= 32'h30f1badd;
    11'b01011010110: data <= 32'h3fd535ab;
    11'b01011010111: data <= 32'h41043ec8;
    11'b01011011000: data <= 32'h3d153d3a;
    11'b01011011001: data <= 32'hafd3b676;
    11'b01011011010: data <= 32'hb78bbce7;
    11'b01011011011: data <= 32'hb5d2b75d;
    11'b01011011100: data <= 32'hb8032ae3;
    11'b01011011101: data <= 32'hb57abc5a;
    11'b01011011110: data <= 32'h386fc0fc;
    11'b01011011111: data <= 32'h3c7dbfe6;
    11'b01011100000: data <= 32'h32e93142;
    11'b01011100001: data <= 32'hbd363e50;
    11'b01011100010: data <= 32'hbe4d3cc1;
    11'b01011100011: data <= 32'hb8cc342c;
    11'b01011100100: data <= 32'hb4742aa3;
    11'b01011100101: data <= 32'hbd503033;
    11'b01011100110: data <= 32'hbfa8b221;
    11'b01011100111: data <= 32'hb68db4d2;
    11'b01011101000: data <= 32'h3f993877;
    11'b01011101001: data <= 32'h40e43e47;
    11'b01011101010: data <= 32'h3b903d80;
    11'b01011101011: data <= 32'hb7153576;
    11'b01011101100: data <= 32'hb5512d4c;
    11'b01011101101: data <= 32'h354f39ea;
    11'b01011101110: data <= 32'h3590384b;
    11'b01011101111: data <= 32'h3117bd37;
    11'b01011110000: data <= 32'h3907c1be;
    11'b01011110001: data <= 32'h3cd0c02f;
    11'b01011110010: data <= 32'h3a6331b4;
    11'b01011110011: data <= 32'hb30b3d0d;
    11'b01011110100: data <= 32'hb8913595;
    11'b01011110101: data <= 32'hb4f3ba04;
    11'b01011110110: data <= 32'hba5fb8b5;
    11'b01011110111: data <= 32'hc0492863;
    11'b01011111000: data <= 32'hc0f0afda;
    11'b01011111001: data <= 32'hb944b8af;
    11'b01011111010: data <= 32'h3e20b17e;
    11'b01011111011: data <= 32'h3e983afd;
    11'b01011111100: data <= 32'ha9ce3d56;
    11'b01011111101: data <= 32'hbc413c7a;
    11'b01011111110: data <= 32'hb4ed3ce6;
    11'b01011111111: data <= 32'h39793e76;
    11'b01100000000: data <= 32'h37593b8c;
    11'b01100000001: data <= 32'hb193bc18;
    11'b01100000010: data <= 32'h33d3c0a1;
    11'b01100000011: data <= 32'h3d80bd50;
    11'b01100000100: data <= 32'h3ef43917;
    11'b01100000101: data <= 32'h3c533c2d;
    11'b01100000110: data <= 32'h3704b53a;
    11'b01100000111: data <= 32'h2e4fbd1f;
    11'b01100001000: data <= 32'hb9dcb906;
    11'b01100001001: data <= 32'hbfe0323c;
    11'b01100001010: data <= 32'hc02db5f8;
    11'b01100001011: data <= 32'hb776be1f;
    11'b01100001100: data <= 32'h3c78bdd2;
    11'b01100001101: data <= 32'h39c4ad0b;
    11'b01100001110: data <= 32'hbb3f3c59;
    11'b01100001111: data <= 32'hbd8c3d7f;
    11'b01100010000: data <= 32'hb3c23df7;
    11'b01100010001: data <= 32'h38483eab;
    11'b01100010010: data <= 32'hb4c23c2a;
    11'b01100010011: data <= 32'hbd19b786;
    11'b01100010100: data <= 32'hb82abd23;
    11'b01100010101: data <= 32'h3d8cb515;
    11'b01100010110: data <= 32'h40b73c5f;
    11'b01100010111: data <= 32'h3f153b8e;
    11'b01100011000: data <= 32'h3ae1b6ea;
    11'b01100011001: data <= 32'h3682bb16;
    11'b01100011010: data <= 32'hb0d230ef;
    11'b01100011011: data <= 32'hbc0a39bd;
    11'b01100011100: data <= 32'hbc90b915;
    11'b01100011101: data <= 32'habd3c0f0;
    11'b01100011110: data <= 32'h3af2c0f8;
    11'b01100011111: data <= 32'h348bb9eb;
    11'b01100100000: data <= 32'hbba739d3;
    11'b01100100001: data <= 32'hbbf03b66;
    11'b01100100010: data <= 32'h29ef3a20;
    11'b01100100011: data <= 32'h300d3ba7;
    11'b01100100100: data <= 32'hbda13aba;
    11'b01100100101: data <= 32'hc0fe1f6e;
    11'b01100100110: data <= 32'hbd17b824;
    11'b01100100111: data <= 32'h3c9430a1;
    11'b01100101000: data <= 32'h406c3c36;
    11'b01100101001: data <= 32'h3dac3a95;
    11'b01100101010: data <= 32'h37b6a693;
    11'b01100101011: data <= 32'h378631e8;
    11'b01100101100: data <= 32'h38823d7c;
    11'b01100101101: data <= 32'h25273dac;
    11'b01100101110: data <= 32'hb646b8fa;
    11'b01100101111: data <= 32'h2f9dc17a;
    11'b01100110000: data <= 32'h3a53c12e;
    11'b01100110001: data <= 32'h3850b9bd;
    11'b01100110010: data <= 32'hafd2372c;
    11'b01100110011: data <= 32'h265b2c4f;
    11'b01100110100: data <= 32'h3898b667;
    11'b01100110101: data <= 32'hafed2d83;
    11'b01100110110: data <= 32'hc02e38f9;
    11'b01100110111: data <= 32'hc21e3273;
    11'b01100111000: data <= 32'hbe42b7e0;
    11'b01100111001: data <= 32'h3a22b53f;
    11'b01100111010: data <= 32'h3d8c35bf;
    11'b01100111011: data <= 32'h34c8384a;
    11'b01100111100: data <= 32'hb583374d;
    11'b01100111101: data <= 32'h35dd3cb4;
    11'b01100111110: data <= 32'h3c0b408d;
    11'b01100111111: data <= 32'h36b53fae;
    11'b01101000000: data <= 32'hb75db483;
    11'b01101000001: data <= 32'hb3b4c048;
    11'b01101000010: data <= 32'h39c7bee6;
    11'b01101000011: data <= 32'h3ca7ad68;
    11'b01101000100: data <= 32'h3c0b35a4;
    11'b01101000101: data <= 32'h3c50b972;
    11'b01101000110: data <= 32'h3c83bcc7;
    11'b01101000111: data <= 32'h2a7cb324;
    11'b01101001000: data <= 32'hbf7239da;
    11'b01101001001: data <= 32'hc1353189;
    11'b01101001010: data <= 32'hbcf3bc74;
    11'b01101001011: data <= 32'h3758bdb3;
    11'b01101001100: data <= 32'h366fb929;
    11'b01101001101: data <= 32'hba732e6c;
    11'b01101001110: data <= 32'hbb843867;
    11'b01101001111: data <= 32'h35b03d7e;
    11'b01101010000: data <= 32'h3c3c4091;
    11'b01101010001: data <= 32'ha2e93fba;
    11'b01101010010: data <= 32'hbd6e321f;
    11'b01101010011: data <= 32'hbc38bc3e;
    11'b01101010100: data <= 32'h381eb7d4;
    11'b01101010101: data <= 32'h3e513920;
    11'b01101010110: data <= 32'h3e77359e;
    11'b01101010111: data <= 32'h3df4bba9;
    11'b01101011000: data <= 32'h3d9fbc79;
    11'b01101011001: data <= 32'h38b4356f;
    11'b01101011010: data <= 32'hbada3d2b;
    11'b01101011011: data <= 32'hbdd230b3;
    11'b01101011100: data <= 32'hb896bf42;
    11'b01101011101: data <= 32'h3533c0b6;
    11'b01101011110: data <= 32'hb1d7bd4d;
    11'b01101011111: data <= 32'hbcaeb49d;
    11'b01101100000: data <= 32'hba412e87;
    11'b01101100001: data <= 32'h394f38d1;
    11'b01101100010: data <= 32'h3b213d9b;
    11'b01101100011: data <= 32'hbae33df9;
    11'b01101100100: data <= 32'hc0ef385e;
    11'b01101100101: data <= 32'hbf68b160;
    11'b01101100110: data <= 32'h31f7347f;
    11'b01101100111: data <= 32'h3d8c3ada;
    11'b01101101000: data <= 32'h3cdc3386;
    11'b01101101001: data <= 32'h3bceba4c;
    11'b01101101010: data <= 32'h3d11b541;
    11'b01101101011: data <= 32'h3cbc3db9;
    11'b01101101100: data <= 32'h3480401c;
    11'b01101101101: data <= 32'hb68534b6;
    11'b01101101110: data <= 32'hafa0bff8;
    11'b01101101111: data <= 32'h3480c0d2;
    11'b01101110000: data <= 32'hb0e2bcd3;
    11'b01101110001: data <= 32'hb90db69a;
    11'b01101110010: data <= 32'h2de2b93c;
    11'b01101110011: data <= 32'h3d0db942;
    11'b01101110100: data <= 32'h3a8233e7;
    11'b01101110101: data <= 32'hbda83be9;
    11'b01101110110: data <= 32'hc1f2396b;
    11'b01101110111: data <= 32'hc02c2c49;
    11'b01101111000: data <= 32'hadbd2f77;
    11'b01101111001: data <= 32'h39163546;
    11'b01101111010: data <= 32'h2202afcb;
    11'b01101111011: data <= 32'haf5eb80f;
    11'b01101111100: data <= 32'h3b0537fe;
    11'b01101111101: data <= 32'h3e2d408e;
    11'b01101111110: data <= 32'h3af94115;
    11'b01101111111: data <= 32'hb10438b5;
    11'b01110000000: data <= 32'hb488bdbd;
    11'b01110000001: data <= 32'h30ffbddd;
    11'b01110000010: data <= 32'h3402b561;
    11'b01110000011: data <= 32'h34ecb380;
    11'b01110000100: data <= 32'h3c55bd36;
    11'b01110000101: data <= 32'h3f5bbe81;
    11'b01110000110: data <= 32'h3bfdb635;
    11'b01110000111: data <= 32'hbcc43afc;
    11'b01110001000: data <= 32'hc0e53975;
    11'b01110001001: data <= 32'hbe38b530;
    11'b01110001010: data <= 32'hb0b8ba11;
    11'b01110001011: data <= 32'hb3ebb8d3;
    11'b01110001100: data <= 32'hbd04b8e4;
    11'b01110001101: data <= 32'hbc27b7a4;
    11'b01110001110: data <= 32'h38e9395b;
    11'b01110001111: data <= 32'h3e654074;
    11'b01110010000: data <= 32'h395940c7;
    11'b01110010001: data <= 32'hba733ac6;
    11'b01110010010: data <= 32'hbc08b735;
    11'b01110010011: data <= 32'haff6ad28;
    11'b01110010100: data <= 32'h387039ba;
    11'b01110010101: data <= 32'h3ad228d1;
    11'b01110010110: data <= 32'h3dcabe3c;
    11'b01110010111: data <= 32'h4000bf19;
    11'b01110011000: data <= 32'h3d76ae2a;
    11'b01110011001: data <= 32'hb44d3d46;
    11'b01110011010: data <= 32'hbca639e1;
    11'b01110011011: data <= 32'hb894bb04;
    11'b01110011100: data <= 32'h1d00be63;
    11'b01110011101: data <= 32'hba51bcfd;
    11'b01110011110: data <= 32'hbf5bbb7b;
    11'b01110011111: data <= 32'hbcb2ba77;
    11'b01110100000: data <= 32'h3a39a8c6;
    11'b01110100001: data <= 32'h3e043ce3;
    11'b01110100010: data <= 32'h9c273e9a;
    11'b01110100011: data <= 32'hbf2b3b4d;
    11'b01110100100: data <= 32'hbf163624;
    11'b01110100101: data <= 32'hb6f13b40;
    11'b01110100110: data <= 32'h36cd3cfe;
    11'b01110100111: data <= 32'h37e22e4b;
    11'b01110101000: data <= 32'h3aa7bdcc;
    11'b01110101001: data <= 32'h3e5fbcb6;
    11'b01110101010: data <= 32'h3ebb3abf;
    11'b01110101011: data <= 32'h3a664018;
    11'b01110101100: data <= 32'h2e3e3b36;
    11'b01110101101: data <= 32'h3305bc42;
    11'b01110101110: data <= 32'h3183beab;
    11'b01110101111: data <= 32'hba6cbc2e;
    11'b01110110000: data <= 32'hbe08baa7;
    11'b01110110001: data <= 32'hb7b5bd3f;
    11'b01110110010: data <= 32'h3d55bce5;
    11'b01110110011: data <= 32'h3de4b05e;
    11'b01110110100: data <= 32'hb82e3a5b;
    11'b01110110101: data <= 32'hc0963a67;
    11'b01110110110: data <= 32'hbfc83921;
    11'b01110110111: data <= 32'hb83e3bb5;
    11'b01110111000: data <= 32'haf063b7c;
    11'b01110111001: data <= 32'hb922b248;
    11'b01110111010: data <= 32'hb735bcef;
    11'b01110111011: data <= 32'h3acdb6c9;
    11'b01110111100: data <= 32'h3f1b3ea5;
    11'b01110111101: data <= 32'h3d9140fb;
    11'b01110111110: data <= 32'h38a43c43;
    11'b01110111111: data <= 32'h34e6b974;
    11'b01111000000: data <= 32'h3066ba43;
    11'b01111000001: data <= 32'hb78f81cc;
    11'b01111000010: data <= 32'hb96bb4fa;
    11'b01111000011: data <= 32'h375abeb9;
    11'b01111000100: data <= 32'h3f8ac05b;
    11'b01111000101: data <= 32'h3e4fbc0b;
    11'b01111000110: data <= 32'hb6e03641;
    11'b01111000111: data <= 32'hbf45396f;
    11'b01111001000: data <= 32'hbd093524;
    11'b01111001001: data <= 32'hb44b3348;
    11'b01111001010: data <= 32'hb9bb2d24;
    11'b01111001011: data <= 32'hbf87b961;
    11'b01111001100: data <= 32'hbe78bcac;
    11'b01111001101: data <= 32'h3445b159;
    11'b01111001110: data <= 32'h3eaa3e9c;
    11'b01111001111: data <= 32'h3d00406c;
    11'b01111010000: data <= 32'h2e433c25;
    11'b01111010001: data <= 32'hb4ec28fd;
    11'b01111010010: data <= 32'hb0223895;
    11'b01111010011: data <= 32'hb1763d31;
    11'b01111010100: data <= 32'had9e34e2;
    11'b01111010101: data <= 32'h3adbbef4;
    11'b01111010110: data <= 32'h3fcec0c0;
    11'b01111010111: data <= 32'h3ecbbb49;
    11'b01111011000: data <= 32'h3401397f;
    11'b01111011001: data <= 32'hb88139a3;
    11'b01111011010: data <= 32'ha84cb272;
    11'b01111011011: data <= 32'h33ceb8ea;
    11'b01111011100: data <= 32'hbc22b8b0;
    11'b01111011101: data <= 32'hc103bb75;
    11'b01111011110: data <= 32'hbfdfbd35;
    11'b01111011111: data <= 32'h33a9b945;
    11'b01111100000: data <= 32'h3e153978;
    11'b01111100001: data <= 32'h38fe3cf7;
    11'b01111100010: data <= 32'hbad739e8;
    11'b01111100011: data <= 32'hbc4f3909;
    11'b01111100100: data <= 32'hb6703e5d;
    11'b01111100101: data <= 32'hb0f14022;
    11'b01111100110: data <= 32'hb43f38ce;
    11'b01111100111: data <= 32'h347fbe31;
    11'b01111101000: data <= 32'h3d56bf55;
    11'b01111101001: data <= 32'h3ea5a8f3;
    11'b01111101010: data <= 32'h3c423d98;
    11'b01111101011: data <= 32'h39c53ad3;
    11'b01111101100: data <= 32'h3c11b7d1;
    11'b01111101101: data <= 32'h3982baa8;
    11'b01111101110: data <= 32'hbb77b6db;
    11'b01111101111: data <= 32'hc077b936;
    11'b01111110000: data <= 32'hbd81bde6;
    11'b01111110001: data <= 32'h3a02be5d;
    11'b01111110010: data <= 32'h3deab98c;
    11'b01111110011: data <= 32'h29c82f22;
    11'b01111110100: data <= 32'hbde034f6;
    11'b01111110101: data <= 32'hbd3139ef;
    11'b01111110110: data <= 32'hb5b73ed6;
    11'b01111110111: data <= 32'hb64b3f92;
    11'b01111111000: data <= 32'hbc9e3629;
    11'b01111111001: data <= 32'hbc0cbd48;
    11'b01111111010: data <= 32'h34febc33;
    11'b01111111011: data <= 32'h3da23ae3;
    11'b01111111100: data <= 32'h3ded3f8f;
    11'b01111111101: data <= 32'h3d123b4a;
    11'b01111111110: data <= 32'h3d1fb5c1;
    11'b01111111111: data <= 32'h3a36b1a4;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    