module top_combine(
CLK, rst,
CEB, ssb, sdi,
vmm_load,
output_z_0, output_z_1, output_z_2, output_z_3
);

input  CLK, rst;
input  CEB;
output [31:0] output_z_0, output_z_1, output_z_2, output_z_3;


wire [31:0] output_data_divider1, output_data_divider2, output_data_divider3, output_data_divider4;
wire [31:0] output_data_divider5, output_data_divider6, output_data_divider7, output_data_divider8;
wire [31:0] output_data_divider9, output_data_divider10, output_data_divider11, output_data_divider12;
wire [31:0] output_data_divider13, output_data_divider14, output_data_divider15, output_data_divider16;
wire [31:0] output_data_divider17, output_data_divider18, output_data_divider19, output_data_divider20;
wire [31:0] output_data_divider21, output_data_divider22, output_data_divider23, output_data_divider24;
wire [31:0] output_data_divider25, output_data_divider26, output_data_divider27, output_data_divider28;
wire [31:0] output_data_divider29, output_data_divider30, output_data_divider31, output_data_divider32;
wire [31:0] output_data_divider33, output_data_divider34, output_data_divider35, output_data_divider36;
wire [31:0] output_data_divider37, output_data_divider38, output_data_divider39, output_data_divider40;
wire [31:0] output_data_divider41, output_data_divider42, output_data_divider43, output_data_divider44;
wire [31:0] output_data_divider45, output_data_divider46, output_data_divider47, output_data_divider48;
wire [31:0] output_data_divider49, output_data_divider50, output_data_divider51, output_data_divider52;
wire [31:0] output_data_divider53, output_data_divider54, output_data_divider55, output_data_divider56;
wire [31:0] output_data_divider57, output_data_divider58, output_data_divider59, output_data_divider60;
wire [31:0] output_data_divider61, output_data_divider62, output_data_divider63, output_data_divider64;

StreamData DUT_DATA_Data(
.CLK(CLK),               
.rst(rst),               
.CEB(CEB),  
.output1(output_data_divider1), .output2(output_data_divider2), .output3(output_data_divider3), .output4(output_data_divider4),
.output5(output_data_divider5), .output6(output_data_divider6), .output7(output_data_divider7), .output8(output_data_divider8),
.output9(output_data_divider9), .output10(output_data_divider10), .output11(output_data_divider11), .output12(output_data_divider12),
.output13(output_data_divider13), .output14(output_data_divider14), .output15(output_data_divider15), .output16(output_data_divider16),
.output17(output_data_divider17), .output18(output_data_divider18), .output19(output_data_divider19), .output20(output_data_divider20),
.output21(output_data_divider21), .output22(output_data_divider22), .output23(output_data_divider23), .output24(output_data_divider24),
.output25(output_data_divider25), .output26(output_data_divider26), .output27(output_data_divider27), .output28(output_data_divider28),
.output29(output_data_divider29), .output30(output_data_divider30), .output31(output_data_divider31), .output32(output_data_divider32),
.output33(output_data_divider33), .output34(output_data_divider34), .output35(output_data_divider35), .output36(output_data_divider36),
.output37(output_data_divider37), .output38(output_data_divider38), .output39(output_data_divider39), .output40(output_data_divider40),
.output41(output_data_divider41), .output42(output_data_divider42), .output43(output_data_divider43), .output44(output_data_divider44),
.output45(output_data_divider45), .output46(output_data_divider46), .output47(output_data_divider47), .output48(output_data_divider48),
.output49(output_data_divider49), .output50(output_data_divider50), .output51(output_data_divider51), .output52(output_data_divider52),
.output53(output_data_divider53), .output54(output_data_divider54), .output55(output_data_divider55), .output56(output_data_divider56),
.output57(output_data_divider57), .output58(output_data_divider58), .output59(output_data_divider59), .output60(output_data_divider60),
.output61(output_data_divider61), .output62(output_data_divider62), .output63(output_data_divider63), .output64(output_data_divider64) 
);

wire [15:0] output_z_real1_0;
wire [15:0] output_z_imag1_0;
wire [15:0] output_z_real1_1;
wire [15:0] output_z_imag1_1;
wire [15:0] output_z_real1_2;
wire [15:0] output_z_imag1_2;
wire [15:0] output_z_real1_3;
wire [15:0] output_z_imag1_3;

input ssb;
input [27:0] sdi;
input vmm_load;
wire [9:0] output_real_1_0, output_real_1_1, output_real_1_2, output_real_1_3;
wire [9:0] output_imag_1_0, output_imag_1_1, output_imag_1_2, output_imag_1_3;
wire [9:0] output_real_2_0, output_real_2_1, output_real_2_2, output_real_2_3;
wire [9:0] output_imag_2_0, output_imag_2_1, output_imag_2_2, output_imag_2_3;
wire [9:0] output_real_3_0, output_real_3_1, output_real_3_2, output_real_3_3;
wire [9:0] output_imag_3_0, output_imag_3_1, output_imag_3_2, output_imag_3_3;
wire [9:0] output_real_4_0, output_real_4_1, output_real_4_2, output_real_4_3;
wire [9:0] output_imag_4_0, output_imag_4_1, output_imag_4_2, output_imag_4_3;
wire [9:0] output_real_5_0, output_real_5_1, output_real_5_2, output_real_5_3;
wire [9:0] output_imag_5_0, output_imag_5_1, output_imag_5_2, output_imag_5_3;
wire [9:0] output_real_6_0, output_real_6_1, output_real_6_2, output_real_6_3;
wire [9:0] output_imag_6_0, output_imag_6_1, output_imag_6_2, output_imag_6_3;
wire [9:0] output_real_7_0, output_real_7_1, output_real_7_2, output_real_7_3;
wire [9:0] output_imag_7_0, output_imag_7_1, output_imag_7_2, output_imag_7_3;
wire [9:0] output_real_8_0, output_real_8_1, output_real_8_2, output_real_8_3;
wire [9:0] output_imag_8_0, output_imag_8_1, output_imag_8_2, output_imag_8_3;
wire [9:0] output_real_9_0, output_real_9_1, output_real_9_2, output_real_9_3;
wire [9:0] output_imag_9_0, output_imag_9_1, output_imag_9_2, output_imag_9_3;
wire [9:0] output_real_10_0, output_real_10_1, output_real_10_2, output_real_10_3;
wire [9:0] output_imag_10_0, output_imag_10_1, output_imag_10_2, output_imag_10_3;
wire [9:0] output_real_11_0, output_real_11_1, output_real_11_2, output_real_11_3;
wire [9:0] output_imag_11_0, output_imag_11_1, output_imag_11_2, output_imag_11_3;
wire [9:0] output_real_12_0, output_real_12_1, output_real_12_2, output_real_12_3;
wire [9:0] output_imag_12_0, output_imag_12_1, output_imag_12_2, output_imag_12_3;
wire [9:0] output_real_13_0, output_real_13_1, output_real_13_2, output_real_13_3;
wire [9:0] output_imag_13_0, output_imag_13_1, output_imag_13_2, output_imag_13_3;
wire [9:0] output_real_14_0, output_real_14_1, output_real_14_2, output_real_14_3;
wire [9:0] output_imag_14_0, output_imag_14_1, output_imag_14_2, output_imag_14_3;
wire [9:0] output_real_15_0, output_real_15_1, output_real_15_2, output_real_15_3;
wire [9:0] output_imag_15_0, output_imag_15_1, output_imag_15_2, output_imag_15_3;
wire [9:0] output_real_16_0, output_real_16_1, output_real_16_2, output_real_16_3;
wire [9:0] output_imag_16_0, output_imag_16_1, output_imag_16_2, output_imag_16_3;
wire [9:0] output_real_17_0, output_real_17_1, output_real_17_2, output_real_17_3;
wire [9:0] output_imag_17_0, output_imag_17_1, output_imag_17_2, output_imag_17_3;
wire [9:0] output_real_18_0, output_real_18_1, output_real_18_2, output_real_18_3;
wire [9:0] output_imag_18_0, output_imag_18_1, output_imag_18_2, output_imag_18_3;
wire [9:0] output_real_19_0, output_real_19_1, output_real_19_2, output_real_19_3;
wire [9:0] output_imag_19_0, output_imag_19_1, output_imag_19_2, output_imag_19_3;
wire [9:0] output_real_20_0, output_real_20_1, output_real_20_2, output_real_20_3;
wire [9:0] output_imag_20_0, output_imag_20_1, output_imag_20_2, output_imag_20_3;
wire [9:0] output_real_21_0, output_real_21_1, output_real_21_2, output_real_21_3;
wire [9:0] output_imag_21_0, output_imag_21_1, output_imag_21_2, output_imag_21_3;
wire [9:0] output_real_22_0, output_real_22_1, output_real_22_2, output_real_22_3;
wire [9:0] output_imag_22_0, output_imag_22_1, output_imag_22_2, output_imag_22_3;
wire [9:0] output_real_23_0, output_real_23_1, output_real_23_2, output_real_23_3;
wire [9:0] output_imag_23_0, output_imag_23_1, output_imag_23_2, output_imag_23_3;
wire [9:0] output_real_24_0, output_real_24_1, output_real_24_2, output_real_24_3;
wire [9:0] output_imag_24_0, output_imag_24_1, output_imag_24_2, output_imag_24_3;
wire [9:0] output_real_25_0, output_real_25_1, output_real_25_2, output_real_25_3;
wire [9:0] output_imag_25_0, output_imag_25_1, output_imag_25_2, output_imag_25_3;
wire [9:0] output_real_26_0, output_real_26_1, output_real_26_2, output_real_26_3;
wire [9:0] output_imag_26_0, output_imag_26_1, output_imag_26_2, output_imag_26_3;
wire [9:0] output_real_27_0, output_real_27_1, output_real_27_2, output_real_27_3;
wire [9:0] output_imag_27_0, output_imag_27_1, output_imag_27_2, output_imag_27_3;
wire [9:0] output_real_28_0, output_real_28_1, output_real_28_2, output_real_28_3;
wire [9:0] output_imag_28_0, output_imag_28_1, output_imag_28_2, output_imag_28_3;
wire [9:0] output_real_29_0, output_real_29_1, output_real_29_2, output_real_29_3;
wire [9:0] output_imag_29_0, output_imag_29_1, output_imag_29_2, output_imag_29_3;
wire [9:0] output_real_30_0, output_real_30_1, output_real_30_2, output_real_30_3;
wire [9:0] output_imag_30_0, output_imag_30_1, output_imag_30_2, output_imag_30_3;
wire [9:0] output_real_31_0, output_real_31_1, output_real_31_2, output_real_31_3;
wire [9:0] output_imag_31_0, output_imag_31_1, output_imag_31_2, output_imag_31_3;
wire [9:0] output_real_32_0, output_real_32_1, output_real_32_2, output_real_32_3;
wire [9:0] output_imag_32_0, output_imag_32_1, output_imag_32_2, output_imag_32_3;
wire [9:0] output_real_33_0, output_real_33_1, output_real_33_2, output_real_33_3;
wire [9:0] output_imag_33_0, output_imag_33_1, output_imag_33_2, output_imag_33_3;
wire [9:0] output_real_34_0, output_real_34_1, output_real_34_2, output_real_34_3;
wire [9:0] output_imag_34_0, output_imag_34_1, output_imag_34_2, output_imag_34_3;
wire [9:0] output_real_35_0, output_real_35_1, output_real_35_2, output_real_35_3;
wire [9:0] output_imag_35_0, output_imag_35_1, output_imag_35_2, output_imag_35_3;
wire [9:0] output_real_36_0, output_real_36_1, output_real_36_2, output_real_36_3;
wire [9:0] output_imag_36_0, output_imag_36_1, output_imag_36_2, output_imag_36_3;
wire [9:0] output_real_37_0, output_real_37_1, output_real_37_2, output_real_37_3;
wire [9:0] output_imag_37_0, output_imag_37_1, output_imag_37_2, output_imag_37_3;
wire [9:0] output_real_38_0, output_real_38_1, output_real_38_2, output_real_38_3;
wire [9:0] output_imag_38_0, output_imag_38_1, output_imag_38_2, output_imag_38_3;
wire [9:0] output_real_39_0, output_real_39_1, output_real_39_2, output_real_39_3;
wire [9:0] output_imag_39_0, output_imag_39_1, output_imag_39_2, output_imag_39_3;
wire [9:0] output_real_40_0, output_real_40_1, output_real_40_2, output_real_40_3;
wire [9:0] output_imag_40_0, output_imag_40_1, output_imag_40_2, output_imag_40_3;
wire [9:0] output_real_41_0, output_real_41_1, output_real_41_2, output_real_41_3;
wire [9:0] output_imag_41_0, output_imag_41_1, output_imag_41_2, output_imag_41_3;
wire [9:0] output_real_42_0, output_real_42_1, output_real_42_2, output_real_42_3;
wire [9:0] output_imag_42_0, output_imag_42_1, output_imag_42_2, output_imag_42_3;
wire [9:0] output_real_43_0, output_real_43_1, output_real_43_2, output_real_43_3;
wire [9:0] output_imag_43_0, output_imag_43_1, output_imag_43_2, output_imag_43_3;
wire [9:0] output_real_44_0, output_real_44_1, output_real_44_2, output_real_44_3;
wire [9:0] output_imag_44_0, output_imag_44_1, output_imag_44_2, output_imag_44_3;
wire [9:0] output_real_45_0, output_real_45_1, output_real_45_2, output_real_45_3;
wire [9:0] output_imag_45_0, output_imag_45_1, output_imag_45_2, output_imag_45_3;
wire [9:0] output_real_46_0, output_real_46_1, output_real_46_2, output_real_46_3;
wire [9:0] output_imag_46_0, output_imag_46_1, output_imag_46_2, output_imag_46_3;
wire [9:0] output_real_47_0, output_real_47_1, output_real_47_2, output_real_47_3;
wire [9:0] output_imag_47_0, output_imag_47_1, output_imag_47_2, output_imag_47_3;
wire [9:0] output_real_48_0, output_real_48_1, output_real_48_2, output_real_48_3;
wire [9:0] output_imag_48_0, output_imag_48_1, output_imag_48_2, output_imag_48_3;
wire [9:0] output_real_49_0, output_real_49_1, output_real_49_2, output_real_49_3;
wire [9:0] output_imag_49_0, output_imag_49_1, output_imag_49_2, output_imag_49_3;
wire [9:0] output_real_50_0, output_real_50_1, output_real_50_2, output_real_50_3;
wire [9:0] output_imag_50_0, output_imag_50_1, output_imag_50_2, output_imag_50_3;
wire [9:0] output_real_51_0, output_real_51_1, output_real_51_2, output_real_51_3;
wire [9:0] output_imag_51_0, output_imag_51_1, output_imag_51_2, output_imag_51_3;
wire [9:0] output_real_52_0, output_real_52_1, output_real_52_2, output_real_52_3;
wire [9:0] output_imag_52_0, output_imag_52_1, output_imag_52_2, output_imag_52_3;
wire [9:0] output_real_53_0, output_real_53_1, output_real_53_2, output_real_53_3;
wire [9:0] output_imag_53_0, output_imag_53_1, output_imag_53_2, output_imag_53_3;
wire [9:0] output_real_54_0, output_real_54_1, output_real_54_2, output_real_54_3;
wire [9:0] output_imag_54_0, output_imag_54_1, output_imag_54_2, output_imag_54_3;
wire [9:0] output_real_55_0, output_real_55_1, output_real_55_2, output_real_55_3;
wire [9:0] output_imag_55_0, output_imag_55_1, output_imag_55_2, output_imag_55_3;
wire [9:0] output_real_56_0, output_real_56_1, output_real_56_2, output_real_56_3;
wire [9:0] output_imag_56_0, output_imag_56_1, output_imag_56_2, output_imag_56_3;
wire [9:0] output_real_57_0, output_real_57_1, output_real_57_2, output_real_57_3;
wire [9:0] output_imag_57_0, output_imag_57_1, output_imag_57_2, output_imag_57_3;
wire [9:0] output_real_58_0, output_real_58_1, output_real_58_2, output_real_58_3;
wire [9:0] output_imag_58_0, output_imag_58_1, output_imag_58_2, output_imag_58_3;
wire [9:0] output_real_59_0, output_real_59_1, output_real_59_2, output_real_59_3;
wire [9:0] output_imag_59_0, output_imag_59_1, output_imag_59_2, output_imag_59_3;
wire [9:0] output_real_60_0, output_real_60_1, output_real_60_2, output_real_60_3;
wire [9:0] output_imag_60_0, output_imag_60_1, output_imag_60_2, output_imag_60_3;
wire [9:0] output_real_61_0, output_real_61_1, output_real_61_2, output_real_61_3;
wire [9:0] output_imag_61_0, output_imag_61_1, output_imag_61_2, output_imag_61_3;
wire [9:0] output_real_62_0, output_real_62_1, output_real_62_2, output_real_62_3;
wire [9:0] output_imag_62_0, output_imag_62_1, output_imag_62_2, output_imag_62_3;
wire [9:0] output_real_63_0, output_real_63_1, output_real_63_2, output_real_63_3;
wire [9:0] output_imag_63_0, output_imag_63_1, output_imag_63_2, output_imag_63_3;
wire [9:0] output_real_64_0, output_real_64_1, output_real_64_2, output_real_64_3;
wire [9:0] output_imag_64_0, output_imag_64_1, output_imag_64_2, output_imag_64_3;

pin_update_vmm_input DUT_VMM_INPUT(
.output_real_0_0(output_real_1_0), .output_imag_0_0(output_imag_1_0),
.output_real_1_0(output_real_2_0), .output_imag_1_0(output_imag_2_0),
.output_real_2_0(output_real_3_0), .output_imag_2_0(output_imag_3_0),
.output_real_3_0(output_real_4_0), .output_imag_3_0(output_imag_4_0),
.output_real_4_0(output_real_5_0), .output_imag_4_0(output_imag_5_0),
.output_real_5_0(output_real_6_0), .output_imag_5_0(output_imag_6_0),
.output_real_6_0(output_real_7_0), .output_imag_6_0(output_imag_7_0),
.output_real_7_0(output_real_8_0), .output_imag_7_0(output_imag_8_0),
.output_real_8_0(output_real_9_0), .output_imag_8_0(output_imag_9_0),
.output_real_9_0(output_real_10_0), .output_imag_9_0(output_imag_10_0),
.output_real_10_0(output_real_11_0), .output_imag_10_0(output_imag_11_0),
.output_real_11_0(output_real_12_0), .output_imag_11_0(output_imag_12_0),
.output_real_12_0(output_real_13_0), .output_imag_12_0(output_imag_13_0),
.output_real_13_0(output_real_14_0), .output_imag_13_0(output_imag_14_0),
.output_real_14_0(output_real_15_0), .output_imag_14_0(output_imag_15_0),
.output_real_15_0(output_real_16_0), .output_imag_15_0(output_imag_16_0),
.output_real_16_0(output_real_17_0), .output_imag_16_0(output_imag_17_0),
.output_real_17_0(output_real_18_0), .output_imag_17_0(output_imag_18_0),
.output_real_18_0(output_real_19_0), .output_imag_18_0(output_imag_19_0),
.output_real_19_0(output_real_20_0), .output_imag_19_0(output_imag_20_0),
.output_real_20_0(output_real_21_0), .output_imag_20_0(output_imag_21_0),
.output_real_21_0(output_real_22_0), .output_imag_21_0(output_imag_22_0),
.output_real_22_0(output_real_23_0), .output_imag_22_0(output_imag_23_0),
.output_real_23_0(output_real_24_0), .output_imag_23_0(output_imag_24_0),
.output_real_24_0(output_real_25_0), .output_imag_24_0(output_imag_25_0),
.output_real_25_0(output_real_26_0), .output_imag_25_0(output_imag_26_0),
.output_real_26_0(output_real_27_0), .output_imag_26_0(output_imag_27_0),
.output_real_27_0(output_real_28_0), .output_imag_27_0(output_imag_28_0),
.output_real_28_0(output_real_29_0), .output_imag_28_0(output_imag_29_0),
.output_real_29_0(output_real_30_0), .output_imag_29_0(output_imag_30_0),
.output_real_30_0(output_real_31_0), .output_imag_30_0(output_imag_31_0),
.output_real_31_0(output_real_32_0), .output_imag_31_0(output_imag_32_0),
.output_real_32_0(output_real_33_0), .output_imag_32_0(output_imag_33_0),
.output_real_33_0(output_real_34_0), .output_imag_33_0(output_imag_34_0),
.output_real_34_0(output_real_35_0), .output_imag_34_0(output_imag_35_0),
.output_real_35_0(output_real_36_0), .output_imag_35_0(output_imag_36_0),
.output_real_36_0(output_real_37_0), .output_imag_36_0(output_imag_37_0),
.output_real_37_0(output_real_38_0), .output_imag_37_0(output_imag_38_0),
.output_real_38_0(output_real_39_0), .output_imag_38_0(output_imag_39_0),
.output_real_39_0(output_real_40_0), .output_imag_39_0(output_imag_40_0),
.output_real_40_0(output_real_41_0), .output_imag_40_0(output_imag_41_0),
.output_real_41_0(output_real_42_0), .output_imag_41_0(output_imag_42_0),
.output_real_42_0(output_real_43_0), .output_imag_42_0(output_imag_43_0),
.output_real_43_0(output_real_44_0), .output_imag_43_0(output_imag_44_0),
.output_real_44_0(output_real_45_0), .output_imag_44_0(output_imag_45_0),
.output_real_45_0(output_real_46_0), .output_imag_45_0(output_imag_46_0),
.output_real_46_0(output_real_47_0), .output_imag_46_0(output_imag_47_0),
.output_real_47_0(output_real_48_0), .output_imag_47_0(output_imag_48_0),
.output_real_48_0(output_real_49_0), .output_imag_48_0(output_imag_49_0),
.output_real_49_0(output_real_50_0), .output_imag_49_0(output_imag_50_0),
.output_real_50_0(output_real_51_0), .output_imag_50_0(output_imag_51_0),
.output_real_51_0(output_real_52_0), .output_imag_51_0(output_imag_52_0),
.output_real_52_0(output_real_53_0), .output_imag_52_0(output_imag_53_0),
.output_real_53_0(output_real_54_0), .output_imag_53_0(output_imag_54_0),
.output_real_54_0(output_real_55_0), .output_imag_54_0(output_imag_55_0),
.output_real_55_0(output_real_56_0), .output_imag_55_0(output_imag_56_0),
.output_real_56_0(output_real_57_0), .output_imag_56_0(output_imag_57_0),
.output_real_57_0(output_real_58_0), .output_imag_57_0(output_imag_58_0),
.output_real_58_0(output_real_59_0), .output_imag_58_0(output_imag_59_0),
.output_real_59_0(output_real_60_0), .output_imag_59_0(output_imag_60_0),
.output_real_60_0(output_real_61_0), .output_imag_60_0(output_imag_61_0),
.output_real_61_0(output_real_62_0), .output_imag_61_0(output_imag_62_0),
.output_real_62_0(output_real_63_0), .output_imag_62_0(output_imag_63_0),
.output_real_63_0(output_real_64_0), .output_imag_63_0(output_imag_64_0),
.output_real_0_1(output_real_1_1), .output_imag_0_1(output_imag_1_1),
.output_real_1_1(output_real_2_1), .output_imag_1_1(output_imag_2_1),
.output_real_2_1(output_real_3_1), .output_imag_2_1(output_imag_3_1),
.output_real_3_1(output_real_4_1), .output_imag_3_1(output_imag_4_1),
.output_real_4_1(output_real_5_1), .output_imag_4_1(output_imag_5_1),
.output_real_5_1(output_real_6_1), .output_imag_5_1(output_imag_6_1),
.output_real_6_1(output_real_7_1), .output_imag_6_1(output_imag_7_1),
.output_real_7_1(output_real_8_1), .output_imag_7_1(output_imag_8_1),
.output_real_8_1(output_real_9_1), .output_imag_8_1(output_imag_9_1),
.output_real_9_1(output_real_10_1), .output_imag_9_1(output_imag_10_1),
.output_real_10_1(output_real_11_1), .output_imag_10_1(output_imag_11_1),
.output_real_11_1(output_real_12_1), .output_imag_11_1(output_imag_12_1),
.output_real_12_1(output_real_13_1), .output_imag_12_1(output_imag_13_1),
.output_real_13_1(output_real_14_1), .output_imag_13_1(output_imag_14_1),
.output_real_14_1(output_real_15_1), .output_imag_14_1(output_imag_15_1),
.output_real_15_1(output_real_16_1), .output_imag_15_1(output_imag_16_1),
.output_real_16_1(output_real_17_1), .output_imag_16_1(output_imag_17_1),
.output_real_17_1(output_real_18_1), .output_imag_17_1(output_imag_18_1),
.output_real_18_1(output_real_19_1), .output_imag_18_1(output_imag_19_1),
.output_real_19_1(output_real_20_1), .output_imag_19_1(output_imag_20_1),
.output_real_20_1(output_real_21_1), .output_imag_20_1(output_imag_21_1),
.output_real_21_1(output_real_22_1), .output_imag_21_1(output_imag_22_1),
.output_real_22_1(output_real_23_1), .output_imag_22_1(output_imag_23_1),
.output_real_23_1(output_real_24_1), .output_imag_23_1(output_imag_24_1),
.output_real_24_1(output_real_25_1), .output_imag_24_1(output_imag_25_1),
.output_real_25_1(output_real_26_1), .output_imag_25_1(output_imag_26_1),
.output_real_26_1(output_real_27_1), .output_imag_26_1(output_imag_27_1),
.output_real_27_1(output_real_28_1), .output_imag_27_1(output_imag_28_1),
.output_real_28_1(output_real_29_1), .output_imag_28_1(output_imag_29_1),
.output_real_29_1(output_real_30_1), .output_imag_29_1(output_imag_30_1),
.output_real_30_1(output_real_31_1), .output_imag_30_1(output_imag_31_1),
.output_real_31_1(output_real_32_1), .output_imag_31_1(output_imag_32_1),
.output_real_32_1(output_real_33_1), .output_imag_32_1(output_imag_33_1),
.output_real_33_1(output_real_34_1), .output_imag_33_1(output_imag_34_1),
.output_real_34_1(output_real_35_1), .output_imag_34_1(output_imag_35_1),
.output_real_35_1(output_real_36_1), .output_imag_35_1(output_imag_36_1),
.output_real_36_1(output_real_37_1), .output_imag_36_1(output_imag_37_1),
.output_real_37_1(output_real_38_1), .output_imag_37_1(output_imag_38_1),
.output_real_38_1(output_real_39_1), .output_imag_38_1(output_imag_39_1),
.output_real_39_1(output_real_40_1), .output_imag_39_1(output_imag_40_1),
.output_real_40_1(output_real_41_1), .output_imag_40_1(output_imag_41_1),
.output_real_41_1(output_real_42_1), .output_imag_41_1(output_imag_42_1),
.output_real_42_1(output_real_43_1), .output_imag_42_1(output_imag_43_1),
.output_real_43_1(output_real_44_1), .output_imag_43_1(output_imag_44_1),
.output_real_44_1(output_real_45_1), .output_imag_44_1(output_imag_45_1),
.output_real_45_1(output_real_46_1), .output_imag_45_1(output_imag_46_1),
.output_real_46_1(output_real_47_1), .output_imag_46_1(output_imag_47_1),
.output_real_47_1(output_real_48_1), .output_imag_47_1(output_imag_48_1),
.output_real_48_1(output_real_49_1), .output_imag_48_1(output_imag_49_1),
.output_real_49_1(output_real_50_1), .output_imag_49_1(output_imag_50_1),
.output_real_50_1(output_real_51_1), .output_imag_50_1(output_imag_51_1),
.output_real_51_1(output_real_52_1), .output_imag_51_1(output_imag_52_1),
.output_real_52_1(output_real_53_1), .output_imag_52_1(output_imag_53_1),
.output_real_53_1(output_real_54_1), .output_imag_53_1(output_imag_54_1),
.output_real_54_1(output_real_55_1), .output_imag_54_1(output_imag_55_1),
.output_real_55_1(output_real_56_1), .output_imag_55_1(output_imag_56_1),
.output_real_56_1(output_real_57_1), .output_imag_56_1(output_imag_57_1),
.output_real_57_1(output_real_58_1), .output_imag_57_1(output_imag_58_1),
.output_real_58_1(output_real_59_1), .output_imag_58_1(output_imag_59_1),
.output_real_59_1(output_real_60_1), .output_imag_59_1(output_imag_60_1),
.output_real_60_1(output_real_61_1), .output_imag_60_1(output_imag_61_1),
.output_real_61_1(output_real_62_1), .output_imag_61_1(output_imag_62_1),
.output_real_62_1(output_real_63_1), .output_imag_62_1(output_imag_63_1),
.output_real_63_1(output_real_64_1), .output_imag_63_1(output_imag_64_1),
.output_real_0_2(output_real_1_2), .output_imag_0_2(output_imag_1_2),
.output_real_1_2(output_real_2_2), .output_imag_1_2(output_imag_2_2),
.output_real_2_2(output_real_3_2), .output_imag_2_2(output_imag_3_2),
.output_real_3_2(output_real_4_2), .output_imag_3_2(output_imag_4_2),
.output_real_4_2(output_real_5_2), .output_imag_4_2(output_imag_5_2),
.output_real_5_2(output_real_6_2), .output_imag_5_2(output_imag_6_2),
.output_real_6_2(output_real_7_2), .output_imag_6_2(output_imag_7_2),
.output_real_7_2(output_real_8_2), .output_imag_7_2(output_imag_8_2),
.output_real_8_2(output_real_9_2), .output_imag_8_2(output_imag_9_2),
.output_real_9_2(output_real_10_2), .output_imag_9_2(output_imag_10_2),
.output_real_10_2(output_real_11_2), .output_imag_10_2(output_imag_11_2),
.output_real_11_2(output_real_12_2), .output_imag_11_2(output_imag_12_2),
.output_real_12_2(output_real_13_2), .output_imag_12_2(output_imag_13_2),
.output_real_13_2(output_real_14_2), .output_imag_13_2(output_imag_14_2),
.output_real_14_2(output_real_15_2), .output_imag_14_2(output_imag_15_2),
.output_real_15_2(output_real_16_2), .output_imag_15_2(output_imag_16_2),
.output_real_16_2(output_real_17_2), .output_imag_16_2(output_imag_17_2),
.output_real_17_2(output_real_18_2), .output_imag_17_2(output_imag_18_2),
.output_real_18_2(output_real_19_2), .output_imag_18_2(output_imag_19_2),
.output_real_19_2(output_real_20_2), .output_imag_19_2(output_imag_20_2),
.output_real_20_2(output_real_21_2), .output_imag_20_2(output_imag_21_2),
.output_real_21_2(output_real_22_2), .output_imag_21_2(output_imag_22_2),
.output_real_22_2(output_real_23_2), .output_imag_22_2(output_imag_23_2),
.output_real_23_2(output_real_24_2), .output_imag_23_2(output_imag_24_2),
.output_real_24_2(output_real_25_2), .output_imag_24_2(output_imag_25_2),
.output_real_25_2(output_real_26_2), .output_imag_25_2(output_imag_26_2),
.output_real_26_2(output_real_27_2), .output_imag_26_2(output_imag_27_2),
.output_real_27_2(output_real_28_2), .output_imag_27_2(output_imag_28_2),
.output_real_28_2(output_real_29_2), .output_imag_28_2(output_imag_29_2),
.output_real_29_2(output_real_30_2), .output_imag_29_2(output_imag_30_2),
.output_real_30_2(output_real_31_2), .output_imag_30_2(output_imag_31_2),
.output_real_31_2(output_real_32_2), .output_imag_31_2(output_imag_32_2),
.output_real_32_2(output_real_33_2), .output_imag_32_2(output_imag_33_2),
.output_real_33_2(output_real_34_2), .output_imag_33_2(output_imag_34_2),
.output_real_34_2(output_real_35_2), .output_imag_34_2(output_imag_35_2),
.output_real_35_2(output_real_36_2), .output_imag_35_2(output_imag_36_2),
.output_real_36_2(output_real_37_2), .output_imag_36_2(output_imag_37_2),
.output_real_37_2(output_real_38_2), .output_imag_37_2(output_imag_38_2),
.output_real_38_2(output_real_39_2), .output_imag_38_2(output_imag_39_2),
.output_real_39_2(output_real_40_2), .output_imag_39_2(output_imag_40_2),
.output_real_40_2(output_real_41_2), .output_imag_40_2(output_imag_41_2),
.output_real_41_2(output_real_42_2), .output_imag_41_2(output_imag_42_2),
.output_real_42_2(output_real_43_2), .output_imag_42_2(output_imag_43_2),
.output_real_43_2(output_real_44_2), .output_imag_43_2(output_imag_44_2),
.output_real_44_2(output_real_45_2), .output_imag_44_2(output_imag_45_2),
.output_real_45_2(output_real_46_2), .output_imag_45_2(output_imag_46_2),
.output_real_46_2(output_real_47_2), .output_imag_46_2(output_imag_47_2),
.output_real_47_2(output_real_48_2), .output_imag_47_2(output_imag_48_2),
.output_real_48_2(output_real_49_2), .output_imag_48_2(output_imag_49_2),
.output_real_49_2(output_real_50_2), .output_imag_49_2(output_imag_50_2),
.output_real_50_2(output_real_51_2), .output_imag_50_2(output_imag_51_2),
.output_real_51_2(output_real_52_2), .output_imag_51_2(output_imag_52_2),
.output_real_52_2(output_real_53_2), .output_imag_52_2(output_imag_53_2),
.output_real_53_2(output_real_54_2), .output_imag_53_2(output_imag_54_2),
.output_real_54_2(output_real_55_2), .output_imag_54_2(output_imag_55_2),
.output_real_55_2(output_real_56_2), .output_imag_55_2(output_imag_56_2),
.output_real_56_2(output_real_57_2), .output_imag_56_2(output_imag_57_2),
.output_real_57_2(output_real_58_2), .output_imag_57_2(output_imag_58_2),
.output_real_58_2(output_real_59_2), .output_imag_58_2(output_imag_59_2),
.output_real_59_2(output_real_60_2), .output_imag_59_2(output_imag_60_2),
.output_real_60_2(output_real_61_2), .output_imag_60_2(output_imag_61_2),
.output_real_61_2(output_real_62_2), .output_imag_61_2(output_imag_62_2),
.output_real_62_2(output_real_63_2), .output_imag_62_2(output_imag_63_2),
.output_real_63_2(output_real_64_2), .output_imag_63_2(output_imag_64_2),
.output_real_0_3(output_real_1_3), .output_imag_0_3(output_imag_1_3),
.output_real_1_3(output_real_2_3), .output_imag_1_3(output_imag_2_3),
.output_real_2_3(output_real_3_3), .output_imag_2_3(output_imag_3_3),
.output_real_3_3(output_real_4_3), .output_imag_3_3(output_imag_4_3),
.output_real_4_3(output_real_5_3), .output_imag_4_3(output_imag_5_3),
.output_real_5_3(output_real_6_3), .output_imag_5_3(output_imag_6_3),
.output_real_6_3(output_real_7_3), .output_imag_6_3(output_imag_7_3),
.output_real_7_3(output_real_8_3), .output_imag_7_3(output_imag_8_3),
.output_real_8_3(output_real_9_3), .output_imag_8_3(output_imag_9_3),
.output_real_9_3(output_real_10_3), .output_imag_9_3(output_imag_10_3),
.output_real_10_3(output_real_11_3), .output_imag_10_3(output_imag_11_3),
.output_real_11_3(output_real_12_3), .output_imag_11_3(output_imag_12_3),
.output_real_12_3(output_real_13_3), .output_imag_12_3(output_imag_13_3),
.output_real_13_3(output_real_14_3), .output_imag_13_3(output_imag_14_3),
.output_real_14_3(output_real_15_3), .output_imag_14_3(output_imag_15_3),
.output_real_15_3(output_real_16_3), .output_imag_15_3(output_imag_16_3),
.output_real_16_3(output_real_17_3), .output_imag_16_3(output_imag_17_3),
.output_real_17_3(output_real_18_3), .output_imag_17_3(output_imag_18_3),
.output_real_18_3(output_real_19_3), .output_imag_18_3(output_imag_19_3),
.output_real_19_3(output_real_20_3), .output_imag_19_3(output_imag_20_3),
.output_real_20_3(output_real_21_3), .output_imag_20_3(output_imag_21_3),
.output_real_21_3(output_real_22_3), .output_imag_21_3(output_imag_22_3),
.output_real_22_3(output_real_23_3), .output_imag_22_3(output_imag_23_3),
.output_real_23_3(output_real_24_3), .output_imag_23_3(output_imag_24_3),
.output_real_24_3(output_real_25_3), .output_imag_24_3(output_imag_25_3),
.output_real_25_3(output_real_26_3), .output_imag_25_3(output_imag_26_3),
.output_real_26_3(output_real_27_3), .output_imag_26_3(output_imag_27_3),
.output_real_27_3(output_real_28_3), .output_imag_27_3(output_imag_28_3),
.output_real_28_3(output_real_29_3), .output_imag_28_3(output_imag_29_3),
.output_real_29_3(output_real_30_3), .output_imag_29_3(output_imag_30_3),
.output_real_30_3(output_real_31_3), .output_imag_30_3(output_imag_31_3),
.output_real_31_3(output_real_32_3), .output_imag_31_3(output_imag_32_3),
.output_real_32_3(output_real_33_3), .output_imag_32_3(output_imag_33_3),
.output_real_33_3(output_real_34_3), .output_imag_33_3(output_imag_34_3),
.output_real_34_3(output_real_35_3), .output_imag_34_3(output_imag_35_3),
.output_real_35_3(output_real_36_3), .output_imag_35_3(output_imag_36_3),
.output_real_36_3(output_real_37_3), .output_imag_36_3(output_imag_37_3),
.output_real_37_3(output_real_38_3), .output_imag_37_3(output_imag_38_3),
.output_real_38_3(output_real_39_3), .output_imag_38_3(output_imag_39_3),
.output_real_39_3(output_real_40_3), .output_imag_39_3(output_imag_40_3),
.output_real_40_3(output_real_41_3), .output_imag_40_3(output_imag_41_3),
.output_real_41_3(output_real_42_3), .output_imag_41_3(output_imag_42_3),
.output_real_42_3(output_real_43_3), .output_imag_42_3(output_imag_43_3),
.output_real_43_3(output_real_44_3), .output_imag_43_3(output_imag_44_3),
.output_real_44_3(output_real_45_3), .output_imag_44_3(output_imag_45_3),
.output_real_45_3(output_real_46_3), .output_imag_45_3(output_imag_46_3),
.output_real_46_3(output_real_47_3), .output_imag_46_3(output_imag_47_3),
.output_real_47_3(output_real_48_3), .output_imag_47_3(output_imag_48_3),
.output_real_48_3(output_real_49_3), .output_imag_48_3(output_imag_49_3),
.output_real_49_3(output_real_50_3), .output_imag_49_3(output_imag_50_3),
.output_real_50_3(output_real_51_3), .output_imag_50_3(output_imag_51_3),
.output_real_51_3(output_real_52_3), .output_imag_51_3(output_imag_52_3),
.output_real_52_3(output_real_53_3), .output_imag_52_3(output_imag_53_3),
.output_real_53_3(output_real_54_3), .output_imag_53_3(output_imag_54_3),
.output_real_54_3(output_real_55_3), .output_imag_54_3(output_imag_55_3),
.output_real_55_3(output_real_56_3), .output_imag_55_3(output_imag_56_3),
.output_real_56_3(output_real_57_3), .output_imag_56_3(output_imag_57_3),
.output_real_57_3(output_real_58_3), .output_imag_57_3(output_imag_58_3),
.output_real_58_3(output_real_59_3), .output_imag_58_3(output_imag_59_3),
.output_real_59_3(output_real_60_3), .output_imag_59_3(output_imag_60_3),
.output_real_60_3(output_real_61_3), .output_imag_60_3(output_imag_61_3),
.output_real_61_3(output_real_62_3), .output_imag_61_3(output_imag_62_3),
.output_real_62_3(output_real_63_3), .output_imag_62_3(output_imag_63_3),
.output_real_63_3(output_real_64_3), .output_imag_63_3(output_imag_64_3),
.ssb(ssb),
.sdi(sdi),
.vmm_load(vmm_load),
.CLK(CLK),
.rst(rst)
);


vmm_adder DUT_VMM_ADDER0(
.CLK(CLK),               
.rst(rst), 
.input_a_real1_vmm0(output_data_divider1[31:16]), .input_a_real2_vmm0(output_data_divider2[31:16]), .input_a_real3_vmm0(output_data_divider3[31:16]), .input_a_real4_vmm0(output_data_divider4[31:16]),
.input_a_imag1_vmm0(output_data_divider1[15:0]),  .input_a_imag2_vmm0(output_data_divider2[15:0]),  .input_a_imag3_vmm0(output_data_divider3[15:0]),  .input_a_imag4_vmm0(output_data_divider4[15:0]),  
.input_a_real5_vmm0(output_data_divider5[31:16]), .input_a_real6_vmm0(output_data_divider6[31:16]), .input_a_real7_vmm0(output_data_divider7[31:16]), .input_a_real8_vmm0(output_data_divider8[31:16]),
.input_a_imag5_vmm0(output_data_divider5[15:0]),  .input_a_imag6_vmm0(output_data_divider6[15:0]),  .input_a_imag7_vmm0(output_data_divider7[15:0]),  .input_a_imag8_vmm0(output_data_divider8[15:0]),  
.input_a_real9_vmm0(output_data_divider9[31:16]), .input_a_real10_vmm0(output_data_divider10[31:16]), .input_a_real11_vmm0(output_data_divider11[31:16]), .input_a_real12_vmm0(output_data_divider12[31:16]),
.input_a_imag9_vmm0(output_data_divider9[15:0]),  .input_a_imag10_vmm0(output_data_divider10[15:0]),  .input_a_imag11_vmm0(output_data_divider11[15:0]),  .input_a_imag12_vmm0(output_data_divider12[15:0]),  
.input_a_real13_vmm0(output_data_divider13[31:16]), .input_a_real14_vmm0(output_data_divider14[31:16]), .input_a_real15_vmm0(output_data_divider15[31:16]), .input_a_real16_vmm0(output_data_divider16[31:16]),
.input_a_imag13_vmm0(output_data_divider13[15:0]),  .input_a_imag14_vmm0(output_data_divider14[15:0]),  .input_a_imag15_vmm0(output_data_divider15[15:0]),  .input_a_imag16_vmm0(output_data_divider16[15:0]),  
.input_a_real1_vmm1(output_data_divider17[31:16]), .input_a_real2_vmm1(output_data_divider18[31:16]), .input_a_real3_vmm1(output_data_divider19[31:16]), .input_a_real4_vmm1(output_data_divider20[31:16]),
.input_a_imag1_vmm1(output_data_divider17[15:0]),  .input_a_imag2_vmm1(output_data_divider18[15:0]),  .input_a_imag3_vmm1(output_data_divider19[15:0]),  .input_a_imag4_vmm1(output_data_divider20[15:0]),  
.input_a_real5_vmm1(output_data_divider21[31:16]), .input_a_real6_vmm1(output_data_divider22[31:16]), .input_a_real7_vmm1(output_data_divider23[31:16]), .input_a_real8_vmm1(output_data_divider24[31:16]),
.input_a_imag5_vmm1(output_data_divider21[15:0]),  .input_a_imag6_vmm1(output_data_divider22[15:0]),  .input_a_imag7_vmm1(output_data_divider23[15:0]),  .input_a_imag8_vmm1(output_data_divider24[15:0]),  
.input_a_real9_vmm1(output_data_divider25[31:16]), .input_a_real10_vmm1(output_data_divider26[31:16]), .input_a_real11_vmm1(output_data_divider27[31:16]), .input_a_real12_vmm1(output_data_divider28[31:16]),
.input_a_imag9_vmm1(output_data_divider25[15:0]),  .input_a_imag10_vmm1(output_data_divider26[15:0]),  .input_a_imag11_vmm1(output_data_divider27[15:0]),  .input_a_imag12_vmm1(output_data_divider28[15:0]),  
.input_a_real13_vmm1(output_data_divider29[31:16]), .input_a_real14_vmm1(output_data_divider30[31:16]), .input_a_real15_vmm1(output_data_divider31[31:16]), .input_a_real16_vmm1(output_data_divider32[31:16]),
.input_a_imag13_vmm1(output_data_divider29[15:0]),  .input_a_imag14_vmm1(output_data_divider30[15:0]),  .input_a_imag15_vmm1(output_data_divider31[15:0]),  .input_a_imag16_vmm1(output_data_divider32[15:0]),  
.input_a_real1_vmm2(output_data_divider33[31:16]), .input_a_real2_vmm2(output_data_divider34[31:16]), .input_a_real3_vmm2(output_data_divider35[31:16]), .input_a_real4_vmm2(output_data_divider36[31:16]),
.input_a_imag1_vmm2(output_data_divider33[15:0]),  .input_a_imag2_vmm2(output_data_divider34[15:0]),  .input_a_imag3_vmm2(output_data_divider35[15:0]),  .input_a_imag4_vmm2(output_data_divider36[15:0]),  
.input_a_real5_vmm2(output_data_divider37[31:16]), .input_a_real6_vmm2(output_data_divider38[31:16]), .input_a_real7_vmm2(output_data_divider39[31:16]), .input_a_real8_vmm2(output_data_divider40[31:16]),
.input_a_imag5_vmm2(output_data_divider37[15:0]),  .input_a_imag6_vmm2(output_data_divider38[15:0]),  .input_a_imag7_vmm2(output_data_divider39[15:0]),  .input_a_imag8_vmm2(output_data_divider40[15:0]),  
.input_a_real9_vmm2(output_data_divider41[31:16]), .input_a_real10_vmm2(output_data_divider42[31:16]), .input_a_real11_vmm2(output_data_divider43[31:16]), .input_a_real12_vmm2(output_data_divider44[31:16]),
.input_a_imag9_vmm2(output_data_divider41[15:0]),  .input_a_imag10_vmm2(output_data_divider42[15:0]),  .input_a_imag11_vmm2(output_data_divider43[15:0]),  .input_a_imag12_vmm2(output_data_divider44[15:0]),  
.input_a_real13_vmm2(output_data_divider45[31:16]), .input_a_real14_vmm2(output_data_divider46[31:16]), .input_a_real15_vmm2(output_data_divider47[31:16]), .input_a_real16_vmm2(output_data_divider48[31:16]),
.input_a_imag13_vmm2(output_data_divider45[15:0]),  .input_a_imag14_vmm2(output_data_divider46[15:0]),  .input_a_imag15_vmm2(output_data_divider47[15:0]),  .input_a_imag16_vmm2(output_data_divider48[15:0]),  
.input_a_real1_vmm3(output_data_divider49[31:16]), .input_a_real2_vmm3(output_data_divider50[31:16]), .input_a_real3_vmm3(output_data_divider51[31:16]), .input_a_real4_vmm3(output_data_divider52[31:16]),
.input_a_imag1_vmm3(output_data_divider49[15:0]),  .input_a_imag2_vmm3(output_data_divider50[15:0]),  .input_a_imag3_vmm3(output_data_divider51[15:0]),  .input_a_imag4_vmm3(output_data_divider52[15:0]),  
.input_a_real5_vmm3(output_data_divider53[31:16]), .input_a_real6_vmm3(output_data_divider54[31:16]), .input_a_real7_vmm3(output_data_divider55[31:16]), .input_a_real8_vmm3(output_data_divider56[31:16]),
.input_a_imag5_vmm3(output_data_divider53[15:0]),  .input_a_imag6_vmm3(output_data_divider54[15:0]),  .input_a_imag7_vmm3(output_data_divider55[15:0]),  .input_a_imag8_vmm3(output_data_divider56[15:0]),  
.input_a_real9_vmm3(output_data_divider57[31:16]), .input_a_real10_vmm3(output_data_divider58[31:16]), .input_a_real11_vmm3(output_data_divider59[31:16]), .input_a_real12_vmm3(output_data_divider60[31:16]),
.input_a_imag9_vmm3(output_data_divider57[15:0]),  .input_a_imag10_vmm3(output_data_divider58[15:0]),  .input_a_imag11_vmm3(output_data_divider59[15:0]),  .input_a_imag12_vmm3(output_data_divider60[15:0]),  
.input_a_real13_vmm3(output_data_divider61[31:16]), .input_a_real14_vmm3(output_data_divider62[31:16]), .input_a_real15_vmm3(output_data_divider63[31:16]), .input_a_real16_vmm3(output_data_divider64[31:16]),
.input_a_imag13_vmm3(output_data_divider61[15:0]),  .input_a_imag14_vmm3(output_data_divider62[15:0]),  .input_a_imag15_vmm3(output_data_divider63[15:0]),  .input_a_imag16_vmm3(output_data_divider64[15:0]), 
.input_b_real1_vmm0(output_real_1_0), .input_b_real2_vmm0(output_real_2_0), .input_b_real3_vmm0(output_real_3_0), .input_b_real4_vmm0(output_real_4_0),
.input_b_imag1_vmm0(output_imag_1_0),   .input_b_imag2_vmm0(output_imag_2_0),   .input_b_imag3_vmm0(output_imag_3_0),   .input_b_imag4_vmm0(output_imag_4_0),  
.input_b_real5_vmm0(output_real_5_0), .input_b_real6_vmm0(output_real_6_0), .input_b_real7_vmm0(output_real_7_0), .input_b_real8_vmm0(output_real_8_0),
.input_b_imag5_vmm0(output_imag_5_0),   .input_b_imag6_vmm0(output_imag_6_0),   .input_b_imag7_vmm0(output_imag_7_0),   .input_b_imag8_vmm0(output_imag_8_0),  
.input_b_real9_vmm0(output_real_9_0), .input_b_real10_vmm0(output_real_10_0), .input_b_real11_vmm0(output_real_11_0), .input_b_real12_vmm0(output_real_12_0),
.input_b_imag9_vmm0(output_imag_9_0),   .input_b_imag10_vmm0(output_imag_10_0),   .input_b_imag11_vmm0(output_imag_11_0),   .input_b_imag12_vmm0(output_imag_12_0),  
.input_b_real13_vmm0(output_real_13_0), .input_b_real14_vmm0(output_real_14_0), .input_b_real15_vmm0(output_real_15_0), .input_b_real16_vmm0(output_real_16_0),
.input_b_imag13_vmm0(output_imag_13_0),   .input_b_imag14_vmm0(output_imag_14_0),   .input_b_imag15_vmm0(output_imag_15_0),   .input_b_imag16_vmm0(output_imag_16_0),  
.input_b_real1_vmm1(output_real_17_0), .input_b_real2_vmm1(output_real_18_0), .input_b_real3_vmm1(output_real_19_0), .input_b_real4_vmm1(output_real_20_0),
.input_b_imag1_vmm1(output_imag_17_0),   .input_b_imag2_vmm1(output_imag_18_0),   .input_b_imag3_vmm1(output_imag_19_0),   .input_b_imag4_vmm1(output_imag_20_0),  
.input_b_real5_vmm1(output_real_21_0), .input_b_real6_vmm1(output_real_22_0), .input_b_real7_vmm1(output_real_23_0), .input_b_real8_vmm1(output_real_24_0),
.input_b_imag5_vmm1(output_imag_21_0),   .input_b_imag6_vmm1(output_imag_22_0),   .input_b_imag7_vmm1(output_imag_23_0),   .input_b_imag8_vmm1(output_imag_24_0),  
.input_b_real9_vmm1(output_real_25_0), .input_b_real10_vmm1(output_real_26_0), .input_b_real11_vmm1(output_real_27_0), .input_b_real12_vmm1(output_real_28_0),
.input_b_imag9_vmm1(output_imag_25_0),   .input_b_imag10_vmm1(output_imag_26_0),   .input_b_imag11_vmm1(output_imag_27_0),   .input_b_imag12_vmm1(output_imag_28_0),  
.input_b_real13_vmm1(output_real_29_0), .input_b_real14_vmm1(output_real_30_0), .input_b_real15_vmm1(output_real_31_0), .input_b_real16_vmm1(output_real_32_0),
.input_b_imag13_vmm1(output_imag_29_0),   .input_b_imag14_vmm1(output_imag_30_0),   .input_b_imag15_vmm1(output_imag_31_0),   .input_b_imag16_vmm1(output_imag_32_0),  
.input_b_real1_vmm2(output_real_33_0), .input_b_real2_vmm2(output_real_34_0), .input_b_real3_vmm2(output_real_35_0), .input_b_real4_vmm2(output_real_36_0),
.input_b_imag1_vmm2(output_imag_33_0),   .input_b_imag2_vmm2(output_imag_34_0),   .input_b_imag3_vmm2(output_imag_35_0),   .input_b_imag4_vmm2(output_imag_36_0),  
.input_b_real5_vmm2(output_real_37_0), .input_b_real6_vmm2(output_real_38_0), .input_b_real7_vmm2(output_real_39_0), .input_b_real8_vmm2(output_real_40_0),
.input_b_imag5_vmm2(output_imag_37_0),   .input_b_imag6_vmm2(output_imag_38_0),   .input_b_imag7_vmm2(output_imag_39_0),   .input_b_imag8_vmm2(output_imag_40_0),  
.input_b_real9_vmm2(output_real_41_0), .input_b_real10_vmm2(output_real_42_0), .input_b_real11_vmm2(output_real_43_0), .input_b_real12_vmm2(output_real_44_0),
.input_b_imag9_vmm2(output_imag_41_0),   .input_b_imag10_vmm2(output_imag_42_0),   .input_b_imag11_vmm2(output_imag_43_0),   .input_b_imag12_vmm2(output_imag_44_0),  
.input_b_real13_vmm2(output_real_45_0), .input_b_real14_vmm2(output_real_46_0), .input_b_real15_vmm2(output_real_47_0), .input_b_real16_vmm2(output_real_48_0),
.input_b_imag13_vmm2(output_imag_45_0),   .input_b_imag14_vmm2(output_imag_46_0),   .input_b_imag15_vmm2(output_imag_47_0),   .input_b_imag16_vmm2(output_imag_48_0),  
.input_b_real1_vmm3(output_real_49_0), .input_b_real2_vmm3(output_real_50_0), .input_b_real3_vmm3(output_real_51_0), .input_b_real4_vmm3(output_real_52_0),
.input_b_imag1_vmm3(output_imag_49_0),   .input_b_imag2_vmm3(output_imag_50_0),   .input_b_imag3_vmm3(output_imag_51_0),   .input_b_imag4_vmm3(output_imag_52_0),  
.input_b_real5_vmm3(output_real_53_0), .input_b_real6_vmm3(output_real_54_0), .input_b_real7_vmm3(output_real_55_0), .input_b_real8_vmm3(output_real_56_0),
.input_b_imag5_vmm3(output_imag_53_0),   .input_b_imag6_vmm3(output_imag_54_0),   .input_b_imag7_vmm3(output_imag_55_0),   .input_b_imag8_vmm3(output_imag_56_0),  
.input_b_real9_vmm3(output_real_57_0), .input_b_real10_vmm3(output_real_58_0), .input_b_real11_vmm3(output_real_59_0), .input_b_real12_vmm3(output_real_60_0),
.input_b_imag9_vmm3(output_imag_57_0),   .input_b_imag10_vmm3(output_imag_58_0),   .input_b_imag11_vmm3(output_imag_59_0),   .input_b_imag12_vmm3(output_imag_60_0),  
.input_b_real13_vmm3(output_real_61_0), .input_b_real14_vmm3(output_real_62_0), .input_b_real15_vmm3(output_real_63_0), .input_b_real16_vmm3(output_real_64_0),
.input_b_imag13_vmm3(output_imag_61_0),   .input_b_imag14_vmm3(output_imag_62_0),   .input_b_imag15_vmm3(output_imag_63_0),   .input_b_imag16_vmm3(output_imag_64_0),  
.output_z_real(output_z_real1_0),
.output_z_imag(output_z_imag1_0)
);

vmm_adder DUT_VMM_ADDER1(
.CLK(CLK),               
.rst(rst), 
.input_a_real1_vmm0(output_data_divider1[31:16]), .input_a_real2_vmm0(output_data_divider2[31:16]), .input_a_real3_vmm0(output_data_divider3[31:16]), .input_a_real4_vmm0(output_data_divider4[31:16]),
.input_a_imag1_vmm0(output_data_divider1[15:0]),  .input_a_imag2_vmm0(output_data_divider2[15:0]),  .input_a_imag3_vmm0(output_data_divider3[15:0]),  .input_a_imag4_vmm0(output_data_divider4[15:0]),  
.input_a_real5_vmm0(output_data_divider5[31:16]), .input_a_real6_vmm0(output_data_divider6[31:16]), .input_a_real7_vmm0(output_data_divider7[31:16]), .input_a_real8_vmm0(output_data_divider8[31:16]),
.input_a_imag5_vmm0(output_data_divider5[15:0]),  .input_a_imag6_vmm0(output_data_divider6[15:0]),  .input_a_imag7_vmm0(output_data_divider7[15:0]),  .input_a_imag8_vmm0(output_data_divider8[15:0]),  
.input_a_real9_vmm0(output_data_divider9[31:16]), .input_a_real10_vmm0(output_data_divider10[31:16]), .input_a_real11_vmm0(output_data_divider11[31:16]), .input_a_real12_vmm0(output_data_divider12[31:16]),
.input_a_imag9_vmm0(output_data_divider9[15:0]),  .input_a_imag10_vmm0(output_data_divider10[15:0]),  .input_a_imag11_vmm0(output_data_divider11[15:0]),  .input_a_imag12_vmm0(output_data_divider12[15:0]),  
.input_a_real13_vmm0(output_data_divider13[31:16]), .input_a_real14_vmm0(output_data_divider14[31:16]), .input_a_real15_vmm0(output_data_divider15[31:16]), .input_a_real16_vmm0(output_data_divider16[31:16]),
.input_a_imag13_vmm0(output_data_divider13[15:0]),  .input_a_imag14_vmm0(output_data_divider14[15:0]),  .input_a_imag15_vmm0(output_data_divider15[15:0]),  .input_a_imag16_vmm0(output_data_divider16[15:0]),  
.input_a_real1_vmm1(output_data_divider17[31:16]), .input_a_real2_vmm1(output_data_divider18[31:16]), .input_a_real3_vmm1(output_data_divider19[31:16]), .input_a_real4_vmm1(output_data_divider20[31:16]),
.input_a_imag1_vmm1(output_data_divider17[15:0]),  .input_a_imag2_vmm1(output_data_divider18[15:0]),  .input_a_imag3_vmm1(output_data_divider19[15:0]),  .input_a_imag4_vmm1(output_data_divider20[15:0]),  
.input_a_real5_vmm1(output_data_divider21[31:16]), .input_a_real6_vmm1(output_data_divider22[31:16]), .input_a_real7_vmm1(output_data_divider23[31:16]), .input_a_real8_vmm1(output_data_divider24[31:16]),
.input_a_imag5_vmm1(output_data_divider21[15:0]),  .input_a_imag6_vmm1(output_data_divider22[15:0]),  .input_a_imag7_vmm1(output_data_divider23[15:0]),  .input_a_imag8_vmm1(output_data_divider24[15:0]),  
.input_a_real9_vmm1(output_data_divider25[31:16]), .input_a_real10_vmm1(output_data_divider26[31:16]), .input_a_real11_vmm1(output_data_divider27[31:16]), .input_a_real12_vmm1(output_data_divider28[31:16]),
.input_a_imag9_vmm1(output_data_divider25[15:0]),  .input_a_imag10_vmm1(output_data_divider26[15:0]),  .input_a_imag11_vmm1(output_data_divider27[15:0]),  .input_a_imag12_vmm1(output_data_divider28[15:0]),  
.input_a_real13_vmm1(output_data_divider29[31:16]), .input_a_real14_vmm1(output_data_divider30[31:16]), .input_a_real15_vmm1(output_data_divider31[31:16]), .input_a_real16_vmm1(output_data_divider32[31:16]),
.input_a_imag13_vmm1(output_data_divider29[15:0]),  .input_a_imag14_vmm1(output_data_divider30[15:0]),  .input_a_imag15_vmm1(output_data_divider31[15:0]),  .input_a_imag16_vmm1(output_data_divider32[15:0]),  
.input_a_real1_vmm2(output_data_divider33[31:16]), .input_a_real2_vmm2(output_data_divider34[31:16]), .input_a_real3_vmm2(output_data_divider35[31:16]), .input_a_real4_vmm2(output_data_divider36[31:16]),
.input_a_imag1_vmm2(output_data_divider33[15:0]),  .input_a_imag2_vmm2(output_data_divider34[15:0]),  .input_a_imag3_vmm2(output_data_divider35[15:0]),  .input_a_imag4_vmm2(output_data_divider36[15:0]),  
.input_a_real5_vmm2(output_data_divider37[31:16]), .input_a_real6_vmm2(output_data_divider38[31:16]), .input_a_real7_vmm2(output_data_divider39[31:16]), .input_a_real8_vmm2(output_data_divider40[31:16]),
.input_a_imag5_vmm2(output_data_divider37[15:0]),  .input_a_imag6_vmm2(output_data_divider38[15:0]),  .input_a_imag7_vmm2(output_data_divider39[15:0]),  .input_a_imag8_vmm2(output_data_divider40[15:0]),  
.input_a_real9_vmm2(output_data_divider41[31:16]), .input_a_real10_vmm2(output_data_divider42[31:16]), .input_a_real11_vmm2(output_data_divider43[31:16]), .input_a_real12_vmm2(output_data_divider44[31:16]),
.input_a_imag9_vmm2(output_data_divider41[15:0]),  .input_a_imag10_vmm2(output_data_divider42[15:0]),  .input_a_imag11_vmm2(output_data_divider43[15:0]),  .input_a_imag12_vmm2(output_data_divider44[15:0]),  
.input_a_real13_vmm2(output_data_divider45[31:16]), .input_a_real14_vmm2(output_data_divider46[31:16]), .input_a_real15_vmm2(output_data_divider47[31:16]), .input_a_real16_vmm2(output_data_divider48[31:16]),
.input_a_imag13_vmm2(output_data_divider45[15:0]),  .input_a_imag14_vmm2(output_data_divider46[15:0]),  .input_a_imag15_vmm2(output_data_divider47[15:0]),  .input_a_imag16_vmm2(output_data_divider48[15:0]),  
.input_a_real1_vmm3(output_data_divider49[31:16]), .input_a_real2_vmm3(output_data_divider50[31:16]), .input_a_real3_vmm3(output_data_divider51[31:16]), .input_a_real4_vmm3(output_data_divider52[31:16]),
.input_a_imag1_vmm3(output_data_divider49[15:0]),  .input_a_imag2_vmm3(output_data_divider50[15:0]),  .input_a_imag3_vmm3(output_data_divider51[15:0]),  .input_a_imag4_vmm3(output_data_divider52[15:0]),  
.input_a_real5_vmm3(output_data_divider53[31:16]), .input_a_real6_vmm3(output_data_divider54[31:16]), .input_a_real7_vmm3(output_data_divider55[31:16]), .input_a_real8_vmm3(output_data_divider56[31:16]),
.input_a_imag5_vmm3(output_data_divider53[15:0]),  .input_a_imag6_vmm3(output_data_divider54[15:0]),  .input_a_imag7_vmm3(output_data_divider55[15:0]),  .input_a_imag8_vmm3(output_data_divider56[15:0]),  
.input_a_real9_vmm3(output_data_divider57[31:16]), .input_a_real10_vmm3(output_data_divider58[31:16]), .input_a_real11_vmm3(output_data_divider59[31:16]), .input_a_real12_vmm3(output_data_divider60[31:16]),
.input_a_imag9_vmm3(output_data_divider57[15:0]),  .input_a_imag10_vmm3(output_data_divider58[15:0]),  .input_a_imag11_vmm3(output_data_divider59[15:0]),  .input_a_imag12_vmm3(output_data_divider60[15:0]),  
.input_a_real13_vmm3(output_data_divider61[31:16]), .input_a_real14_vmm3(output_data_divider62[31:16]), .input_a_real15_vmm3(output_data_divider63[31:16]), .input_a_real16_vmm3(output_data_divider64[31:16]),
.input_a_imag13_vmm3(output_data_divider61[15:0]),  .input_a_imag14_vmm3(output_data_divider62[15:0]),  .input_a_imag15_vmm3(output_data_divider63[15:0]),  .input_a_imag16_vmm3(output_data_divider64[15:0]),   
.input_b_real1_vmm0(output_real_1_1), .input_b_real2_vmm0(output_real_2_1), .input_b_real3_vmm0(output_real_3_1), .input_b_real4_vmm0(output_real_4_1),
.input_b_imag1_vmm0(output_imag_1_1),   .input_b_imag2_vmm0(output_imag_2_1),   .input_b_imag3_vmm0(output_imag_3_1),   .input_b_imag4_vmm0(output_imag_4_1),  
.input_b_real5_vmm0(output_real_5_1), .input_b_real6_vmm0(output_real_6_1), .input_b_real7_vmm0(output_real_7_1), .input_b_real8_vmm0(output_real_8_1),
.input_b_imag5_vmm0(output_imag_5_1),   .input_b_imag6_vmm0(output_imag_6_1),   .input_b_imag7_vmm0(output_imag_7_1),   .input_b_imag8_vmm0(output_imag_8_1),  
.input_b_real9_vmm0(output_real_9_1), .input_b_real10_vmm0(output_real_10_1), .input_b_real11_vmm0(output_real_11_1), .input_b_real12_vmm0(output_real_12_1),
.input_b_imag9_vmm0(output_imag_9_1),   .input_b_imag10_vmm0(output_imag_10_1),   .input_b_imag11_vmm0(output_imag_11_1),   .input_b_imag12_vmm0(output_imag_12_1),  
.input_b_real13_vmm0(output_real_13_1), .input_b_real14_vmm0(output_real_14_1), .input_b_real15_vmm0(output_real_15_1), .input_b_real16_vmm0(output_real_16_1),
.input_b_imag13_vmm0(output_imag_13_1),   .input_b_imag14_vmm0(output_imag_14_1),   .input_b_imag15_vmm0(output_imag_15_1),   .input_b_imag16_vmm0(output_imag_16_1),  
.input_b_real1_vmm1(output_real_17_1), .input_b_real2_vmm1(output_real_18_1), .input_b_real3_vmm1(output_real_19_1), .input_b_real4_vmm1(output_real_20_1),
.input_b_imag1_vmm1(output_imag_17_1),   .input_b_imag2_vmm1(output_imag_18_1),   .input_b_imag3_vmm1(output_imag_19_1),   .input_b_imag4_vmm1(output_imag_20_1),  
.input_b_real5_vmm1(output_real_21_1), .input_b_real6_vmm1(output_real_22_1), .input_b_real7_vmm1(output_real_23_1), .input_b_real8_vmm1(output_real_24_1),
.input_b_imag5_vmm1(output_imag_21_1),   .input_b_imag6_vmm1(output_imag_22_1),   .input_b_imag7_vmm1(output_imag_23_1),   .input_b_imag8_vmm1(output_imag_24_1),  
.input_b_real9_vmm1(output_real_25_1), .input_b_real10_vmm1(output_real_26_1), .input_b_real11_vmm1(output_real_27_1), .input_b_real12_vmm1(output_real_28_1),
.input_b_imag9_vmm1(output_imag_25_1),   .input_b_imag10_vmm1(output_imag_26_1),   .input_b_imag11_vmm1(output_imag_27_1),   .input_b_imag12_vmm1(output_imag_28_1),  
.input_b_real13_vmm1(output_real_29_1), .input_b_real14_vmm1(output_real_30_1), .input_b_real15_vmm1(output_real_31_1), .input_b_real16_vmm1(output_real_32_1),
.input_b_imag13_vmm1(output_imag_29_1),   .input_b_imag14_vmm1(output_imag_30_1),   .input_b_imag15_vmm1(output_imag_31_1),   .input_b_imag16_vmm1(output_imag_32_1),  
.input_b_real1_vmm2(output_real_33_1), .input_b_real2_vmm2(output_real_34_1), .input_b_real3_vmm2(output_real_35_1), .input_b_real4_vmm2(output_real_36_1),
.input_b_imag1_vmm2(output_imag_33_1),   .input_b_imag2_vmm2(output_imag_34_1),   .input_b_imag3_vmm2(output_imag_35_1),   .input_b_imag4_vmm2(output_imag_36_1),  
.input_b_real5_vmm2(output_real_37_1), .input_b_real6_vmm2(output_real_38_1), .input_b_real7_vmm2(output_real_39_1), .input_b_real8_vmm2(output_real_40_1),
.input_b_imag5_vmm2(output_imag_37_1),   .input_b_imag6_vmm2(output_imag_38_1),   .input_b_imag7_vmm2(output_imag_39_1),   .input_b_imag8_vmm2(output_imag_40_1),  
.input_b_real9_vmm2(output_real_41_1), .input_b_real10_vmm2(output_real_42_1), .input_b_real11_vmm2(output_real_43_1), .input_b_real12_vmm2(output_real_44_1),
.input_b_imag9_vmm2(output_imag_41_1),   .input_b_imag10_vmm2(output_imag_42_1),   .input_b_imag11_vmm2(output_imag_43_1),   .input_b_imag12_vmm2(output_imag_44_1),  
.input_b_real13_vmm2(output_real_45_1), .input_b_real14_vmm2(output_real_46_1), .input_b_real15_vmm2(output_real_47_1), .input_b_real16_vmm2(output_real_48_1),
.input_b_imag13_vmm2(output_imag_45_1),   .input_b_imag14_vmm2(output_imag_46_1),   .input_b_imag15_vmm2(output_imag_47_1),   .input_b_imag16_vmm2(output_imag_48_1),  
.input_b_real1_vmm3(output_real_49_1), .input_b_real2_vmm3(output_real_50_1), .input_b_real3_vmm3(output_real_51_1), .input_b_real4_vmm3(output_real_52_1),
.input_b_imag1_vmm3(output_imag_49_1),   .input_b_imag2_vmm3(output_imag_50_1),   .input_b_imag3_vmm3(output_imag_51_1),   .input_b_imag4_vmm3(output_imag_52_1),  
.input_b_real5_vmm3(output_real_53_1), .input_b_real6_vmm3(output_real_54_1), .input_b_real7_vmm3(output_real_55_1), .input_b_real8_vmm3(output_real_56_1),
.input_b_imag5_vmm3(output_imag_53_1),   .input_b_imag6_vmm3(output_imag_54_1),   .input_b_imag7_vmm3(output_imag_55_1),   .input_b_imag8_vmm3(output_imag_56_1),  
.input_b_real9_vmm3(output_real_57_1), .input_b_real10_vmm3(output_real_58_1), .input_b_real11_vmm3(output_real_59_1), .input_b_real12_vmm3(output_real_60_1),
.input_b_imag9_vmm3(output_imag_57_1),   .input_b_imag10_vmm3(output_imag_58_1),   .input_b_imag11_vmm3(output_imag_59_1),   .input_b_imag12_vmm3(output_imag_60_1),  
.input_b_real13_vmm3(output_real_61_1), .input_b_real14_vmm3(output_real_62_1), .input_b_real15_vmm3(output_real_63_1), .input_b_real16_vmm3(output_real_64_1),
.input_b_imag13_vmm3(output_imag_61_1),   .input_b_imag14_vmm3(output_imag_62_1),   .input_b_imag15_vmm3(output_imag_63_1),   .input_b_imag16_vmm3(output_imag_64_1),
.output_z_real(output_z_real1_1),
.output_z_imag(output_z_imag1_1)
);

vmm_adder DUT_VMM_ADDER2(
.CLK(CLK),               
.rst(rst), 
.input_a_real1_vmm0(output_data_divider1[31:16]), .input_a_real2_vmm0(output_data_divider2[31:16]), .input_a_real3_vmm0(output_data_divider3[31:16]), .input_a_real4_vmm0(output_data_divider4[31:16]),
.input_a_imag1_vmm0(output_data_divider1[15:0]),  .input_a_imag2_vmm0(output_data_divider2[15:0]),  .input_a_imag3_vmm0(output_data_divider3[15:0]),  .input_a_imag4_vmm0(output_data_divider4[15:0]),  
.input_a_real5_vmm0(output_data_divider5[31:16]), .input_a_real6_vmm0(output_data_divider6[31:16]), .input_a_real7_vmm0(output_data_divider7[31:16]), .input_a_real8_vmm0(output_data_divider8[31:16]),
.input_a_imag5_vmm0(output_data_divider5[15:0]),  .input_a_imag6_vmm0(output_data_divider6[15:0]),  .input_a_imag7_vmm0(output_data_divider7[15:0]),  .input_a_imag8_vmm0(output_data_divider8[15:0]),  
.input_a_real9_vmm0(output_data_divider9[31:16]), .input_a_real10_vmm0(output_data_divider10[31:16]), .input_a_real11_vmm0(output_data_divider11[31:16]), .input_a_real12_vmm0(output_data_divider12[31:16]),
.input_a_imag9_vmm0(output_data_divider9[15:0]),  .input_a_imag10_vmm0(output_data_divider10[15:0]),  .input_a_imag11_vmm0(output_data_divider11[15:0]),  .input_a_imag12_vmm0(output_data_divider12[15:0]),  
.input_a_real13_vmm0(output_data_divider13[31:16]), .input_a_real14_vmm0(output_data_divider14[31:16]), .input_a_real15_vmm0(output_data_divider15[31:16]), .input_a_real16_vmm0(output_data_divider16[31:16]),
.input_a_imag13_vmm0(output_data_divider13[15:0]),  .input_a_imag14_vmm0(output_data_divider14[15:0]),  .input_a_imag15_vmm0(output_data_divider15[15:0]),  .input_a_imag16_vmm0(output_data_divider16[15:0]),  
.input_a_real1_vmm1(output_data_divider17[31:16]), .input_a_real2_vmm1(output_data_divider18[31:16]), .input_a_real3_vmm1(output_data_divider19[31:16]), .input_a_real4_vmm1(output_data_divider20[31:16]),
.input_a_imag1_vmm1(output_data_divider17[15:0]),  .input_a_imag2_vmm1(output_data_divider18[15:0]),  .input_a_imag3_vmm1(output_data_divider19[15:0]),  .input_a_imag4_vmm1(output_data_divider20[15:0]),  
.input_a_real5_vmm1(output_data_divider21[31:16]), .input_a_real6_vmm1(output_data_divider22[31:16]), .input_a_real7_vmm1(output_data_divider23[31:16]), .input_a_real8_vmm1(output_data_divider24[31:16]),
.input_a_imag5_vmm1(output_data_divider21[15:0]),  .input_a_imag6_vmm1(output_data_divider22[15:0]),  .input_a_imag7_vmm1(output_data_divider23[15:0]),  .input_a_imag8_vmm1(output_data_divider24[15:0]),  
.input_a_real9_vmm1(output_data_divider25[31:16]), .input_a_real10_vmm1(output_data_divider26[31:16]), .input_a_real11_vmm1(output_data_divider27[31:16]), .input_a_real12_vmm1(output_data_divider28[31:16]),
.input_a_imag9_vmm1(output_data_divider25[15:0]),  .input_a_imag10_vmm1(output_data_divider26[15:0]),  .input_a_imag11_vmm1(output_data_divider27[15:0]),  .input_a_imag12_vmm1(output_data_divider28[15:0]),  
.input_a_real13_vmm1(output_data_divider29[31:16]), .input_a_real14_vmm1(output_data_divider30[31:16]), .input_a_real15_vmm1(output_data_divider31[31:16]), .input_a_real16_vmm1(output_data_divider32[31:16]),
.input_a_imag13_vmm1(output_data_divider29[15:0]),  .input_a_imag14_vmm1(output_data_divider30[15:0]),  .input_a_imag15_vmm1(output_data_divider31[15:0]),  .input_a_imag16_vmm1(output_data_divider32[15:0]),  
.input_a_real1_vmm2(output_data_divider33[31:16]), .input_a_real2_vmm2(output_data_divider34[31:16]), .input_a_real3_vmm2(output_data_divider35[31:16]), .input_a_real4_vmm2(output_data_divider36[31:16]),
.input_a_imag1_vmm2(output_data_divider33[15:0]),  .input_a_imag2_vmm2(output_data_divider34[15:0]),  .input_a_imag3_vmm2(output_data_divider35[15:0]),  .input_a_imag4_vmm2(output_data_divider36[15:0]),  
.input_a_real5_vmm2(output_data_divider37[31:16]), .input_a_real6_vmm2(output_data_divider38[31:16]), .input_a_real7_vmm2(output_data_divider39[31:16]), .input_a_real8_vmm2(output_data_divider40[31:16]),
.input_a_imag5_vmm2(output_data_divider37[15:0]),  .input_a_imag6_vmm2(output_data_divider38[15:0]),  .input_a_imag7_vmm2(output_data_divider39[15:0]),  .input_a_imag8_vmm2(output_data_divider40[15:0]),  
.input_a_real9_vmm2(output_data_divider41[31:16]), .input_a_real10_vmm2(output_data_divider42[31:16]), .input_a_real11_vmm2(output_data_divider43[31:16]), .input_a_real12_vmm2(output_data_divider44[31:16]),
.input_a_imag9_vmm2(output_data_divider41[15:0]),  .input_a_imag10_vmm2(output_data_divider42[15:0]),  .input_a_imag11_vmm2(output_data_divider43[15:0]),  .input_a_imag12_vmm2(output_data_divider44[15:0]),  
.input_a_real13_vmm2(output_data_divider45[31:16]), .input_a_real14_vmm2(output_data_divider46[31:16]), .input_a_real15_vmm2(output_data_divider47[31:16]), .input_a_real16_vmm2(output_data_divider48[31:16]),
.input_a_imag13_vmm2(output_data_divider45[15:0]),  .input_a_imag14_vmm2(output_data_divider46[15:0]),  .input_a_imag15_vmm2(output_data_divider47[15:0]),  .input_a_imag16_vmm2(output_data_divider48[15:0]),  
.input_a_real1_vmm3(output_data_divider49[31:16]), .input_a_real2_vmm3(output_data_divider50[31:16]), .input_a_real3_vmm3(output_data_divider51[31:16]), .input_a_real4_vmm3(output_data_divider52[31:16]),
.input_a_imag1_vmm3(output_data_divider49[15:0]),  .input_a_imag2_vmm3(output_data_divider50[15:0]),  .input_a_imag3_vmm3(output_data_divider51[15:0]),  .input_a_imag4_vmm3(output_data_divider52[15:0]),  
.input_a_real5_vmm3(output_data_divider53[31:16]), .input_a_real6_vmm3(output_data_divider54[31:16]), .input_a_real7_vmm3(output_data_divider55[31:16]), .input_a_real8_vmm3(output_data_divider56[31:16]),
.input_a_imag5_vmm3(output_data_divider53[15:0]),  .input_a_imag6_vmm3(output_data_divider54[15:0]),  .input_a_imag7_vmm3(output_data_divider55[15:0]),  .input_a_imag8_vmm3(output_data_divider56[15:0]),  
.input_a_real9_vmm3(output_data_divider57[31:16]), .input_a_real10_vmm3(output_data_divider58[31:16]), .input_a_real11_vmm3(output_data_divider59[31:16]), .input_a_real12_vmm3(output_data_divider60[31:16]),
.input_a_imag9_vmm3(output_data_divider57[15:0]),  .input_a_imag10_vmm3(output_data_divider58[15:0]),  .input_a_imag11_vmm3(output_data_divider59[15:0]),  .input_a_imag12_vmm3(output_data_divider60[15:0]),  
.input_a_real13_vmm3(output_data_divider61[31:16]), .input_a_real14_vmm3(output_data_divider62[31:16]), .input_a_real15_vmm3(output_data_divider63[31:16]), .input_a_real16_vmm3(output_data_divider64[31:16]),
.input_a_imag13_vmm3(output_data_divider61[15:0]),  .input_a_imag14_vmm3(output_data_divider62[15:0]),  .input_a_imag15_vmm3(output_data_divider63[15:0]),  .input_a_imag16_vmm3(output_data_divider64[15:0]),  
.input_b_real1_vmm0(output_real_1_2), .input_b_real2_vmm0(output_real_2_2), .input_b_real3_vmm0(output_real_3_2), .input_b_real4_vmm0(output_real_4_2),
.input_b_imag1_vmm0(output_imag_1_2),   .input_b_imag2_vmm0(output_imag_2_2),   .input_b_imag3_vmm0(output_imag_3_2),   .input_b_imag4_vmm0(output_imag_4_2),  
.input_b_real5_vmm0(output_real_5_2), .input_b_real6_vmm0(output_real_6_2), .input_b_real7_vmm0(output_real_7_2), .input_b_real8_vmm0(output_real_8_2),
.input_b_imag5_vmm0(output_imag_5_2),   .input_b_imag6_vmm0(output_imag_6_2),   .input_b_imag7_vmm0(output_imag_7_2),   .input_b_imag8_vmm0(output_imag_8_2),  
.input_b_real9_vmm0(output_real_9_2), .input_b_real10_vmm0(output_real_10_2), .input_b_real11_vmm0(output_real_11_2), .input_b_real12_vmm0(output_real_12_2),
.input_b_imag9_vmm0(output_imag_9_2),   .input_b_imag10_vmm0(output_imag_10_2),   .input_b_imag11_vmm0(output_imag_11_2),   .input_b_imag12_vmm0(output_imag_12_2),  
.input_b_real13_vmm0(output_real_13_2), .input_b_real14_vmm0(output_real_14_2), .input_b_real15_vmm0(output_real_15_2), .input_b_real16_vmm0(output_real_16_2),
.input_b_imag13_vmm0(output_imag_13_2),   .input_b_imag14_vmm0(output_imag_14_2),   .input_b_imag15_vmm0(output_imag_15_2),   .input_b_imag16_vmm0(output_imag_16_2),  
.input_b_real1_vmm1(output_real_17_2), .input_b_real2_vmm1(output_real_18_2), .input_b_real3_vmm1(output_real_19_2), .input_b_real4_vmm1(output_real_20_2),
.input_b_imag1_vmm1(output_imag_17_2),   .input_b_imag2_vmm1(output_imag_18_2),   .input_b_imag3_vmm1(output_imag_19_2),   .input_b_imag4_vmm1(output_imag_20_2),  
.input_b_real5_vmm1(output_real_21_2), .input_b_real6_vmm1(output_real_22_2), .input_b_real7_vmm1(output_real_23_2), .input_b_real8_vmm1(output_real_24_2),
.input_b_imag5_vmm1(output_imag_21_2),   .input_b_imag6_vmm1(output_imag_22_2),   .input_b_imag7_vmm1(output_imag_23_2),   .input_b_imag8_vmm1(output_imag_24_2),  
.input_b_real9_vmm1(output_real_25_2), .input_b_real10_vmm1(output_real_26_2), .input_b_real11_vmm1(output_real_27_2), .input_b_real12_vmm1(output_real_28_2),
.input_b_imag9_vmm1(output_imag_25_2),   .input_b_imag10_vmm1(output_imag_26_2),   .input_b_imag11_vmm1(output_imag_27_2),   .input_b_imag12_vmm1(output_imag_28_2),  
.input_b_real13_vmm1(output_real_29_2), .input_b_real14_vmm1(output_real_30_2), .input_b_real15_vmm1(output_real_31_2), .input_b_real16_vmm1(output_real_32_2),
.input_b_imag13_vmm1(output_imag_29_2),   .input_b_imag14_vmm1(output_imag_30_2),   .input_b_imag15_vmm1(output_imag_31_2),   .input_b_imag16_vmm1(output_imag_32_2),  
.input_b_real1_vmm2(output_real_33_2), .input_b_real2_vmm2(output_real_34_2), .input_b_real3_vmm2(output_real_35_2), .input_b_real4_vmm2(output_real_36_2),
.input_b_imag1_vmm2(output_imag_33_2),   .input_b_imag2_vmm2(output_imag_34_2),   .input_b_imag3_vmm2(output_imag_35_2),   .input_b_imag4_vmm2(output_imag_36_2),  
.input_b_real5_vmm2(output_real_37_2), .input_b_real6_vmm2(output_real_38_2), .input_b_real7_vmm2(output_real_39_2), .input_b_real8_vmm2(output_real_40_2),
.input_b_imag5_vmm2(output_imag_37_2),   .input_b_imag6_vmm2(output_imag_38_2),   .input_b_imag7_vmm2(output_imag_39_2),   .input_b_imag8_vmm2(output_imag_40_2),  
.input_b_real9_vmm2(output_real_41_2), .input_b_real10_vmm2(output_real_42_2), .input_b_real11_vmm2(output_real_43_2), .input_b_real12_vmm2(output_real_44_2),
.input_b_imag9_vmm2(output_imag_41_2),   .input_b_imag10_vmm2(output_imag_42_2),   .input_b_imag11_vmm2(output_imag_43_2),   .input_b_imag12_vmm2(output_imag_44_2),  
.input_b_real13_vmm2(output_real_45_2), .input_b_real14_vmm2(output_real_46_2), .input_b_real15_vmm2(output_real_47_2), .input_b_real16_vmm2(output_real_48_2),
.input_b_imag13_vmm2(output_imag_45_2),   .input_b_imag14_vmm2(output_imag_46_2),   .input_b_imag15_vmm2(output_imag_47_2),   .input_b_imag16_vmm2(output_imag_48_2),  
.input_b_real1_vmm3(output_real_49_2), .input_b_real2_vmm3(output_real_50_2), .input_b_real3_vmm3(output_real_51_2), .input_b_real4_vmm3(output_real_52_2),
.input_b_imag1_vmm3(output_imag_49_2),   .input_b_imag2_vmm3(output_imag_50_2),   .input_b_imag3_vmm3(output_imag_51_2),   .input_b_imag4_vmm3(output_imag_52_2),  
.input_b_real5_vmm3(output_real_53_2), .input_b_real6_vmm3(output_real_54_2), .input_b_real7_vmm3(output_real_55_2), .input_b_real8_vmm3(output_real_56_2),
.input_b_imag5_vmm3(output_imag_53_2),   .input_b_imag6_vmm3(output_imag_54_2),   .input_b_imag7_vmm3(output_imag_55_2),   .input_b_imag8_vmm3(output_imag_56_2),  
.input_b_real9_vmm3(output_real_57_2), .input_b_real10_vmm3(output_real_58_2), .input_b_real11_vmm3(output_real_59_2), .input_b_real12_vmm3(output_real_60_2),
.input_b_imag9_vmm3(output_imag_57_2),   .input_b_imag10_vmm3(output_imag_58_2),   .input_b_imag11_vmm3(output_imag_59_2),   .input_b_imag12_vmm3(output_imag_60_2),  
.input_b_real13_vmm3(output_real_61_2), .input_b_real14_vmm3(output_real_62_2), .input_b_real15_vmm3(output_real_63_2), .input_b_real16_vmm3(output_real_64_2),
.input_b_imag13_vmm3(output_imag_61_2),   .input_b_imag14_vmm3(output_imag_62_2),   .input_b_imag15_vmm3(output_imag_63_2),   .input_b_imag16_vmm3(output_imag_64_2), 
.output_z_real(output_z_real1_2),
.output_z_imag(output_z_imag1_2)
);

vmm_adder DUT_VMM_ADDER3(
.CLK(CLK),               
.rst(rst), 
.input_a_real1_vmm0(output_data_divider1[31:16]), .input_a_real2_vmm0(output_data_divider2[31:16]), .input_a_real3_vmm0(output_data_divider3[31:16]), .input_a_real4_vmm0(output_data_divider4[31:16]),
.input_a_imag1_vmm0(output_data_divider1[15:0]),  .input_a_imag2_vmm0(output_data_divider2[15:0]),  .input_a_imag3_vmm0(output_data_divider3[15:0]),  .input_a_imag4_vmm0(output_data_divider4[15:0]),  
.input_a_real5_vmm0(output_data_divider5[31:16]), .input_a_real6_vmm0(output_data_divider6[31:16]), .input_a_real7_vmm0(output_data_divider7[31:16]), .input_a_real8_vmm0(output_data_divider8[31:16]),
.input_a_imag5_vmm0(output_data_divider5[15:0]),  .input_a_imag6_vmm0(output_data_divider6[15:0]),  .input_a_imag7_vmm0(output_data_divider7[15:0]),  .input_a_imag8_vmm0(output_data_divider8[15:0]),  
.input_a_real9_vmm0(output_data_divider9[31:16]), .input_a_real10_vmm0(output_data_divider10[31:16]), .input_a_real11_vmm0(output_data_divider11[31:16]), .input_a_real12_vmm0(output_data_divider12[31:16]),
.input_a_imag9_vmm0(output_data_divider9[15:0]),  .input_a_imag10_vmm0(output_data_divider10[15:0]),  .input_a_imag11_vmm0(output_data_divider11[15:0]),  .input_a_imag12_vmm0(output_data_divider12[15:0]),  
.input_a_real13_vmm0(output_data_divider13[31:16]), .input_a_real14_vmm0(output_data_divider14[31:16]), .input_a_real15_vmm0(output_data_divider15[31:16]), .input_a_real16_vmm0(output_data_divider16[31:16]),
.input_a_imag13_vmm0(output_data_divider13[15:0]),  .input_a_imag14_vmm0(output_data_divider14[15:0]),  .input_a_imag15_vmm0(output_data_divider15[15:0]),  .input_a_imag16_vmm0(output_data_divider16[15:0]),  
.input_a_real1_vmm1(output_data_divider17[31:16]), .input_a_real2_vmm1(output_data_divider18[31:16]), .input_a_real3_vmm1(output_data_divider19[31:16]), .input_a_real4_vmm1(output_data_divider20[31:16]),
.input_a_imag1_vmm1(output_data_divider17[15:0]),  .input_a_imag2_vmm1(output_data_divider18[15:0]),  .input_a_imag3_vmm1(output_data_divider19[15:0]),  .input_a_imag4_vmm1(output_data_divider20[15:0]),  
.input_a_real5_vmm1(output_data_divider21[31:16]), .input_a_real6_vmm1(output_data_divider22[31:16]), .input_a_real7_vmm1(output_data_divider23[31:16]), .input_a_real8_vmm1(output_data_divider24[31:16]),
.input_a_imag5_vmm1(output_data_divider21[15:0]),  .input_a_imag6_vmm1(output_data_divider22[15:0]),  .input_a_imag7_vmm1(output_data_divider23[15:0]),  .input_a_imag8_vmm1(output_data_divider24[15:0]),  
.input_a_real9_vmm1(output_data_divider25[31:16]), .input_a_real10_vmm1(output_data_divider26[31:16]), .input_a_real11_vmm1(output_data_divider27[31:16]), .input_a_real12_vmm1(output_data_divider28[31:16]),
.input_a_imag9_vmm1(output_data_divider25[15:0]),  .input_a_imag10_vmm1(output_data_divider26[15:0]),  .input_a_imag11_vmm1(output_data_divider27[15:0]),  .input_a_imag12_vmm1(output_data_divider28[15:0]),  
.input_a_real13_vmm1(output_data_divider29[31:16]), .input_a_real14_vmm1(output_data_divider30[31:16]), .input_a_real15_vmm1(output_data_divider31[31:16]), .input_a_real16_vmm1(output_data_divider32[31:16]),
.input_a_imag13_vmm1(output_data_divider29[15:0]),  .input_a_imag14_vmm1(output_data_divider30[15:0]),  .input_a_imag15_vmm1(output_data_divider31[15:0]),  .input_a_imag16_vmm1(output_data_divider32[15:0]),  
.input_a_real1_vmm2(output_data_divider33[31:16]), .input_a_real2_vmm2(output_data_divider34[31:16]), .input_a_real3_vmm2(output_data_divider35[31:16]), .input_a_real4_vmm2(output_data_divider36[31:16]),
.input_a_imag1_vmm2(output_data_divider33[15:0]),  .input_a_imag2_vmm2(output_data_divider34[15:0]),  .input_a_imag3_vmm2(output_data_divider35[15:0]),  .input_a_imag4_vmm2(output_data_divider36[15:0]),  
.input_a_real5_vmm2(output_data_divider37[31:16]), .input_a_real6_vmm2(output_data_divider38[31:16]), .input_a_real7_vmm2(output_data_divider39[31:16]), .input_a_real8_vmm2(output_data_divider40[31:16]),
.input_a_imag5_vmm2(output_data_divider37[15:0]),  .input_a_imag6_vmm2(output_data_divider38[15:0]),  .input_a_imag7_vmm2(output_data_divider39[15:0]),  .input_a_imag8_vmm2(output_data_divider40[15:0]),  
.input_a_real9_vmm2(output_data_divider41[31:16]), .input_a_real10_vmm2(output_data_divider42[31:16]), .input_a_real11_vmm2(output_data_divider43[31:16]), .input_a_real12_vmm2(output_data_divider44[31:16]),
.input_a_imag9_vmm2(output_data_divider41[15:0]),  .input_a_imag10_vmm2(output_data_divider42[15:0]),  .input_a_imag11_vmm2(output_data_divider43[15:0]),  .input_a_imag12_vmm2(output_data_divider44[15:0]),  
.input_a_real13_vmm2(output_data_divider45[31:16]), .input_a_real14_vmm2(output_data_divider46[31:16]), .input_a_real15_vmm2(output_data_divider47[31:16]), .input_a_real16_vmm2(output_data_divider48[31:16]),
.input_a_imag13_vmm2(output_data_divider45[15:0]),  .input_a_imag14_vmm2(output_data_divider46[15:0]),  .input_a_imag15_vmm2(output_data_divider47[15:0]),  .input_a_imag16_vmm2(output_data_divider48[15:0]),  
.input_a_real1_vmm3(output_data_divider49[31:16]), .input_a_real2_vmm3(output_data_divider50[31:16]), .input_a_real3_vmm3(output_data_divider51[31:16]), .input_a_real4_vmm3(output_data_divider52[31:16]),
.input_a_imag1_vmm3(output_data_divider49[15:0]),  .input_a_imag2_vmm3(output_data_divider50[15:0]),  .input_a_imag3_vmm3(output_data_divider51[15:0]),  .input_a_imag4_vmm3(output_data_divider52[15:0]),  
.input_a_real5_vmm3(output_data_divider53[31:16]), .input_a_real6_vmm3(output_data_divider54[31:16]), .input_a_real7_vmm3(output_data_divider55[31:16]), .input_a_real8_vmm3(output_data_divider56[31:16]),
.input_a_imag5_vmm3(output_data_divider53[15:0]),  .input_a_imag6_vmm3(output_data_divider54[15:0]),  .input_a_imag7_vmm3(output_data_divider55[15:0]),  .input_a_imag8_vmm3(output_data_divider56[15:0]),  
.input_a_real9_vmm3(output_data_divider57[31:16]), .input_a_real10_vmm3(output_data_divider58[31:16]), .input_a_real11_vmm3(output_data_divider59[31:16]), .input_a_real12_vmm3(output_data_divider60[31:16]),
.input_a_imag9_vmm3(output_data_divider57[15:0]),  .input_a_imag10_vmm3(output_data_divider58[15:0]),  .input_a_imag11_vmm3(output_data_divider59[15:0]),  .input_a_imag12_vmm3(output_data_divider60[15:0]),  
.input_a_real13_vmm3(output_data_divider61[31:16]), .input_a_real14_vmm3(output_data_divider62[31:16]), .input_a_real15_vmm3(output_data_divider63[31:16]), .input_a_real16_vmm3(output_data_divider64[31:16]),
.input_a_imag13_vmm3(output_data_divider61[15:0]),  .input_a_imag14_vmm3(output_data_divider62[15:0]),  .input_a_imag15_vmm3(output_data_divider63[15:0]),  .input_a_imag16_vmm3(output_data_divider64[15:0]),  
.input_b_real1_vmm0(output_real_1_3), .input_b_real2_vmm0(output_real_2_3), .input_b_real3_vmm0(output_real_3_3), .input_b_real4_vmm0(output_real_4_3),
.input_b_imag1_vmm0(output_imag_1_3),   .input_b_imag2_vmm0(output_imag_2_3),   .input_b_imag3_vmm0(output_imag_3_3),   .input_b_imag4_vmm0(output_imag_4_3),  
.input_b_real5_vmm0(output_real_5_3), .input_b_real6_vmm0(output_real_6_3), .input_b_real7_vmm0(output_real_7_3), .input_b_real8_vmm0(output_real_8_3),
.input_b_imag5_vmm0(output_imag_5_3),   .input_b_imag6_vmm0(output_imag_6_3),   .input_b_imag7_vmm0(output_imag_7_3),   .input_b_imag8_vmm0(output_imag_8_3),  
.input_b_real9_vmm0(output_real_9_3), .input_b_real10_vmm0(output_real_10_3), .input_b_real11_vmm0(output_real_11_3), .input_b_real12_vmm0(output_real_12_3),
.input_b_imag9_vmm0(output_imag_9_3),   .input_b_imag10_vmm0(output_imag_10_3),   .input_b_imag11_vmm0(output_imag_11_3),   .input_b_imag12_vmm0(output_imag_12_3),  
.input_b_real13_vmm0(output_real_13_3), .input_b_real14_vmm0(output_real_14_3), .input_b_real15_vmm0(output_real_15_3), .input_b_real16_vmm0(output_real_16_3),
.input_b_imag13_vmm0(output_imag_13_3),   .input_b_imag14_vmm0(output_imag_14_3),   .input_b_imag15_vmm0(output_imag_15_3),   .input_b_imag16_vmm0(output_imag_16_3),  
.input_b_real1_vmm1(output_real_17_3), .input_b_real2_vmm1(output_real_18_3), .input_b_real3_vmm1(output_real_19_3), .input_b_real4_vmm1(output_real_20_3),
.input_b_imag1_vmm1(output_imag_17_3),   .input_b_imag2_vmm1(output_imag_18_3),   .input_b_imag3_vmm1(output_imag_19_3),   .input_b_imag4_vmm1(output_imag_20_3),  
.input_b_real5_vmm1(output_real_21_3), .input_b_real6_vmm1(output_real_22_3), .input_b_real7_vmm1(output_real_23_3), .input_b_real8_vmm1(output_real_24_3),
.input_b_imag5_vmm1(output_imag_21_3),   .input_b_imag6_vmm1(output_imag_22_3),   .input_b_imag7_vmm1(output_imag_23_3),   .input_b_imag8_vmm1(output_imag_24_3),  
.input_b_real9_vmm1(output_real_25_3), .input_b_real10_vmm1(output_real_26_3), .input_b_real11_vmm1(output_real_27_3), .input_b_real12_vmm1(output_real_28_3),
.input_b_imag9_vmm1(output_imag_25_3),   .input_b_imag10_vmm1(output_imag_26_3),   .input_b_imag11_vmm1(output_imag_27_3),   .input_b_imag12_vmm1(output_imag_28_3),  
.input_b_real13_vmm1(output_real_29_3), .input_b_real14_vmm1(output_real_30_3), .input_b_real15_vmm1(output_real_31_3), .input_b_real16_vmm1(output_real_32_3),
.input_b_imag13_vmm1(output_imag_29_3),   .input_b_imag14_vmm1(output_imag_30_3),   .input_b_imag15_vmm1(output_imag_31_3),   .input_b_imag16_vmm1(output_imag_32_3),  
.input_b_real1_vmm2(output_real_33_3), .input_b_real2_vmm2(output_real_34_3), .input_b_real3_vmm2(output_real_35_3), .input_b_real4_vmm2(output_real_36_3),
.input_b_imag1_vmm2(output_imag_33_3),   .input_b_imag2_vmm2(output_imag_34_3),   .input_b_imag3_vmm2(output_imag_35_3),   .input_b_imag4_vmm2(output_imag_36_3),  
.input_b_real5_vmm2(output_real_37_3), .input_b_real6_vmm2(output_real_38_3), .input_b_real7_vmm2(output_real_39_3), .input_b_real8_vmm2(output_real_40_3),
.input_b_imag5_vmm2(output_imag_37_3),   .input_b_imag6_vmm2(output_imag_38_3),   .input_b_imag7_vmm2(output_imag_39_3),   .input_b_imag8_vmm2(output_imag_40_3),  
.input_b_real9_vmm2(output_real_41_3), .input_b_real10_vmm2(output_real_42_3), .input_b_real11_vmm2(output_real_43_3), .input_b_real12_vmm2(output_real_44_3),
.input_b_imag9_vmm2(output_imag_41_3),   .input_b_imag10_vmm2(output_imag_42_3),   .input_b_imag11_vmm2(output_imag_43_3),   .input_b_imag12_vmm2(output_imag_44_3),  
.input_b_real13_vmm2(output_real_45_3), .input_b_real14_vmm2(output_real_46_3), .input_b_real15_vmm2(output_real_47_3), .input_b_real16_vmm2(output_real_48_3),
.input_b_imag13_vmm2(output_imag_45_3),   .input_b_imag14_vmm2(output_imag_46_3),   .input_b_imag15_vmm2(output_imag_47_3),   .input_b_imag16_vmm2(output_imag_48_3),  
.input_b_real1_vmm3(output_real_49_3), .input_b_real2_vmm3(output_real_50_3), .input_b_real3_vmm3(output_real_51_3), .input_b_real4_vmm3(output_real_52_3),
.input_b_imag1_vmm3(output_imag_49_3),   .input_b_imag2_vmm3(output_imag_50_3),   .input_b_imag3_vmm3(output_imag_51_3),   .input_b_imag4_vmm3(output_imag_52_3),  
.input_b_real5_vmm3(output_real_53_3), .input_b_real6_vmm3(output_real_54_3), .input_b_real7_vmm3(output_real_55_3), .input_b_real8_vmm3(output_real_56_3),
.input_b_imag5_vmm3(output_imag_53_3),   .input_b_imag6_vmm3(output_imag_54_3),   .input_b_imag7_vmm3(output_imag_55_3),   .input_b_imag8_vmm3(output_imag_56_3),  
.input_b_real9_vmm3(output_real_57_3), .input_b_real10_vmm3(output_real_58_3), .input_b_real11_vmm3(output_real_59_3), .input_b_real12_vmm3(output_real_60_3),
.input_b_imag9_vmm3(output_imag_57_3),   .input_b_imag10_vmm3(output_imag_58_3),   .input_b_imag11_vmm3(output_imag_59_3),   .input_b_imag12_vmm3(output_imag_60_3),  
.input_b_real13_vmm3(output_real_61_3), .input_b_real14_vmm3(output_real_62_3), .input_b_real15_vmm3(output_real_63_3), .input_b_real16_vmm3(output_real_64_3),
.input_b_imag13_vmm3(output_imag_61_3),   .input_b_imag14_vmm3(output_imag_62_3),   .input_b_imag15_vmm3(output_imag_63_3),   .input_b_imag16_vmm3(output_imag_64_3),
.output_z_real(output_z_real1_3),
.output_z_imag(output_z_imag1_3)
);

assign output_z_0 = {output_z_real1_0, output_z_imag1_0};
assign output_z_1 = {output_z_real1_1, output_z_imag1_1};
assign output_z_2 = {output_z_real1_2, output_z_imag1_2};
assign output_z_3 = {output_z_real1_3, output_z_imag1_3};
//assign output_z_3 = 16'd0;

endmodule
