
module memory_rom_59(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hb66dbe19;
    11'b00000000001: data <= 32'hb507bb2c;
    11'b00000000010: data <= 32'h32b73ac1;
    11'b00000000011: data <= 32'hb54e3f5c;
    11'b00000000100: data <= 32'hbe52396b;
    11'b00000000101: data <= 32'hbfedbcf5;
    11'b00000000110: data <= 32'hbd00bdb3;
    11'b00000000111: data <= 32'hb7f63272;
    11'b00000001000: data <= 32'hb0d73d5b;
    11'b00000001001: data <= 32'h38243a61;
    11'b00000001010: data <= 32'h3e0f2c31;
    11'b00000001011: data <= 32'h3dff39b6;
    11'b00000001100: data <= 32'ha8153f8d;
    11'b00000001101: data <= 32'hbd5e3ee5;
    11'b00000001110: data <= 32'hb92532a6;
    11'b00000001111: data <= 32'h3cbfbc17;
    11'b00000010000: data <= 32'h3f06bcde;
    11'b00000010001: data <= 32'h3927bc9a;
    11'b00000010010: data <= 32'haf79bce4;
    11'b00000010011: data <= 32'h397eb9a6;
    11'b00000010100: data <= 32'h3e303818;
    11'b00000010101: data <= 32'h38fd3c06;
    11'b00000010110: data <= 32'hbd97b106;
    11'b00000010111: data <= 32'hc0abbe6f;
    11'b00000011000: data <= 32'hbe6dbda8;
    11'b00000011001: data <= 32'hb8d32676;
    11'b00000011010: data <= 32'hb3e93880;
    11'b00000011011: data <= 32'h27edb557;
    11'b00000011100: data <= 32'h38a9b9ac;
    11'b00000011101: data <= 32'h385c3a44;
    11'b00000011110: data <= 32'hb81e413c;
    11'b00000011111: data <= 32'hbd404106;
    11'b00000100000: data <= 32'hb8ab3950;
    11'b00000100001: data <= 32'h3a50b9f7;
    11'b00000100010: data <= 32'h3bd7b9ab;
    11'b00000100011: data <= 32'h2fdeb473;
    11'b00000100100: data <= 32'h31c0b569;
    11'b00000100101: data <= 32'h3edfb4ce;
    11'b00000100110: data <= 32'h415d3532;
    11'b00000100111: data <= 32'h3d4a3915;
    11'b00000101000: data <= 32'hbc60b221;
    11'b00000101001: data <= 32'hbff4bcf7;
    11'b00000101010: data <= 32'hbbc4bc9f;
    11'b00000101011: data <= 32'h2b9db68d;
    11'b00000101100: data <= 32'haa0eb8d1;
    11'b00000101101: data <= 32'hb66ebe8e;
    11'b00000101110: data <= 32'haf9cbe07;
    11'b00000101111: data <= 32'h2fb838bf;
    11'b00000110000: data <= 32'hb7de4133;
    11'b00000110001: data <= 32'hbcf6408b;
    11'b00000110010: data <= 32'hbc1f3537;
    11'b00000110011: data <= 32'hb4fdb9a5;
    11'b00000110100: data <= 32'hb474a99f;
    11'b00000110101: data <= 32'hb8e13996;
    11'b00000110110: data <= 32'h326f35e8;
    11'b00000110111: data <= 32'h4036affc;
    11'b00000111000: data <= 32'h41d73494;
    11'b00000111001: data <= 32'h3d693b8e;
    11'b00000111010: data <= 32'hbadf396a;
    11'b00000111011: data <= 32'hbcd9b2ca;
    11'b00000111100: data <= 32'h305cb906;
    11'b00000111101: data <= 32'h3b38b988;
    11'b00000111110: data <= 32'h314abd81;
    11'b00000111111: data <= 32'hb89fc0a6;
    11'b00001000000: data <= 32'hae60bf78;
    11'b00001000001: data <= 32'h391b3420;
    11'b00001000010: data <= 32'h32e03f8d;
    11'b00001000011: data <= 32'hbbd23cfa;
    11'b00001000100: data <= 32'hbe3fb79e;
    11'b00001000101: data <= 32'hbd7eba97;
    11'b00001000110: data <= 32'hbd143629;
    11'b00001000111: data <= 32'hbcae3c4b;
    11'b00001001000: data <= 32'haf013439;
    11'b00001001001: data <= 32'h3e81b816;
    11'b00001001010: data <= 32'h405b3389;
    11'b00001001011: data <= 32'h3a203e84;
    11'b00001001100: data <= 32'hba5e3f88;
    11'b00001001101: data <= 32'hb8163b31;
    11'b00001001110: data <= 32'h3b43aa53;
    11'b00001001111: data <= 32'h3cc9b864;
    11'b00001010000: data <= 32'h281fbcfe;
    11'b00001010001: data <= 32'hb86dbffb;
    11'b00001010010: data <= 32'h388abe71;
    11'b00001010011: data <= 32'h3f40a580;
    11'b00001010100: data <= 32'h3d183bd9;
    11'b00001010101: data <= 32'hb8593221;
    11'b00001010110: data <= 32'hbed8bc40;
    11'b00001010111: data <= 32'hbea8baad;
    11'b00001011000: data <= 32'hbd883711;
    11'b00001011001: data <= 32'hbd0138ff;
    11'b00001011010: data <= 32'hb88cb98d;
    11'b00001011011: data <= 32'h3913bd8d;
    11'b00001011100: data <= 32'h3c202705;
    11'b00001011101: data <= 32'h2c75403d;
    11'b00001011110: data <= 32'hba7d4130;
    11'b00001011111: data <= 32'hb3ef3d96;
    11'b00001100000: data <= 32'h3a9f3452;
    11'b00001100001: data <= 32'h38d8a800;
    11'b00001100010: data <= 32'hb8a7b52d;
    11'b00001100011: data <= 32'hb860bb98;
    11'b00001100100: data <= 32'h3d53bc05;
    11'b00001100101: data <= 32'h41b8b0af;
    11'b00001100110: data <= 32'h401736f8;
    11'b00001100111: data <= 32'hb073b0cd;
    11'b00001101000: data <= 32'hbd40bb2b;
    11'b00001101001: data <= 32'hbbd3b803;
    11'b00001101010: data <= 32'hb8be34c7;
    11'b00001101011: data <= 32'hbb09b40f;
    11'b00001101100: data <= 32'hbb75bf9d;
    11'b00001101101: data <= 32'hb2dac091;
    11'b00001101110: data <= 32'h3501b511;
    11'b00001101111: data <= 32'hafe24002;
    11'b00001110000: data <= 32'hb986409a;
    11'b00001110001: data <= 32'hb6963bc1;
    11'b00001110010: data <= 32'h26d831a9;
    11'b00001110011: data <= 32'hb861388e;
    11'b00001110100: data <= 32'hbdba3a38;
    11'b00001110101: data <= 32'hb9cd2898;
    11'b00001110110: data <= 32'h3e56b8cf;
    11'b00001110111: data <= 32'h4218b27c;
    11'b00001111000: data <= 32'h400d37a6;
    11'b00001111001: data <= 32'h21043689;
    11'b00001111010: data <= 32'hb8a9228d;
    11'b00001111011: data <= 32'h339730e8;
    11'b00001111100: data <= 32'h380e3410;
    11'b00001111101: data <= 32'hb6eebadd;
    11'b00001111110: data <= 32'hbc63c114;
    11'b00001111111: data <= 32'hb709c146;
    11'b00010000000: data <= 32'h381db8f4;
    11'b00010000001: data <= 32'h37133d40;
    11'b00010000010: data <= 32'hb4d93cb6;
    11'b00010000011: data <= 32'hb96cac26;
    11'b00010000100: data <= 32'hbaadb175;
    11'b00010000101: data <= 32'hbdf73bba;
    11'b00010000110: data <= 32'hc0103d80;
    11'b00010000111: data <= 32'hbc3d33f8;
    11'b00010001000: data <= 32'h3c61ba93;
    11'b00010001001: data <= 32'h4070b5ce;
    11'b00010001010: data <= 32'h3cf33b14;
    11'b00010001011: data <= 32'hb0853d8c;
    11'b00010001100: data <= 32'h2cb83c4c;
    11'b00010001101: data <= 32'h3cd73a7e;
    11'b00010001110: data <= 32'h3c7a37a7;
    11'b00010001111: data <= 32'hb608b982;
    11'b00010010000: data <= 32'hbca2c047;
    11'b00010010001: data <= 32'haad0c06f;
    11'b00010010010: data <= 32'h3dc2b9b0;
    11'b00010010011: data <= 32'h3dc73745;
    11'b00010010100: data <= 32'h33b9abb8;
    11'b00010010101: data <= 32'hb98abbbe;
    11'b00010010110: data <= 32'hbc34b646;
    11'b00010010111: data <= 32'hbe313c54;
    11'b00010011000: data <= 32'hbffc3cce;
    11'b00010011001: data <= 32'hbd7ab70e;
    11'b00010011010: data <= 32'h30acbe83;
    11'b00010011011: data <= 32'h3b3ab997;
    11'b00010011100: data <= 32'h336a3cc7;
    11'b00010011101: data <= 32'hb6293ff8;
    11'b00010011110: data <= 32'h35f03e1f;
    11'b00010011111: data <= 32'h3d983c45;
    11'b00010100000: data <= 32'h3a813b29;
    11'b00010100001: data <= 32'hbb333290;
    11'b00010100010: data <= 32'hbd24bb88;
    11'b00010100011: data <= 32'h37fabd46;
    11'b00010100100: data <= 32'h40b4b8c7;
    11'b00010100101: data <= 32'h405eae8e;
    11'b00010100110: data <= 32'h3912b94c;
    11'b00010100111: data <= 32'hb56ebc6a;
    11'b00010101000: data <= 32'hb608b197;
    11'b00010101001: data <= 32'hb9053c46;
    11'b00010101010: data <= 32'hbd6c3877;
    11'b00010101011: data <= 32'hbdfcbdf7;
    11'b00010101100: data <= 32'hb991c100;
    11'b00010101101: data <= 32'hac3abc4f;
    11'b00010101110: data <= 32'hb4833c48;
    11'b00010101111: data <= 32'hb68f3ec3;
    11'b00010110000: data <= 32'h35323bf5;
    11'b00010110001: data <= 32'h3acb39f2;
    11'b00010110010: data <= 32'hb10c3d1b;
    11'b00010110011: data <= 32'hbeeb3d27;
    11'b00010110100: data <= 32'hbe263488;
    11'b00010110101: data <= 32'h3989b8a2;
    11'b00010110110: data <= 32'h4104b79d;
    11'b00010110111: data <= 32'h4029b110;
    11'b00010111000: data <= 32'h38c8b5e1;
    11'b00010111001: data <= 32'h326fb673;
    11'b00010111010: data <= 32'h3a8c3744;
    11'b00010111011: data <= 32'h39953c83;
    11'b00010111100: data <= 32'hb88e2b5c;
    11'b00010111101: data <= 32'hbdd2c027;
    11'b00010111110: data <= 32'hbbfac196;
    11'b00010111111: data <= 32'hb05ebcfc;
    11'b00011000000: data <= 32'h29cd383e;
    11'b00011000001: data <= 32'hac2538a6;
    11'b00011000010: data <= 32'h31d3b3fd;
    11'b00011000011: data <= 32'h302b2bd3;
    11'b00011000100: data <= 32'hbc213dcc;
    11'b00011000101: data <= 32'hc0963fc3;
    11'b00011000110: data <= 32'hbf2b3a2e;
    11'b00011000111: data <= 32'h34f5b83e;
    11'b00011001000: data <= 32'h3ec0b88a;
    11'b00011001001: data <= 32'h3c672f88;
    11'b00011001010: data <= 32'h301c36f6;
    11'b00011001011: data <= 32'h3906388d;
    11'b00011001100: data <= 32'h3f523c65;
    11'b00011001101: data <= 32'h3e5a3d4d;
    11'b00011001110: data <= 32'hb2e23141;
    11'b00011001111: data <= 32'hbdaabeb6;
    11'b00011010000: data <= 32'hb9e6c06b;
    11'b00011010001: data <= 32'h38afbc2f;
    11'b00011010010: data <= 32'h3b75aeb6;
    11'b00011010011: data <= 32'h37a6b97e;
    11'b00011010100: data <= 32'h320dbdba;
    11'b00011010101: data <= 32'hae99b7bc;
    11'b00011010110: data <= 32'hbc563dba;
    11'b00011010111: data <= 32'hc0413f88;
    11'b00011011000: data <= 32'hbf6534ee;
    11'b00011011001: data <= 32'hb6e2bcc4;
    11'b00011011010: data <= 32'h3591bb38;
    11'b00011011011: data <= 32'hb1d435e2;
    11'b00011011100: data <= 32'hb7503c0d;
    11'b00011011101: data <= 32'h3a1a3c0c;
    11'b00011011110: data <= 32'h403f3d09;
    11'b00011011111: data <= 32'h3e1d3e27;
    11'b00011100000: data <= 32'hb87b3afe;
    11'b00011100001: data <= 32'hbe20b761;
    11'b00011100010: data <= 32'hb45cbc2a;
    11'b00011100011: data <= 32'h3db9b8a5;
    11'b00011100100: data <= 32'h3e98b79b;
    11'b00011100101: data <= 32'h3a7cbd89;
    11'b00011100110: data <= 32'h3648bf55;
    11'b00011100111: data <= 32'h36b5b7ad;
    11'b00011101000: data <= 32'hb0cc3d8d;
    11'b00011101001: data <= 32'hbcf23d5f;
    11'b00011101010: data <= 32'hbe81b921;
    11'b00011101011: data <= 32'hbc47c00e;
    11'b00011101100: data <= 32'hb9abbd00;
    11'b00011101101: data <= 32'hbbdb356d;
    11'b00011101110: data <= 32'hb9e13a9c;
    11'b00011101111: data <= 32'h39493776;
    11'b00011110000: data <= 32'h3ec039b5;
    11'b00011110001: data <= 32'h39853e59;
    11'b00011110010: data <= 32'hbd583eff;
    11'b00011110011: data <= 32'hbf183abc;
    11'b00011110100: data <= 32'ha80b10b3;
    11'b00011110101: data <= 32'h3eaab161;
    11'b00011110110: data <= 32'h3e28b722;
    11'b00011110111: data <= 32'h38b5bcd4;
    11'b00011111000: data <= 32'h390fbd32;
    11'b00011111001: data <= 32'h3da52c82;
    11'b00011111010: data <= 32'h3cfc3dcc;
    11'b00011111011: data <= 32'hb0773ab0;
    11'b00011111100: data <= 32'hbd0bbd15;
    11'b00011111101: data <= 32'hbd05c0a3;
    11'b00011111110: data <= 32'hbb33bd16;
    11'b00011111111: data <= 32'hbad72b78;
    11'b00100000000: data <= 32'hb803ae03;
    11'b00100000001: data <= 32'h382dbab9;
    11'b00100000010: data <= 32'h3bf9b46f;
    11'b00100000011: data <= 32'hb2533da9;
    11'b00100000100: data <= 32'hbf9c4084;
    11'b00100000101: data <= 32'hbfaf3dcf;
    11'b00100000110: data <= 32'hb25b348e;
    11'b00100000111: data <= 32'h3c0faecd;
    11'b00100001000: data <= 32'h380bb145;
    11'b00100001001: data <= 32'hb1b2b763;
    11'b00100001010: data <= 32'h39aab58b;
    11'b00100001011: data <= 32'h408639bd;
    11'b00100001100: data <= 32'h40833e4f;
    11'b00100001101: data <= 32'h37ba3a31;
    11'b00100001110: data <= 32'hbc17bc16;
    11'b00100001111: data <= 32'hbbc4bec4;
    11'b00100010000: data <= 32'hb41aba5d;
    11'b00100010001: data <= 32'ha643b363;
    11'b00100010010: data <= 32'h2888bcc4;
    11'b00100010011: data <= 32'h37e2c049;
    11'b00100010100: data <= 32'h3920bc78;
    11'b00100010101: data <= 32'hb60b3c9f;
    11'b00100010110: data <= 32'hbed6404d;
    11'b00100010111: data <= 32'hbeee3c54;
    11'b00100011000: data <= 32'hb8e0b47d;
    11'b00100011001: data <= 32'hb0dfb6a4;
    11'b00100011010: data <= 32'hbb2d2e64;
    11'b00100011011: data <= 32'hbc53323e;
    11'b00100011100: data <= 32'h38803278;
    11'b00100011101: data <= 32'h40f73af6;
    11'b00100011110: data <= 32'h409c3e57;
    11'b00100011111: data <= 32'h34643cb9;
    11'b00100100000: data <= 32'hbc53261b;
    11'b00100100001: data <= 32'hb801b68a;
    11'b00100100010: data <= 32'h390b13df;
    11'b00100100011: data <= 32'h3a2eb4aa;
    11'b00100100100: data <= 32'h3604bf2f;
    11'b00100100101: data <= 32'h3847c155;
    11'b00100100110: data <= 32'h3b29bd2c;
    11'b00100100111: data <= 32'h363a3c11;
    11'b00100101000: data <= 32'hb9b93e6b;
    11'b00100101001: data <= 32'hbcb52fea;
    11'b00100101010: data <= 32'hbb5abcac;
    11'b00100101011: data <= 32'hbc66ba3c;
    11'b00100101100: data <= 32'hbf573217;
    11'b00100101101: data <= 32'hbe553398;
    11'b00100101110: data <= 32'h3530b1d8;
    11'b00100101111: data <= 32'h401033b5;
    11'b00100110000: data <= 32'h3df13d43;
    11'b00100110001: data <= 32'hb82b3ede;
    11'b00100110010: data <= 32'hbd5c3cd2;
    11'b00100110011: data <= 32'hb19e3a44;
    11'b00100110100: data <= 32'h3c383972;
    11'b00100110101: data <= 32'h3a83ad35;
    11'b00100110110: data <= 32'h2df9be61;
    11'b00100110111: data <= 32'h37bcc05b;
    11'b00100111000: data <= 32'h3e36ba14;
    11'b00100111001: data <= 32'h3e9d3c58;
    11'b00100111010: data <= 32'h384f3c29;
    11'b00100111011: data <= 32'hb812b947;
    11'b00100111100: data <= 32'hbb0abe68;
    11'b00100111101: data <= 32'hbd03ba1e;
    11'b00100111110: data <= 32'hbf233150;
    11'b00100111111: data <= 32'hbda4b5d7;
    11'b00101000000: data <= 32'h318fbd69;
    11'b00101000001: data <= 32'h3d35bb3f;
    11'b00101000010: data <= 32'h37a03a85;
    11'b00101000011: data <= 32'hbcde3fdb;
    11'b00101000100: data <= 32'hbde53f0e;
    11'b00101000101: data <= 32'haff23cb1;
    11'b00101000110: data <= 32'h39993ad7;
    11'b00101000111: data <= 32'had1433bf;
    11'b00101001000: data <= 32'hba90ba92;
    11'b00101001001: data <= 32'h330dbc8e;
    11'b00101001010: data <= 32'h403b1503;
    11'b00101001011: data <= 32'h41333ce2;
    11'b00101001100: data <= 32'h3d2d3a62;
    11'b00101001101: data <= 32'haea6b975;
    11'b00101001110: data <= 32'hb81dbc79;
    11'b00101001111: data <= 32'hb8b4b10c;
    11'b00101010000: data <= 32'hbb3532cf;
    11'b00101010001: data <= 32'hba44bca2;
    11'b00101010010: data <= 32'h3141c12a;
    11'b00101010011: data <= 32'h3a6abf9c;
    11'b00101010100: data <= 32'h2a383567;
    11'b00101010101: data <= 32'hbcb23eef;
    11'b00101010110: data <= 32'hbcb63d7d;
    11'b00101010111: data <= 32'hb2cf38be;
    11'b00101011000: data <= 32'hb11237da;
    11'b00101011001: data <= 32'hbd9c37c2;
    11'b00101011010: data <= 32'hbf97aab5;
    11'b00101011011: data <= 32'hb1fbb5e4;
    11'b00101011100: data <= 32'h405734fa;
    11'b00101011101: data <= 32'h413f3c9a;
    11'b00101011110: data <= 32'h3c6f3b3d;
    11'b00101011111: data <= 32'hb18e2aef;
    11'b00101100000: data <= 32'haae72d00;
    11'b00101100001: data <= 32'h362c3a97;
    11'b00101100010: data <= 32'h2db7372f;
    11'b00101100011: data <= 32'hb489be41;
    11'b00101100100: data <= 32'h3120c228;
    11'b00101100101: data <= 32'h3a4bc047;
    11'b00101100110: data <= 32'h38173117;
    11'b00101100111: data <= 32'hb4793cb2;
    11'b00101101000: data <= 32'hb700357e;
    11'b00101101001: data <= 32'hb26bb751;
    11'b00101101010: data <= 32'hbb05a6dc;
    11'b00101101011: data <= 32'hc0a038c0;
    11'b00101101100: data <= 32'hc1003336;
    11'b00101101101: data <= 32'hb828b753;
    11'b00101101110: data <= 32'h3eb5b287;
    11'b00101101111: data <= 32'h3efc39a9;
    11'b00101110000: data <= 32'h31df3c6e;
    11'b00101110001: data <= 32'hb88f3be0;
    11'b00101110010: data <= 32'h34563cf9;
    11'b00101110011: data <= 32'h3c0d3e93;
    11'b00101110100: data <= 32'h369e3a78;
    11'b00101110101: data <= 32'hb6f3bd26;
    11'b00101110110: data <= 32'ha953c116;
    11'b00101110111: data <= 32'h3c73be0e;
    11'b00101111000: data <= 32'h3e083572;
    11'b00101111001: data <= 32'h3b8e38f0;
    11'b00101111010: data <= 32'h3675b8ec;
    11'b00101111011: data <= 32'h293abca2;
    11'b00101111100: data <= 32'hbb64b117;
    11'b00101111101: data <= 32'hc0753986;
    11'b00101111110: data <= 32'hc08fab64;
    11'b00101111111: data <= 32'hb8bfbd65;
    11'b00110000000: data <= 32'h3ba3bd3f;
    11'b00110000001: data <= 32'h38af22eb;
    11'b00110000010: data <= 32'hba1f3c6d;
    11'b00110000011: data <= 32'hbae83d9e;
    11'b00110000100: data <= 32'h369c3e74;
    11'b00110000101: data <= 32'h3baa3f46;
    11'b00110000110: data <= 32'hb2423c67;
    11'b00110000111: data <= 32'hbd2eb819;
    11'b00110001000: data <= 32'hb80dbd7f;
    11'b00110001001: data <= 32'h3d92b828;
    11'b00110001010: data <= 32'h40923923;
    11'b00110001011: data <= 32'h3ec434fd;
    11'b00110001100: data <= 32'h3ae4bb56;
    11'b00110001101: data <= 32'h36debbb6;
    11'b00110001110: data <= 32'hb3ac360b;
    11'b00110001111: data <= 32'hbcf33b7a;
    11'b00110010000: data <= 32'hbdc9b865;
    11'b00110010001: data <= 32'hb6fdc0c6;
    11'b00110010010: data <= 32'h36a1c09d;
    11'b00110010011: data <= 32'hae7db886;
    11'b00110010100: data <= 32'hbc0f3a5e;
    11'b00110010101: data <= 32'hb9453bc3;
    11'b00110010110: data <= 32'h38113b95;
    11'b00110010111: data <= 32'h36973d25;
    11'b00110011000: data <= 32'hbd3c3cc4;
    11'b00110011001: data <= 32'hc0c13478;
    11'b00110011010: data <= 32'hbc39b5d8;
    11'b00110011011: data <= 32'h3d422d82;
    11'b00110011100: data <= 32'h407c3983;
    11'b00110011101: data <= 32'h3dc63417;
    11'b00110011110: data <= 32'h395db7ee;
    11'b00110011111: data <= 32'h3a1f1eef;
    11'b00110100000: data <= 32'h39fc3d74;
    11'b00110100001: data <= 32'ha8023d61;
    11'b00110100010: data <= 32'hb938ba31;
    11'b00110100011: data <= 32'hb4c6c196;
    11'b00110100100: data <= 32'h3432c103;
    11'b00110100101: data <= 32'h2a35b966;
    11'b00110100110: data <= 32'hb5d03522;
    11'b00110100111: data <= 32'h2cf0acb8;
    11'b00110101000: data <= 32'h39bbb4bb;
    11'b00110101001: data <= 32'hadbb37c3;
    11'b00110101010: data <= 32'hc0383c8e;
    11'b00110101011: data <= 32'hc1ed3954;
    11'b00110101100: data <= 32'hbd7eb0c0;
    11'b00110101101: data <= 32'h3ae1b150;
    11'b00110101110: data <= 32'h3d5e344c;
    11'b00110101111: data <= 32'h3591340d;
    11'b00110110000: data <= 32'h216831f6;
    11'b00110110001: data <= 32'h3b603c2f;
    11'b00110110010: data <= 32'h3dd74061;
    11'b00110110011: data <= 32'h38b73efa;
    11'b00110110100: data <= 32'hb82cb7d0;
    11'b00110110101: data <= 32'hb738c073;
    11'b00110110110: data <= 32'h362fbef0;
    11'b00110110111: data <= 32'h3a2fb428;
    11'b00110111000: data <= 32'h39b9aca1;
    11'b00110111001: data <= 32'h3b8bbc66;
    11'b00110111010: data <= 32'h3c32bd21;
    11'b00110111011: data <= 32'hacf72b29;
    11'b00110111100: data <= 32'hbfef3ca0;
    11'b00110111101: data <= 32'hc1423891;
    11'b00110111110: data <= 32'hbd03ba03;
    11'b00110111111: data <= 32'h348cbc6d;
    11'b00111000000: data <= 32'h2ffab754;
    11'b00111000001: data <= 32'hbafd2f7e;
    11'b00111000010: data <= 32'hb8b83801;
    11'b00111000011: data <= 32'h3ba73d74;
    11'b00111000100: data <= 32'h3e4c4093;
    11'b00111000101: data <= 32'h34733f90;
    11'b00111000110: data <= 32'hbcc3314d;
    11'b00111000111: data <= 32'hbb8ebc04;
    11'b00111001000: data <= 32'h3801b7b6;
    11'b00111001001: data <= 32'h3d9e35a6;
    11'b00111001010: data <= 32'h3d99b3ed;
    11'b00111001011: data <= 32'h3d70be35;
    11'b00111001100: data <= 32'h3d65bd91;
    11'b00111001101: data <= 32'h38273602;
    11'b00111001110: data <= 32'hbb903da9;
    11'b00111001111: data <= 32'hbe3b3438;
    11'b00111010000: data <= 32'hba54be6e;
    11'b00111010001: data <= 32'haf02c00e;
    11'b00111010010: data <= 32'hb993bc1e;
    11'b00111010011: data <= 32'hbdbdb142;
    11'b00111010100: data <= 32'hb90a2f4b;
    11'b00111010101: data <= 32'h3c2d393c;
    11'b00111010110: data <= 32'h3ce13e2e;
    11'b00111010111: data <= 32'hb9003ec7;
    11'b00111011000: data <= 32'hc05e3a6e;
    11'b00111011001: data <= 32'hbe0d2ff9;
    11'b00111011010: data <= 32'h3655370e;
    11'b00111011011: data <= 32'h3d753960;
    11'b00111011100: data <= 32'h3c71b454;
    11'b00111011101: data <= 32'h3bf9bd4a;
    11'b00111011110: data <= 32'h3db9b93f;
    11'b00111011111: data <= 32'h3d6e3d04;
    11'b00111100000: data <= 32'h35e63f71;
    11'b00111100001: data <= 32'hb71f2f32;
    11'b00111100010: data <= 32'hb5acbfea;
    11'b00111100011: data <= 32'hb262c05f;
    11'b00111100100: data <= 32'hb9e3bc07;
    11'b00111100101: data <= 32'hbc2ab6e4;
    11'b00111100110: data <= 32'ha5e7ba5e;
    11'b00111100111: data <= 32'h3d2fb97c;
    11'b00111101000: data <= 32'h3aa236ec;
    11'b00111101001: data <= 32'hbd6c3d4e;
    11'b00111101010: data <= 32'hc1763c66;
    11'b00111101011: data <= 32'hbef73830;
    11'b00111101100: data <= 32'h2e433789;
    11'b00111101101: data <= 32'h38983695;
    11'b00111101110: data <= 32'hac9db503;
    11'b00111101111: data <= 32'h2951ba40;
    11'b00111110000: data <= 32'h3d11347a;
    11'b00111110001: data <= 32'h3fd44016;
    11'b00111110010: data <= 32'h3ca6406c;
    11'b00111110011: data <= 32'ha0ef34b6;
    11'b00111110100: data <= 32'hb4fbbdf8;
    11'b00111110101: data <= 32'hae80bd59;
    11'b00111110110: data <= 32'hb18eb528;
    11'b00111110111: data <= 32'hae46b819;
    11'b00111111000: data <= 32'h3a6abeca;
    11'b00111111001: data <= 32'h3e79bf58;
    11'b00111111010: data <= 32'h3a52b51e;
    11'b00111111011: data <= 32'hbd213c71;
    11'b00111111100: data <= 32'hc0a93c08;
    11'b00111111101: data <= 32'hbd882e2a;
    11'b00111111110: data <= 32'hb204b4d0;
    11'b00111111111: data <= 32'hb825b432;
    11'b01000000000: data <= 32'hbdceb784;
    11'b01000000001: data <= 32'hbb28b773;
    11'b01000000010: data <= 32'h3c2338fe;
    11'b01000000011: data <= 32'h4019402e;
    11'b01000000100: data <= 32'h3c234053;
    11'b01000000101: data <= 32'hb7a13985;
    11'b01000000110: data <= 32'hb9d5b640;
    11'b01000000111: data <= 32'ha6892c46;
    11'b01000001000: data <= 32'h36a3390f;
    11'b01000001001: data <= 32'h38aeb653;
    11'b01000001010: data <= 32'h3cbec035;
    11'b01000001011: data <= 32'h3f14c045;
    11'b01000001100: data <= 32'h3cadb38c;
    11'b01000001101: data <= 32'hb5ac3d0d;
    11'b01000001110: data <= 32'hbc7a39f3;
    11'b01000001111: data <= 32'hb8a7b970;
    11'b01000010000: data <= 32'hb45ebcc3;
    11'b01000010001: data <= 32'hbd1aba81;
    11'b01000010010: data <= 32'hc06ab936;
    11'b01000010011: data <= 32'hbcd0b973;
    11'b01000010100: data <= 32'h3bda2284;
    11'b01000010101: data <= 32'h3eed3ce7;
    11'b01000010110: data <= 32'h33a83e92;
    11'b01000010111: data <= 32'hbda13c0e;
    11'b01000011000: data <= 32'hbd203949;
    11'b01000011001: data <= 32'hacc83cc2;
    11'b01000011010: data <= 32'h37f53d04;
    11'b01000011011: data <= 32'h360cb3a4;
    11'b01000011100: data <= 32'h39c3bf99;
    11'b01000011101: data <= 32'h3e3abe1e;
    11'b01000011110: data <= 32'h3ecd3864;
    11'b01000011111: data <= 32'h3afc3ec1;
    11'b01000100000: data <= 32'h32473892;
    11'b01000100001: data <= 32'h31f9bc82;
    11'b01000100010: data <= 32'hb0a7bda8;
    11'b01000100011: data <= 32'hbd4db9b6;
    11'b01000100100: data <= 32'hbfddb94c;
    11'b01000100101: data <= 32'hb9d0bd38;
    11'b01000100110: data <= 32'h3cccbcf2;
    11'b01000100111: data <= 32'h3d61ad94;
    11'b01000101000: data <= 32'hb8373b5f;
    11'b01000101001: data <= 32'hc0013c3b;
    11'b01000101010: data <= 32'hbdd33c38;
    11'b01000101011: data <= 32'hb1363d94;
    11'b01000101100: data <= 32'ha8da3ca8;
    11'b01000101101: data <= 32'hb9b6b33c;
    11'b01000101110: data <= 32'hb6cabd84;
    11'b01000101111: data <= 32'h3c20b8c1;
    11'b01000110000: data <= 32'h400b3d79;
    11'b01000110001: data <= 32'h3e974004;
    11'b01000110010: data <= 32'h3a9f38b9;
    11'b01000110011: data <= 32'h3727bae3;
    11'b01000110100: data <= 32'h2919b938;
    11'b01000110101: data <= 32'hba5430a2;
    11'b01000110110: data <= 32'hbc3bb63d;
    11'b01000110111: data <= 32'h2ed8bfa8;
    11'b01000111000: data <= 32'h3e08c0b6;
    11'b01000111001: data <= 32'h3cbfbc36;
    11'b01000111010: data <= 32'hb91a3714;
    11'b01000111011: data <= 32'hbebf3ab9;
    11'b01000111100: data <= 32'hbb933942;
    11'b01000111101: data <= 32'haf45398b;
    11'b01000111110: data <= 32'hbab13815;
    11'b01000111111: data <= 32'hc01bb60a;
    11'b01001000000: data <= 32'hbe59bbdf;
    11'b01001000001: data <= 32'h37f2ae71;
    11'b01001000010: data <= 32'h3fc93dfe;
    11'b01001000011: data <= 32'h3e2d3f58;
    11'b01001000100: data <= 32'h376e396f;
    11'b01001000101: data <= 32'h2d92a9aa;
    11'b01001000110: data <= 32'h2ff239a7;
    11'b01001000111: data <= 32'hb10d3d55;
    11'b01001001000: data <= 32'hb42b2bba;
    11'b01001001001: data <= 32'h3894c03d;
    11'b01001001010: data <= 32'h3e46c158;
    11'b01001001011: data <= 32'h3d2ebc6c;
    11'b01001001100: data <= 32'h24ed37de;
    11'b01001001101: data <= 32'hb8313868;
    11'b01001001110: data <= 32'h2d99b072;
    11'b01001001111: data <= 32'h30f4b467;
    11'b01001010000: data <= 32'hbd76af63;
    11'b01001010001: data <= 32'hc1a5b803;
    11'b01001010010: data <= 32'hc021bbc8;
    11'b01001010011: data <= 32'h34aab75d;
    11'b01001010100: data <= 32'h3e503987;
    11'b01001010101: data <= 32'h39f43c5e;
    11'b01001010110: data <= 32'hb80f3921;
    11'b01001010111: data <= 32'hb8343a13;
    11'b01001011000: data <= 32'h2ed03f5d;
    11'b01001011001: data <= 32'h2eeb404f;
    11'b01001011010: data <= 32'hb3a336b1;
    11'b01001011011: data <= 32'h31a1bf56;
    11'b01001011100: data <= 32'h3c9ec025;
    11'b01001011101: data <= 32'h3de1b50d;
    11'b01001011110: data <= 32'h3be63ba4;
    11'b01001011111: data <= 32'h3a6835cf;
    11'b01001100000: data <= 32'h3c58b9d6;
    11'b01001100001: data <= 32'h3841b99d;
    11'b01001100010: data <= 32'hbd35ae26;
    11'b01001100011: data <= 32'hc131b579;
    11'b01001100100: data <= 32'hbe7cbd07;
    11'b01001100101: data <= 32'h3821bdc7;
    11'b01001100110: data <= 32'h3cb9b903;
    11'b01001100111: data <= 32'hb03b2fad;
    11'b01001101000: data <= 32'hbd203648;
    11'b01001101001: data <= 32'hba513c0a;
    11'b01001101010: data <= 32'h30e94024;
    11'b01001101011: data <= 32'haf7b4048;
    11'b01001101100: data <= 32'hbc46376c;
    11'b01001101101: data <= 32'hbbb6bd30;
    11'b01001101110: data <= 32'h35e8bc37;
    11'b01001101111: data <= 32'h3ddc393d;
    11'b01001110000: data <= 32'h3e5b3d78;
    11'b01001110001: data <= 32'h3ddd347c;
    11'b01001110010: data <= 32'h3de0b9ec;
    11'b01001110011: data <= 32'h3a62b243;
    11'b01001110100: data <= 32'hb9eb39f6;
    11'b01001110101: data <= 32'hbe8431f1;
    11'b01001110110: data <= 32'hb952be16;
    11'b01001110111: data <= 32'h3b55c0bc;
    11'b01001111000: data <= 32'h3b9bbe88;
    11'b01001111001: data <= 32'hb7cbb839;
    11'b01001111010: data <= 32'hbcd72928;
    11'b01001111011: data <= 32'hb5013881;
    11'b01001111100: data <= 32'h37153d55;
    11'b01001111101: data <= 32'hb8873d9b;
    11'b01001111110: data <= 32'hc0643363;
    11'b01001111111: data <= 32'hc058bad4;
    11'b01010000000: data <= 32'hb5ffb58f;
    11'b01010000001: data <= 32'h3ccf3c17;
    11'b01010000010: data <= 32'h3da63cfc;
    11'b01010000011: data <= 32'h3c5b30e8;
    11'b01010000100: data <= 32'h3c44b448;
    11'b01010000101: data <= 32'h3a953b8a;
    11'b01010000110: data <= 32'hacb93feb;
    11'b01010000111: data <= 32'hb9333b02;
    11'b01010001000: data <= 32'h271cbdf7;
    11'b01010001001: data <= 32'h3c33c12b;
    11'b01010001010: data <= 32'h3afdbec6;
    11'b01010001011: data <= 32'hb12ab7c6;
    11'b01010001100: data <= 32'hb46cb332;
    11'b01010001101: data <= 32'h3a1cb428;
    11'b01010001110: data <= 32'h3bc532d1;
    11'b01010001111: data <= 32'hba943881;
    11'b01010010000: data <= 32'hc1b02412;
    11'b01010010001: data <= 32'hc15ab984;
    11'b01010010010: data <= 32'hb91db64a;
    11'b01010010011: data <= 32'h3a813734;
    11'b01010010100: data <= 32'h38a5378c;
    11'b01010010101: data <= 32'h9e50b0f0;
    11'b01010010110: data <= 32'h343b3390;
    11'b01010010111: data <= 32'h39a13fc2;
    11'b01010011000: data <= 32'h34fd41b3;
    11'b01010011001: data <= 32'hb55e3d62;
    11'b01010011010: data <= 32'hb003bc8c;
    11'b01010011011: data <= 32'h38fdbfc6;
    11'b01010011100: data <= 32'h3a40ba75;
    11'b01010011101: data <= 32'h37d03053;
    11'b01010011110: data <= 32'h3b2db501;
    11'b01010011111: data <= 32'h3f50bb8b;
    11'b01010100000: data <= 32'h3e0ab7b8;
    11'b01010100001: data <= 32'hb9203555;
    11'b01010100010: data <= 32'hc120311f;
    11'b01010100011: data <= 32'hc055b9ca;
    11'b01010100100: data <= 32'hb4bfbc33;
    11'b01010100101: data <= 32'h3803b99b;
    11'b01010100110: data <= 32'hb5e9b8a0;
    11'b01010100111: data <= 32'hbc19b8df;
    11'b01010101000: data <= 32'hb4003526;
    11'b01010101001: data <= 32'h39aa4035;
    11'b01010101010: data <= 32'h3500419a;
    11'b01010101011: data <= 32'hbab03d47;
    11'b01010101100: data <= 32'hbc55b94a;
    11'b01010101101: data <= 32'hb3b5bae4;
    11'b01010101110: data <= 32'h384a362b;
    11'b01010101111: data <= 32'h3b103a5c;
    11'b01010110000: data <= 32'h3df2b544;
    11'b01010110001: data <= 32'h406cbc9a;
    11'b01010110010: data <= 32'h3f0ab4cc;
    11'b01010110011: data <= 32'haed53bce;
    11'b01010110100: data <= 32'hbe273a10;
    11'b01010110101: data <= 32'hbc0cb9d3;
    11'b01010110110: data <= 32'h3574beec;
    11'b01010110111: data <= 32'h35adbe7b;
    11'b01010111000: data <= 32'hbb2abd0b;
    11'b01010111001: data <= 32'hbd14bc04;
    11'b01010111010: data <= 32'h219bb057;
    11'b01010111011: data <= 32'h3c323d3e;
    11'b01010111100: data <= 32'h30223f91;
    11'b01010111101: data <= 32'hbec93af4;
    11'b01010111110: data <= 32'hc062b4f9;
    11'b01010111111: data <= 32'hbc329ef2;
    11'b01011000000: data <= 32'h31863c3e;
    11'b01011000001: data <= 32'h39353b40;
    11'b01011000010: data <= 32'h3c3ab7bf;
    11'b01011000011: data <= 32'h3eb5bb83;
    11'b01011000100: data <= 32'h3e64386d;
    11'b01011000101: data <= 32'h37784032;
    11'b01011000110: data <= 32'hb6e23e21;
    11'b01011000111: data <= 32'ha548b85d;
    11'b01011001000: data <= 32'h39c9bf65;
    11'b01011001001: data <= 32'h346cbe83;
    11'b01011001010: data <= 32'hba8ebc84;
    11'b01011001011: data <= 32'hb910bc82;
    11'b01011001100: data <= 32'h3bb0bb08;
    11'b01011001101: data <= 32'h3eb12d0d;
    11'b01011001110: data <= 32'h2c2c3a25;
    11'b01011001111: data <= 32'hc0693647;
    11'b01011010000: data <= 32'hc149b18c;
    11'b01011010001: data <= 32'hbd1131d6;
    11'b01011010010: data <= 32'hb01e3a60;
    11'b01011010011: data <= 32'haff13470;
    11'b01011010100: data <= 32'hb065bb1c;
    11'b01011010101: data <= 32'h38e3b941;
    11'b01011010110: data <= 32'h3cdb3d84;
    11'b01011010111: data <= 32'h3a6741d4;
    11'b01011011000: data <= 32'h2e813ffe;
    11'b01011011001: data <= 32'h30a3b312;
    11'b01011011010: data <= 32'h377ebced;
    11'b01011011011: data <= 32'h2e32b93a;
    11'b01011011100: data <= 32'hb694b45b;
    11'b01011011101: data <= 32'h3579bbb0;
    11'b01011011110: data <= 32'h3fe2bdf8;
    11'b01011011111: data <= 32'h407eba86;
    11'b01011100000: data <= 32'h345e32ca;
    11'b01011100001: data <= 32'hbfab3561;
    11'b01011100010: data <= 32'hc01bb077;
    11'b01011100011: data <= 32'hb9cab31a;
    11'b01011100100: data <= 32'hb2b3b028;
    11'b01011100101: data <= 32'hbbffb9b4;
    11'b01011100110: data <= 32'hbd5abda7;
    11'b01011100111: data <= 32'hb373b934;
    11'b01011101000: data <= 32'h3beb3e04;
    11'b01011101001: data <= 32'h3abd4199;
    11'b01011101010: data <= 32'hb0a23f41;
    11'b01011101011: data <= 32'hb8822b71;
    11'b01011101100: data <= 32'hb52eb308;
    11'b01011101101: data <= 32'hb3c039a9;
    11'b01011101110: data <= 32'hb09639b6;
    11'b01011101111: data <= 32'h3ae4b9d1;
    11'b01011110000: data <= 32'h409bbedc;
    11'b01011110001: data <= 32'h40c5bb10;
    11'b01011110010: data <= 32'h393b38a7;
    11'b01011110011: data <= 32'hbb983ab7;
    11'b01011110100: data <= 32'hb9f4a90d;
    11'b01011110101: data <= 32'h3362b9e5;
    11'b01011110110: data <= 32'hadffbb9a;
    11'b01011110111: data <= 32'hbe10bd70;
    11'b01011111000: data <= 32'hbf4fbefe;
    11'b01011111001: data <= 32'hb442bc05;
    11'b01011111010: data <= 32'h3cd53a06;
    11'b01011111011: data <= 32'h3a173f00;
    11'b01011111100: data <= 32'hba793c41;
    11'b01011111101: data <= 32'hbe2c3098;
    11'b01011111110: data <= 32'hbc6a38df;
    11'b01011111111: data <= 32'hb8c53e7c;
    11'b01100000000: data <= 32'hb53a3c8f;
    11'b01100000001: data <= 32'h3747b9d3;
    11'b01100000010: data <= 32'h3e99be5f;
    11'b01100000011: data <= 32'h3fd2b3d4;
    11'b01100000100: data <= 32'h3bc53e30;
    11'b01100000101: data <= 32'h2fcf3e5a;
    11'b01100000110: data <= 32'h37b031a2;
    11'b01100000111: data <= 32'h3b92bacd;
    11'b01100001000: data <= 32'h233dbbad;
    11'b01100001001: data <= 32'hbe0ebc87;
    11'b01100001010: data <= 32'hbdadbe94;
    11'b01100001011: data <= 32'h37febe0e;
    11'b01100001100: data <= 32'h3f32b6ff;
    11'b01100001101: data <= 32'h3a17366b;
    11'b01100001110: data <= 32'hbd1133aa;
    11'b01100001111: data <= 32'hbfe62c23;
    11'b01100010000: data <= 32'hbd023ad3;
    11'b01100010001: data <= 32'hb9c43e64;
    11'b01100010010: data <= 32'hbb3739cd;
    11'b01100010011: data <= 32'hb995bc56;
    11'b01100010100: data <= 32'h35ecbd94;
    11'b01100010101: data <= 32'h3ce037d4;
    11'b01100010110: data <= 32'h3c4140a5;
    11'b01100010111: data <= 32'h39864003;
    11'b01100011000: data <= 32'h3b303606;
    11'b01100011001: data <= 32'h3b85b63e;
    11'b01100011010: data <= 32'hae06a543;
    11'b01100011011: data <= 32'hbccdad30;
    11'b01100011100: data <= 32'hb88fbc8b;
    11'b01100011101: data <= 32'h3dcabf7e;
    11'b01100011110: data <= 32'h40b1bd68;
    11'b01100011111: data <= 32'h3b2bb6a9;
    11'b01100100000: data <= 32'hbc5cae71;
    11'b01100100001: data <= 32'hbda69c90;
    11'b01100100010: data <= 32'hb84d385e;
    11'b01100100011: data <= 32'hb7b63a9f;
    11'b01100100100: data <= 32'hbe17b1cc;
    11'b01100100101: data <= 32'hbfa0be62;
    11'b01100100110: data <= 32'hb9ebbd72;
    11'b01100100111: data <= 32'h396d3975;
    11'b01100101000: data <= 32'h3bbc4074;
    11'b01100101001: data <= 32'h38483eb7;
    11'b01100101010: data <= 32'h35ff35ed;
    11'b01100101011: data <= 32'h342e3613;
    11'b01100101100: data <= 32'hb6cf3d5d;
    11'b01100101101: data <= 32'hbb923caf;
    11'b01100101110: data <= 32'ha5cdb87a;
    11'b01100101111: data <= 32'h3f2cbfaf;
    11'b01100110000: data <= 32'h40bfbdff;
    11'b01100110001: data <= 32'h3c22b41f;
    11'b01100110010: data <= 32'hb57c340b;
    11'b01100110011: data <= 32'haec12d2a;
    11'b01100110100: data <= 32'h396e2ce4;
    11'b01100110101: data <= 32'ha0f124e6;
    11'b01100110110: data <= 32'hbf5abaaa;
    11'b01100110111: data <= 32'hc0edbf6b;
    11'b01100111000: data <= 32'hbc07be16;
    11'b01100111001: data <= 32'h39a43002;
    11'b01100111010: data <= 32'h3acf3cbb;
    11'b01100111011: data <= 32'hac07396c;
    11'b01100111100: data <= 32'hb8712e1e;
    11'b01100111101: data <= 32'hb81a3be9;
    11'b01100111110: data <= 32'hb9e240a1;
    11'b01100111111: data <= 32'hbbe43f6a;
    11'b01101000000: data <= 32'hb442b53e;
    11'b01101000001: data <= 32'h3c99bef3;
    11'b01101000010: data <= 32'h3edabb82;
    11'b01101000011: data <= 32'h3bff38fa;
    11'b01101000100: data <= 32'h38003bcf;
    11'b01101000101: data <= 32'h3cb43469;
    11'b01101000110: data <= 32'h3eafb029;
    11'b01101000111: data <= 32'h35f2afa8;
    11'b01101001000: data <= 32'hbef8b8fd;
    11'b01101001001: data <= 32'hc047be36;
    11'b01101001010: data <= 32'hb5c7becd;
    11'b01101001011: data <= 32'h3cfbbab0;
    11'b01101001100: data <= 32'h3abfb2f8;
    11'b01101001101: data <= 32'hb88fb704;
    11'b01101001110: data <= 32'hbc54b4b2;
    11'b01101001111: data <= 32'hb97a3c71;
    11'b01101010000: data <= 32'hb99940c2;
    11'b01101010001: data <= 32'hbd103e5f;
    11'b01101010010: data <= 32'hbccab8cd;
    11'b01101010011: data <= 32'hb18ebe21;
    11'b01101010100: data <= 32'h396bb20c;
    11'b01101010101: data <= 32'h3a053dd6;
    11'b01101010110: data <= 32'h3b593daf;
    11'b01101010111: data <= 32'h3ebc35b1;
    11'b01101011000: data <= 32'h3f6c2ceb;
    11'b01101011001: data <= 32'h363138e5;
    11'b01101011010: data <= 32'hbda83763;
    11'b01101011011: data <= 32'hbd34b9ff;
    11'b01101011100: data <= 32'h38f0bed0;
    11'b01101011101: data <= 32'h3f45be4f;
    11'b01101011110: data <= 32'h3b25bc84;
    11'b01101011111: data <= 32'hb8cfbc09;
    11'b01101100000: data <= 32'hb9a8b841;
    11'b01101100001: data <= 32'h2aa53a2d;
    11'b01101100010: data <= 32'hb1e93e92;
    11'b01101100011: data <= 32'hbe1c3985;
    11'b01101100100: data <= 32'hc06fbc85;
    11'b01101100101: data <= 32'hbd84bdc7;
    11'b01101100110: data <= 32'hb0203168;
    11'b01101100111: data <= 32'h36fe3e1f;
    11'b01101101000: data <= 32'h39ae3c56;
    11'b01101101001: data <= 32'h3cdc2e72;
    11'b01101101010: data <= 32'h3cdf37ff;
    11'b01101101011: data <= 32'h2ad13f1c;
    11'b01101101100: data <= 32'hbc833f3c;
    11'b01101101101: data <= 32'hb9052f9d;
    11'b01101101110: data <= 32'h3c71bdf3;
    11'b01101101111: data <= 32'h3f68be95;
    11'b01101110000: data <= 32'h3a86bc2c;
    11'b01101110001: data <= 32'hb1bbb9ee;
    11'b01101110010: data <= 32'h3676b78d;
    11'b01101110011: data <= 32'h3d6f348e;
    11'b01101110100: data <= 32'h38c739f5;
    11'b01101110101: data <= 32'hbe2cadc1;
    11'b01101110110: data <= 32'hc157bda7;
    11'b01101110111: data <= 32'hbef0bdb5;
    11'b01101111000: data <= 32'hb386add0;
    11'b01101111001: data <= 32'h341f3971;
    11'b01101111010: data <= 32'h2e2a1436;
    11'b01101111011: data <= 32'h3358b7d8;
    11'b01101111100: data <= 32'h35743a48;
    11'b01101111101: data <= 32'hb4b64142;
    11'b01101111110: data <= 32'hbc1f412f;
    11'b01101111111: data <= 32'hb8d93841;
    11'b01110000000: data <= 32'h3941bcc6;
    11'b01110000001: data <= 32'h3c7dbc3f;
    11'b01110000010: data <= 32'h3787b06b;
    11'b01110000011: data <= 32'h353a2ae2;
    11'b01110000100: data <= 32'h3e32b388;
    11'b01110000101: data <= 32'h40efa59e;
    11'b01110000110: data <= 32'h3cd13601;
    11'b01110000111: data <= 32'hbd2aac47;
    11'b01110001000: data <= 32'hc09ebc41;
    11'b01110001001: data <= 32'hbc5dbd40;
    11'b01110001010: data <= 32'h3569b9b1;
    11'b01110001011: data <= 32'h3486b89b;
    11'b01110001100: data <= 32'hb7b7bcf9;
    11'b01110001101: data <= 32'hb7e2bc94;
    11'b01110001110: data <= 32'ha1da39a6;
    11'b01110001111: data <= 32'hb39d4149;
    11'b01110010000: data <= 32'hbc2f40b9;
    11'b01110010001: data <= 32'hbccf344e;
    11'b01110010010: data <= 32'hb81abc01;
    11'b01110010011: data <= 32'ha9d9b425;
    11'b01110010100: data <= 32'hacc43ae2;
    11'b01110010101: data <= 32'h3809395b;
    11'b01110010110: data <= 32'h3ffbb0d1;
    11'b01110010111: data <= 32'h416ca986;
    11'b01110011000: data <= 32'h3d1d3a4d;
    11'b01110011001: data <= 32'hbb923ad8;
    11'b01110011010: data <= 32'hbdb5b043;
    11'b01110011011: data <= 32'h24c5bbfa;
    11'b01110011100: data <= 32'h3c43bcb7;
    11'b01110011101: data <= 32'h35b7bda7;
    11'b01110011110: data <= 32'hb9a2bf9f;
    11'b01110011111: data <= 32'hb6a9bdfc;
    11'b01110100000: data <= 32'h386f3507;
    11'b01110100001: data <= 32'h363a3f78;
    11'b01110100010: data <= 32'hbbe13d70;
    11'b01110100011: data <= 32'hbfb2b655;
    11'b01110100100: data <= 32'hbe89bb9b;
    11'b01110100101: data <= 32'hbbc6341b;
    11'b01110100110: data <= 32'hb8783cd5;
    11'b01110100111: data <= 32'h326e3816;
    11'b01110101000: data <= 32'h3df4b7ed;
    11'b01110101001: data <= 32'h40042c35;
    11'b01110101010: data <= 32'h3ab53e92;
    11'b01110101011: data <= 32'hb99a4037;
    11'b01110101100: data <= 32'hb8fe3b04;
    11'b01110101101: data <= 32'h3a22b87d;
    11'b01110101110: data <= 32'h3d24bc6f;
    11'b01110101111: data <= 32'h32edbd28;
    11'b01110110000: data <= 32'hb89fbe71;
    11'b01110110001: data <= 32'h3617bd7b;
    11'b01110110010: data <= 32'h3f06b07b;
    11'b01110110011: data <= 32'h3d4d3ae7;
    11'b01110110100: data <= 32'hb9e8358a;
    11'b01110110101: data <= 32'hc065baf5;
    11'b01110110110: data <= 32'hbfccbb30;
    11'b01110110111: data <= 32'hbc5f344a;
    11'b01110111000: data <= 32'hb9c9395d;
    11'b01110111001: data <= 32'hb661b74f;
    11'b01110111010: data <= 32'h36a8bcf9;
    11'b01110111011: data <= 32'h3b652bca;
    11'b01110111100: data <= 32'h34cb4090;
    11'b01110111101: data <= 32'hb8c441b3;
    11'b01110111110: data <= 32'hb5bc3d62;
    11'b01110111111: data <= 32'h38fbb339;
    11'b01111000000: data <= 32'h397eb813;
    11'b01111000001: data <= 32'hb476b4fd;
    11'b01111000010: data <= 32'hb60eb91e;
    11'b01111000011: data <= 32'h3d27bb9e;
    11'b01111000100: data <= 32'h41a4b6e8;
    11'b01111000101: data <= 32'h400d3470;
    11'b01111000110: data <= 32'hb6322c21;
    11'b01111000111: data <= 32'hbf25b95b;
    11'b01111001000: data <= 32'hbcf9b934;
    11'b01111001001: data <= 32'hb618a918;
    11'b01111001010: data <= 32'hb84fb53f;
    11'b01111001011: data <= 32'hbb99be9f;
    11'b01111001100: data <= 32'hb7ebc00d;
    11'b01111001101: data <= 32'h3465b17e;
    11'b01111001110: data <= 32'h31f2406b;
    11'b01111001111: data <= 32'hb8074122;
    11'b01111010000: data <= 32'hb92a3be3;
    11'b01111010001: data <= 32'hb462b10d;
    11'b01111010010: data <= 32'hb6e13440;
    11'b01111010011: data <= 32'hbbd53ad1;
    11'b01111010100: data <= 32'hb66e342a;
    11'b01111010101: data <= 32'h3e78b96e;
    11'b01111010110: data <= 32'h420cb83d;
    11'b01111010111: data <= 32'h40193649;
    11'b01111011000: data <= 32'hafdf399a;
    11'b01111011001: data <= 32'hbb603249;
    11'b01111011010: data <= 32'h2229b13d;
    11'b01111011011: data <= 32'h38eab441;
    11'b01111011100: data <= 32'hb440bc15;
    11'b01111011101: data <= 32'hbce0c094;
    11'b01111011110: data <= 32'hb995c0c0;
    11'b01111011111: data <= 32'h3859b842;
    11'b01111100000: data <= 32'h39d23dbc;
    11'b01111100001: data <= 32'hb4503dbd;
    11'b01111100010: data <= 32'hbc632ce8;
    11'b01111100011: data <= 32'hbce4b4e6;
    11'b01111100100: data <= 32'hbd5c3a72;
    11'b01111100101: data <= 32'hbe0d3dd8;
    11'b01111100110: data <= 32'hb9d63682;
    11'b01111100111: data <= 32'h3c5cbb4f;
    11'b01111101000: data <= 32'h406cb8a7;
    11'b01111101001: data <= 32'h3d953bae;
    11'b01111101010: data <= 32'hac453f06;
    11'b01111101011: data <= 32'haf0c3cc8;
    11'b01111101100: data <= 32'h3c0435e5;
    11'b01111101101: data <= 32'h3c93af67;
    11'b01111101110: data <= 32'hb453bad4;
    11'b01111101111: data <= 32'hbcefbfa2;
    11'b01111110000: data <= 32'hb240c027;
    11'b01111110001: data <= 32'h3e1cba8c;
    11'b01111110010: data <= 32'h3e9b36dd;
    11'b01111110011: data <= 32'h2eff322e;
    11'b01111110100: data <= 32'hbcf4b9b1;
    11'b01111110101: data <= 32'hbde2b6a3;
    11'b01111110110: data <= 32'hbd9a3b7c;
    11'b01111110111: data <= 32'hbe383cdf;
    11'b01111111000: data <= 32'hbcc7b52c;
    11'b01111111001: data <= 32'h24c7be8f;
    11'b01111111010: data <= 32'h3b54b9f2;
    11'b01111111011: data <= 32'h385a3db1;
    11'b01111111100: data <= 32'hb0a040d0;
    11'b01111111101: data <= 32'h34023e83;
    11'b01111111110: data <= 32'h3c9e3918;
    11'b01111111111: data <= 32'h3a6d364a;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    