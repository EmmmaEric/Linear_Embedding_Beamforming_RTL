
module memory_rom_29(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h26e5be56;
    11'b00000000001: data <= 32'ha862bb05;
    11'b00000000010: data <= 32'habc33b9a;
    11'b00000000011: data <= 32'hbb2d3e95;
    11'b00000000100: data <= 32'hbee82dba;
    11'b00000000101: data <= 32'hbe0abf3f;
    11'b00000000110: data <= 32'hba15bea7;
    11'b00000000111: data <= 32'hb84c306a;
    11'b00000001000: data <= 32'hb81d3d03;
    11'b00000001001: data <= 32'h35383b09;
    11'b00000001010: data <= 32'h3ddd3807;
    11'b00000001011: data <= 32'h3caf3ca3;
    11'b00000001100: data <= 32'hb9533f39;
    11'b00000001101: data <= 32'hbf213cd8;
    11'b00000001110: data <= 32'hb89da8d2;
    11'b00000001111: data <= 32'h3e08b92e;
    11'b00000010000: data <= 32'h4003b94f;
    11'b00000010001: data <= 32'h3b1abb81;
    11'b00000010010: data <= 32'h33c5bccc;
    11'b00000010011: data <= 32'h3b3ab6a7;
    11'b00000010100: data <= 32'h3d4a3be6;
    11'b00000010101: data <= 32'h335a3c65;
    11'b00000010110: data <= 32'hbd67b93a;
    11'b00000010111: data <= 32'hbf0bc07d;
    11'b00000011000: data <= 32'hbc62befd;
    11'b00000011001: data <= 32'hb894ad2d;
    11'b00000011010: data <= 32'hb62b373d;
    11'b00000011011: data <= 32'h312db59f;
    11'b00000011100: data <= 32'h3a2fb7a5;
    11'b00000011101: data <= 32'h339e3bf6;
    11'b00000011110: data <= 32'hbd4340c8;
    11'b00000011111: data <= 32'hbfda3fe0;
    11'b00000100000: data <= 32'hb945365b;
    11'b00000100001: data <= 32'h3c17b804;
    11'b00000100010: data <= 32'h3c6eb620;
    11'b00000100011: data <= 32'h3139b370;
    11'b00000100100: data <= 32'h3514b445;
    11'b00000100101: data <= 32'h3f3733e4;
    11'b00000100110: data <= 32'h40ea3c70;
    11'b00000100111: data <= 32'h3bd83b8b;
    11'b00000101000: data <= 32'hbc42b8a4;
    11'b00000101001: data <= 32'hbe1abf20;
    11'b00000101010: data <= 32'hb85bbd56;
    11'b00000101011: data <= 32'h3201b593;
    11'b00000101100: data <= 32'h2f89b919;
    11'b00000101101: data <= 32'h2e0fbee2;
    11'b00000101110: data <= 32'h3529bda6;
    11'b00000101111: data <= 32'hae4b39bc;
    11'b00000110000: data <= 32'hbd1640c2;
    11'b00000110001: data <= 32'hbf563efa;
    11'b00000110010: data <= 32'hbc18ab6f;
    11'b00000110011: data <= 32'hacbbba13;
    11'b00000110100: data <= 32'hb494ad18;
    11'b00000110101: data <= 32'hba463806;
    11'b00000110110: data <= 32'h31743671;
    11'b00000110111: data <= 32'h4045380d;
    11'b00000111000: data <= 32'h415e3c91;
    11'b00000111001: data <= 32'h3b4a3d17;
    11'b00000111010: data <= 32'hbc4c3587;
    11'b00000111011: data <= 32'hbc34b899;
    11'b00000111100: data <= 32'h3606b85f;
    11'b00000111101: data <= 32'h3c3eb6af;
    11'b00000111110: data <= 32'h3825bd56;
    11'b00000111111: data <= 32'h2f55c0d4;
    11'b00001000000: data <= 32'h3762bef0;
    11'b00001000001: data <= 32'h38223851;
    11'b00001000010: data <= 32'hb6433f83;
    11'b00001000011: data <= 32'hbd473a93;
    11'b00001000100: data <= 32'hbd60bbb7;
    11'b00001000101: data <= 32'hbc4fbc97;
    11'b00001000110: data <= 32'hbd622c0f;
    11'b00001000111: data <= 32'hbd9f3987;
    11'b00001001000: data <= 32'hadb8321c;
    11'b00001001001: data <= 32'h3f159c7e;
    11'b00001001010: data <= 32'h3fe43b42;
    11'b00001001011: data <= 32'h31393f33;
    11'b00001001100: data <= 32'hbd513e28;
    11'b00001001101: data <= 32'hb966396d;
    11'b00001001110: data <= 32'h3b8e3262;
    11'b00001001111: data <= 32'h3d1eb2e1;
    11'b00001010000: data <= 32'h3582bcfa;
    11'b00001010001: data <= 32'h2c1fc029;
    11'b00001010010: data <= 32'h3c40bd36;
    11'b00001010011: data <= 32'h3ef738a6;
    11'b00001010100: data <= 32'h3af43d26;
    11'b00001010101: data <= 32'hb916abe9;
    11'b00001010110: data <= 32'hbd61be2f;
    11'b00001010111: data <= 32'hbd6abce4;
    11'b00001011000: data <= 32'hbdd62cc4;
    11'b00001011001: data <= 32'hbd6a3298;
    11'b00001011010: data <= 32'hb468bb06;
    11'b00001011011: data <= 32'h3c30bc75;
    11'b00001011100: data <= 32'h3b7236ae;
    11'b00001011101: data <= 32'hb8f54034;
    11'b00001011110: data <= 32'hbe164071;
    11'b00001011111: data <= 32'hb8853cdd;
    11'b00001100000: data <= 32'h3a02379b;
    11'b00001100001: data <= 32'h385a2ff2;
    11'b00001100010: data <= 32'hb7f6b81c;
    11'b00001100011: data <= 32'hb218bc4b;
    11'b00001100100: data <= 32'h3ea0b838;
    11'b00001100101: data <= 32'h419339d9;
    11'b00001100110: data <= 32'h3efc3bcf;
    11'b00001100111: data <= 32'hb156b413;
    11'b00001101000: data <= 32'hbc07bcfe;
    11'b00001101001: data <= 32'hba36b9af;
    11'b00001101010: data <= 32'hb9453020;
    11'b00001101011: data <= 32'hba23b887;
    11'b00001101100: data <= 32'hb4f0c04c;
    11'b00001101101: data <= 32'h379ec063;
    11'b00001101110: data <= 32'h35adade1;
    11'b00001101111: data <= 32'hb9fb3fc4;
    11'b00001110000: data <= 32'hbd453fdb;
    11'b00001110001: data <= 32'hb9023a0d;
    11'b00001110010: data <= 32'ha6623199;
    11'b00001110011: data <= 32'hb9f23667;
    11'b00001110100: data <= 32'hbe6b3506;
    11'b00001110101: data <= 32'hb8dfb226;
    11'b00001110110: data <= 32'h3f32adff;
    11'b00001110111: data <= 32'h41f339c0;
    11'b00001111000: data <= 32'h3ed43c1d;
    11'b00001111001: data <= 32'hb18135a8;
    11'b00001111010: data <= 32'hb853b106;
    11'b00001111011: data <= 32'h32f233c4;
    11'b00001111100: data <= 32'h365735cc;
    11'b00001111101: data <= 32'hb243bc29;
    11'b00001111110: data <= 32'hb4dcc19a;
    11'b00001111111: data <= 32'h35edc12a;
    11'b00010000000: data <= 32'h3948b538;
    11'b00010000001: data <= 32'h1d533dae;
    11'b00010000010: data <= 32'hb9253bda;
    11'b00010000011: data <= 32'hb8fcb4ce;
    11'b00010000100: data <= 32'hba3ab5f4;
    11'b00010000101: data <= 32'hbf093848;
    11'b00010000110: data <= 32'hc0a939b2;
    11'b00010000111: data <= 32'hbbdaaedc;
    11'b00010001000: data <= 32'h3d86b760;
    11'b00010001001: data <= 32'h406c3578;
    11'b00010001010: data <= 32'h3abe3ce8;
    11'b00010001011: data <= 32'hb8833d1a;
    11'b00010001100: data <= 32'hb1e83c30;
    11'b00010001101: data <= 32'h3bb73c83;
    11'b00010001110: data <= 32'h3b2a39dd;
    11'b00010001111: data <= 32'hb2c1bae2;
    11'b00010010000: data <= 32'hb785c0d8;
    11'b00010010001: data <= 32'h3935c025;
    11'b00010010010: data <= 32'h3e66b1ab;
    11'b00010010011: data <= 32'h3cd73acf;
    11'b00010010100: data <= 32'h3299ab3c;
    11'b00010010101: data <= 32'hb67dbc96;
    11'b00010010110: data <= 32'hbb6eb8f2;
    11'b00010010111: data <= 32'hbf5a3910;
    11'b00010011000: data <= 32'hc07d383e;
    11'b00010011001: data <= 32'hbc67bb10;
    11'b00010011010: data <= 32'h3962be04;
    11'b00010011011: data <= 32'h3c26b540;
    11'b00010011100: data <= 32'hb2013d13;
    11'b00010011101: data <= 32'hbb7f3f30;
    11'b00010011110: data <= 32'ha4623e3e;
    11'b00010011111: data <= 32'h3c363dad;
    11'b00010100000: data <= 32'h374f3c39;
    11'b00010100001: data <= 32'hbbc3b02f;
    11'b00010100010: data <= 32'hbb41bd35;
    11'b00010100011: data <= 32'h3ba8bc4b;
    11'b00010100100: data <= 32'h40e930fd;
    11'b00010100101: data <= 32'h40223810;
    11'b00010100110: data <= 32'h39ebb814;
    11'b00010100111: data <= 32'ha6f4bc98;
    11'b00010101000: data <= 32'hb544b2a8;
    11'b00010101001: data <= 32'hbb8d3ae2;
    11'b00010101010: data <= 32'hbddc2bf1;
    11'b00010101011: data <= 32'hbbaabfc5;
    11'b00010101100: data <= 32'h2dc5c123;
    11'b00010101101: data <= 32'h3318bb90;
    11'b00010101110: data <= 32'hb8f03c0a;
    11'b00010101111: data <= 32'hbadc3df6;
    11'b00010110000: data <= 32'h2cf93c1b;
    11'b00010110001: data <= 32'h38b13bbc;
    11'b00010110010: data <= 32'hb8cf3cb5;
    11'b00010110011: data <= 32'hc0203992;
    11'b00010110100: data <= 32'hbde0b283;
    11'b00010110101: data <= 32'h3b96b566;
    11'b00010110110: data <= 32'h412134b0;
    11'b00010110111: data <= 32'h3fe636dc;
    11'b00010111000: data <= 32'h390bb2be;
    11'b00010111001: data <= 32'h351eb4d8;
    11'b00010111010: data <= 32'h394a39cf;
    11'b00010111011: data <= 32'h34e73d0e;
    11'b00010111100: data <= 32'hb8c7b2f9;
    11'b00010111101: data <= 32'hba40c0fb;
    11'b00010111110: data <= 32'haf9bc1d8;
    11'b00010111111: data <= 32'h3328bc82;
    11'b00011000000: data <= 32'hb01c3883;
    11'b00011000001: data <= 32'hb2e33807;
    11'b00011000010: data <= 32'h3442b288;
    11'b00011000011: data <= 32'h2c0f3075;
    11'b00011000100: data <= 32'hbdf83c82;
    11'b00011000101: data <= 32'hc18c3cae;
    11'b00011000110: data <= 32'hbf5e319b;
    11'b00011000111: data <= 32'h3874b6c2;
    11'b00011001000: data <= 32'h3f24a769;
    11'b00011001001: data <= 32'h3ba93706;
    11'b00011001010: data <= 32'ha4973740;
    11'b00011001011: data <= 32'h37d83a0e;
    11'b00011001100: data <= 32'h3dda3e76;
    11'b00011001101: data <= 32'h3c593ec1;
    11'b00011001110: data <= 32'hb508a30c;
    11'b00011001111: data <= 32'hbae9c02a;
    11'b00011010000: data <= 32'ha468c091;
    11'b00011010001: data <= 32'h3b14ba0c;
    11'b00011010010: data <= 32'h3b47316e;
    11'b00011010011: data <= 32'h3930b89a;
    11'b00011010100: data <= 32'h38afbd47;
    11'b00011010101: data <= 32'ha2a8b6ad;
    11'b00011010110: data <= 32'hbe1c3c72;
    11'b00011010111: data <= 32'hc12e3c99;
    11'b00011011000: data <= 32'hbf20b4f8;
    11'b00011011001: data <= 32'h175bbd19;
    11'b00011011010: data <= 32'h389cb9b6;
    11'b00011011011: data <= 32'hb5463572;
    11'b00011011100: data <= 32'hb9a93ad3;
    11'b00011011101: data <= 32'h38243cda;
    11'b00011011110: data <= 32'h3ec53f5f;
    11'b00011011111: data <= 32'h3b8e3f89;
    11'b00011100000: data <= 32'hbadf38c0;
    11'b00011100001: data <= 32'hbd38bb71;
    11'b00011100010: data <= 32'h2ff9bc2d;
    11'b00011100011: data <= 32'h3e51aec7;
    11'b00011100100: data <= 32'h3ec8a2f8;
    11'b00011100101: data <= 32'h3c9bbc9a;
    11'b00011100110: data <= 32'h3b29be7d;
    11'b00011100111: data <= 32'h3809b3ea;
    11'b00011101000: data <= 32'hb8d43d4d;
    11'b00011101001: data <= 32'hbe5f3adb;
    11'b00011101010: data <= 32'hbd55bcb4;
    11'b00011101011: data <= 32'hb68bc080;
    11'b00011101100: data <= 32'hb584bd50;
    11'b00011101101: data <= 32'hbc432dfb;
    11'b00011101110: data <= 32'hbb2b38ad;
    11'b00011101111: data <= 32'h3898392f;
    11'b00011110000: data <= 32'h3d9e3cd0;
    11'b00011110001: data <= 32'h2ed13ee6;
    11'b00011110010: data <= 32'hbf623cfd;
    11'b00011110011: data <= 32'hbf8a3428;
    11'b00011110100: data <= 32'h2cd614a7;
    11'b00011110101: data <= 32'h3eba3538;
    11'b00011110110: data <= 32'h3e46a6a1;
    11'b00011110111: data <= 32'h3b22bc1b;
    11'b00011111000: data <= 32'h3c00bc14;
    11'b00011111001: data <= 32'h3d53387d;
    11'b00011111010: data <= 32'h39cf3f07;
    11'b00011111011: data <= 32'hb6b63948;
    11'b00011111100: data <= 32'hbab7beb5;
    11'b00011111101: data <= 32'hb82ac123;
    11'b00011111110: data <= 32'hb816bd99;
    11'b00011111111: data <= 32'hbabdb11c;
    11'b00100000000: data <= 32'hb680b42b;
    11'b00100000001: data <= 32'h3a57b93a;
    11'b00100000010: data <= 32'h3bfb2d27;
    11'b00100000011: data <= 32'hb99d3d61;
    11'b00100000100: data <= 32'hc1093e63;
    11'b00100000101: data <= 32'hc05f3a5f;
    11'b00100000110: data <= 32'hb19f328a;
    11'b00100000111: data <= 32'h3c0f321a;
    11'b00100001000: data <= 32'h37cea886;
    11'b00100001001: data <= 32'ha82db809;
    11'b00100001010: data <= 32'h3abdace5;
    11'b00100001011: data <= 32'h3ff63da2;
    11'b00100001100: data <= 32'h3e9e404b;
    11'b00100001101: data <= 32'h31783a38;
    11'b00100001110: data <= 32'hb994bd67;
    11'b00100001111: data <= 32'hb6b1bf80;
    11'b00100010000: data <= 32'ha01bba39;
    11'b00100010001: data <= 32'h29e7b3b5;
    11'b00100010010: data <= 32'h3684bcc3;
    11'b00100010011: data <= 32'h3c72bfa1;
    11'b00100010100: data <= 32'h3b17ba63;
    11'b00100010101: data <= 32'hba4e3c46;
    11'b00100010110: data <= 32'hc0943e31;
    11'b00100010111: data <= 32'hbfa437a3;
    11'b00100011000: data <= 32'hb71ab772;
    11'b00100011001: data <= 32'haa0eb6d0;
    11'b00100011010: data <= 32'hbb73b0ff;
    11'b00100011011: data <= 32'hbc37af8f;
    11'b00100011100: data <= 32'h38a23668;
    11'b00100011101: data <= 32'h40543e69;
    11'b00100011110: data <= 32'h3eba4057;
    11'b00100011111: data <= 32'hb1103c89;
    11'b00100100000: data <= 32'hbc2bb562;
    11'b00100100001: data <= 32'hb4efb814;
    11'b00100100010: data <= 32'h390e3298;
    11'b00100100011: data <= 32'h3a93af20;
    11'b00100100100: data <= 32'h3b1cbec0;
    11'b00100100101: data <= 32'h3d2fc0c4;
    11'b00100100110: data <= 32'h3ccabb02;
    11'b00100100111: data <= 32'h21633c9b;
    11'b00100101000: data <= 32'hbcb73d24;
    11'b00100101001: data <= 32'hbc8ab4d4;
    11'b00100101010: data <= 32'hb83cbd99;
    11'b00100101011: data <= 32'hbafcbc19;
    11'b00100101100: data <= 32'hbf60b530;
    11'b00100101101: data <= 32'hbe16b35f;
    11'b00100101110: data <= 32'h377cab34;
    11'b00100101111: data <= 32'h3f943af0;
    11'b00100110000: data <= 32'h3ba23ed2;
    11'b00100110001: data <= 32'hbc483dd9;
    11'b00100110010: data <= 32'hbe6b39f8;
    11'b00100110011: data <= 32'hb51439b9;
    11'b00100110100: data <= 32'h3abb3b98;
    11'b00100110101: data <= 32'h3a452d61;
    11'b00100110110: data <= 32'h386dbe44;
    11'b00100110111: data <= 32'h3c83bfa5;
    11'b00100111000: data <= 32'h3edab19d;
    11'b00100111001: data <= 32'h3ce73e39;
    11'b00100111010: data <= 32'h31953c4e;
    11'b00100111011: data <= 32'hb4debaeb;
    11'b00100111100: data <= 32'hb652bf24;
    11'b00100111101: data <= 32'hbc19bc2a;
    11'b00100111110: data <= 32'hbf16b58b;
    11'b00100111111: data <= 32'hbcb6ba53;
    11'b00101000000: data <= 32'h391dbcf8;
    11'b00101000001: data <= 32'h3dfcb6dd;
    11'b00101000010: data <= 32'h2fd33bc9;
    11'b00101000011: data <= 32'hbf2a3e21;
    11'b00101000100: data <= 32'hbf7d3cff;
    11'b00101000101: data <= 32'hb6213c5b;
    11'b00101000110: data <= 32'h36cd3c03;
    11'b00101000111: data <= 32'hb1f530c7;
    11'b00101001000: data <= 32'hb843bc40;
    11'b00101001001: data <= 32'h38efbbd5;
    11'b00101001010: data <= 32'h40243998;
    11'b00101001011: data <= 32'h40353fb9;
    11'b00101001100: data <= 32'h3b9e3c36;
    11'b00101001101: data <= 32'h2ca8ba03;
    11'b00101001110: data <= 32'hb1c7bcc9;
    11'b00101001111: data <= 32'hb857b468;
    11'b00101010000: data <= 32'hbb6bad7f;
    11'b00101010001: data <= 32'hb5d1bda5;
    11'b00101010010: data <= 32'h3ba2c0de;
    11'b00101010011: data <= 32'h3d25be08;
    11'b00101010100: data <= 32'hb07d36b2;
    11'b00101010101: data <= 32'hbea73d52;
    11'b00101010110: data <= 32'hbde63b92;
    11'b00101010111: data <= 32'hb55137f3;
    11'b00101011000: data <= 32'hb54f36b6;
    11'b00101011001: data <= 32'hbe2527e8;
    11'b00101011010: data <= 32'hbf0eb8eb;
    11'b00101011011: data <= 32'h290bb5ce;
    11'b00101011100: data <= 32'h401a3bec;
    11'b00101011101: data <= 32'h40473f71;
    11'b00101011110: data <= 32'h39db3c7e;
    11'b00101011111: data <= 32'hb252a7f8;
    11'b00101100000: data <= 32'hab4a2e2d;
    11'b00101100001: data <= 32'h302d3b61;
    11'b00101100010: data <= 32'haa543624;
    11'b00101100011: data <= 32'h32afbeb9;
    11'b00101100100: data <= 32'h3c4ec1d0;
    11'b00101100101: data <= 32'h3d66bee6;
    11'b00101100110: data <= 32'h361f3612;
    11'b00101100111: data <= 32'hb9093c1e;
    11'b00101101000: data <= 32'hb7d630e1;
    11'b00101101001: data <= 32'habf2b806;
    11'b00101101010: data <= 32'hbb3cb421;
    11'b00101101011: data <= 32'hc0e1aea2;
    11'b00101101100: data <= 32'hc0cdb830;
    11'b00101101101: data <= 32'hb3ccb887;
    11'b00101101110: data <= 32'h3eda3571;
    11'b00101101111: data <= 32'h3da03ccc;
    11'b00101110000: data <= 32'hb2c03c5e;
    11'b00101110001: data <= 32'hba8b3a3f;
    11'b00101110010: data <= 32'haaa83d3c;
    11'b00101110011: data <= 32'h38013f75;
    11'b00101110100: data <= 32'h30753a67;
    11'b00101110101: data <= 32'ha821bdd4;
    11'b00101110110: data <= 32'h39eac0e0;
    11'b00101110111: data <= 32'h3e12bc1e;
    11'b00101111000: data <= 32'h3d463a84;
    11'b00101111001: data <= 32'h39a73a88;
    11'b00101111010: data <= 32'h3884b847;
    11'b00101111011: data <= 32'h3572bc5a;
    11'b00101111100: data <= 32'hbb5ab606;
    11'b00101111101: data <= 32'hc0c021d8;
    11'b00101111110: data <= 32'hc034ba13;
    11'b00101111111: data <= 32'hace7bde2;
    11'b00110000000: data <= 32'h3d3bbb73;
    11'b00110000001: data <= 32'h37ac3359;
    11'b00110000010: data <= 32'hbc693ad6;
    11'b00110000011: data <= 32'hbcc43c75;
    11'b00110000100: data <= 32'ha31a3ec9;
    11'b00110000101: data <= 32'h36084002;
    11'b00110000110: data <= 32'hb8723b51;
    11'b00110000111: data <= 32'hbc55bb7d;
    11'b00110001000: data <= 32'ha299bdbc;
    11'b00110001001: data <= 32'h3e29a1c1;
    11'b00110001010: data <= 32'h3ffe3d2e;
    11'b00110001011: data <= 32'h3e0339c1;
    11'b00110001100: data <= 32'h3c4cb970;
    11'b00110001101: data <= 32'h393fba1c;
    11'b00110001110: data <= 32'hb6683575;
    11'b00110001111: data <= 32'hbdee3807;
    11'b00110010000: data <= 32'hbcb2bc20;
    11'b00110010001: data <= 32'h3569c0e2;
    11'b00110010010: data <= 32'h3c33c010;
    11'b00110010011: data <= 32'ha04cb800;
    11'b00110010100: data <= 32'hbcea37ef;
    11'b00110010101: data <= 32'hbadd39fd;
    11'b00110010110: data <= 32'h33f93c4c;
    11'b00110010111: data <= 32'ha81c3d64;
    11'b00110011000: data <= 32'hbeb039b3;
    11'b00110011001: data <= 32'hc0acb75a;
    11'b00110011010: data <= 32'hba65b8fe;
    11'b00110011011: data <= 32'h3d3e382f;
    11'b00110011100: data <= 32'h3fc23d3a;
    11'b00110011101: data <= 32'h3d1638d4;
    11'b00110011110: data <= 32'h3a35b4c3;
    11'b00110011111: data <= 32'h39ce3498;
    11'b00110100000: data <= 32'h34a73e3d;
    11'b00110100001: data <= 32'hb70e3cd5;
    11'b00110100010: data <= 32'hb5f5bc31;
    11'b00110100011: data <= 32'h387dc198;
    11'b00110100100: data <= 32'h3badc082;
    11'b00110100101: data <= 32'h3224b87d;
    11'b00110100110: data <= 32'hb71832a4;
    11'b00110100111: data <= 32'h3084ac25;
    11'b00110101000: data <= 32'h3a28abb4;
    11'b00110101001: data <= 32'hb515375e;
    11'b00110101010: data <= 32'hc0de376b;
    11'b00110101011: data <= 32'hc1feb3ec;
    11'b00110101100: data <= 32'hbca0b834;
    11'b00110101101: data <= 32'h3b7e3013;
    11'b00110101110: data <= 32'h3cb5392d;
    11'b00110101111: data <= 32'h33053518;
    11'b00110110000: data <= 32'ha6d83282;
    11'b00110110001: data <= 32'h38e73d5c;
    11'b00110110010: data <= 32'h3a024114;
    11'b00110110011: data <= 32'h26973efe;
    11'b00110110100: data <= 32'hb5a6b9e6;
    11'b00110110101: data <= 32'h33e7c08f;
    11'b00110110110: data <= 32'h3b0fbde7;
    11'b00110110111: data <= 32'h3a6a2578;
    11'b00110111000: data <= 32'h39bc2e9c;
    11'b00110111001: data <= 32'h3cfeba8e;
    11'b00110111010: data <= 32'h3d5fbb30;
    11'b00110111011: data <= 32'hb23e2d18;
    11'b00110111100: data <= 32'hc09d383a;
    11'b00110111101: data <= 32'hc147b428;
    11'b00110111110: data <= 32'hbb12bc65;
    11'b00110111111: data <= 32'h38f5bb9f;
    11'b00111000000: data <= 32'h3247b61b;
    11'b00111000001: data <= 32'hbb38b028;
    11'b00111000010: data <= 32'hb94935a5;
    11'b00111000011: data <= 32'h389a3e9b;
    11'b00111000100: data <= 32'h3a96414f;
    11'b00111000101: data <= 32'hb5773f3a;
    11'b00111000110: data <= 32'hbcc9b466;
    11'b00111000111: data <= 32'hb87abcea;
    11'b00111001000: data <= 32'h3955b400;
    11'b00111001001: data <= 32'h3d063a0b;
    11'b00111001010: data <= 32'h3db12e88;
    11'b00111001011: data <= 32'h3f0ebc87;
    11'b00111001100: data <= 32'h3ea3bb25;
    11'b00111001101: data <= 32'h34d83897;
    11'b00111001110: data <= 32'hbd793c3e;
    11'b00111001111: data <= 32'hbe1fb47e;
    11'b00111010000: data <= 32'hb35ebf41;
    11'b00111010001: data <= 32'h3789bfcb;
    11'b00111010010: data <= 32'hb6f4bc96;
    11'b00111010011: data <= 32'hbd59b864;
    11'b00111010100: data <= 32'hb886a8bf;
    11'b00111010101: data <= 32'h3adc3bdc;
    11'b00111010110: data <= 32'h39533f63;
    11'b00111010111: data <= 32'hbcb63d90;
    11'b00111011000: data <= 32'hc0a92db0;
    11'b00111011001: data <= 32'hbd9eb4c0;
    11'b00111011010: data <= 32'h352538ad;
    11'b00111011011: data <= 32'h3c813c16;
    11'b00111011100: data <= 32'h3c909fec;
    11'b00111011101: data <= 32'h3d68bbf1;
    11'b00111011110: data <= 32'h3e36b05b;
    11'b00111011111: data <= 32'h3b1c3ea2;
    11'b00111100000: data <= 32'hb31f3f5b;
    11'b00111100001: data <= 32'hb709b052;
    11'b00111100010: data <= 32'h3430c01a;
    11'b00111100011: data <= 32'h36a3c03b;
    11'b00111100100: data <= 32'hb766bc89;
    11'b00111100101: data <= 32'hbadab9af;
    11'b00111100110: data <= 32'h3482ba1e;
    11'b00111100111: data <= 32'h3dd4b3c1;
    11'b00111101000: data <= 32'h389d3980;
    11'b00111101001: data <= 32'hbf243aeb;
    11'b00111101010: data <= 32'hc1dc33a6;
    11'b00111101011: data <= 32'hbee92240;
    11'b00111101100: data <= 32'h24923806;
    11'b00111101101: data <= 32'h36b63847;
    11'b00111101110: data <= 32'h209db5e1;
    11'b00111101111: data <= 32'h34ceb9b5;
    11'b00111110000: data <= 32'h3caa39d8;
    11'b00111110001: data <= 32'h3d0f4126;
    11'b00111110010: data <= 32'h36f640c4;
    11'b00111110011: data <= 32'hae4b3133;
    11'b00111110100: data <= 32'h30bfbe38;
    11'b00111110101: data <= 32'h3472bd0d;
    11'b00111110110: data <= 32'hadbab555;
    11'b00111110111: data <= 32'h2dbdb876;
    11'b00111111000: data <= 32'h3d49bdb2;
    11'b00111111001: data <= 32'h4024bd03;
    11'b00111111010: data <= 32'h39efa4f9;
    11'b00111111011: data <= 32'hbe93399b;
    11'b00111111100: data <= 32'hc1033430;
    11'b00111111101: data <= 32'hbd17b51b;
    11'b00111111110: data <= 32'hac89b563;
    11'b00111111111: data <= 32'hb779b6a8;
    11'b01000000000: data <= 32'hbd14bb14;
    11'b01000000001: data <= 32'hb945b943;
    11'b01000000010: data <= 32'h3aff3bf0;
    11'b01000000011: data <= 32'h3d604144;
    11'b01000000100: data <= 32'h34ea409b;
    11'b01000000101: data <= 32'hb96c36f9;
    11'b01000000110: data <= 32'hb87eb8b4;
    11'b01000000111: data <= 32'ha61f2ee4;
    11'b01000001000: data <= 32'h333839c2;
    11'b01000001001: data <= 32'h39b5b498;
    11'b01000001010: data <= 32'h3f2abedd;
    11'b01000001011: data <= 32'h4097bdeb;
    11'b01000001100: data <= 32'h3c643212;
    11'b01000001101: data <= 32'hba2e3c71;
    11'b01000001110: data <= 32'hbd0f3546;
    11'b01000001111: data <= 32'hb500bae0;
    11'b01000010000: data <= 32'h2bb2bcdf;
    11'b01000010001: data <= 32'hbc39bc94;
    11'b01000010010: data <= 32'hbfb7bd0c;
    11'b01000010011: data <= 32'hbaf3bbad;
    11'b01000010100: data <= 32'h3c0435f2;
    11'b01000010101: data <= 32'h3d103ed5;
    11'b01000010110: data <= 32'hb54f3e68;
    11'b01000010111: data <= 32'hbeab382e;
    11'b01000011000: data <= 32'hbd7e349b;
    11'b01000011001: data <= 32'hb5f63ca4;
    11'b01000011010: data <= 32'h301d3d3d;
    11'b01000011011: data <= 32'h374db2cb;
    11'b01000011100: data <= 32'h3d20be90;
    11'b01000011101: data <= 32'h3fc1bb7b;
    11'b01000011110: data <= 32'h3daf3c67;
    11'b01000011111: data <= 32'h34f13f66;
    11'b01000100000: data <= 32'h28d0381f;
    11'b01000100001: data <= 32'h3828bc4e;
    11'b01000100010: data <= 32'h330dbd8a;
    11'b01000100011: data <= 32'hbc83bc39;
    11'b01000100100: data <= 32'hbeb0bcdf;
    11'b01000100101: data <= 32'hb31ebdd0;
    11'b01000100110: data <= 32'h3e36ba4d;
    11'b01000100111: data <= 32'h3cf7358c;
    11'b01000101000: data <= 32'hbafd39cf;
    11'b01000101001: data <= 32'hc07b36d5;
    11'b01000101010: data <= 32'hbe9038f8;
    11'b01000101011: data <= 32'hb82b3d40;
    11'b01000101100: data <= 32'hb6273c38;
    11'b01000101101: data <= 32'hb8ecb804;
    11'b01000101110: data <= 32'h2979bdc3;
    11'b01000101111: data <= 32'h3cd0b17a;
    11'b01000110000: data <= 32'h3e213fe1;
    11'b01000110001: data <= 32'h3bc440b7;
    11'b01000110010: data <= 32'h38f839ab;
    11'b01000110011: data <= 32'h3962b9d4;
    11'b01000110100: data <= 32'h31d4b8a8;
    11'b01000110101: data <= 32'hbab6ad81;
    11'b01000110110: data <= 32'hbae1b9db;
    11'b01000110111: data <= 32'h39f6bf5b;
    11'b01000111000: data <= 32'h404abf25;
    11'b01000111001: data <= 32'h3d67b8dd;
    11'b01000111010: data <= 32'hbaab342a;
    11'b01000111011: data <= 32'hbf6d350d;
    11'b01000111100: data <= 32'hbc2835ea;
    11'b01000111101: data <= 32'hb4e03915;
    11'b01000111110: data <= 32'hbc033281;
    11'b01000111111: data <= 32'hbf7cbc05;
    11'b01001000000: data <= 32'hbcaabd7d;
    11'b01001000001: data <= 32'h38a630bb;
    11'b01001000010: data <= 32'h3dc1401c;
    11'b01001000011: data <= 32'h3b4b4050;
    11'b01001000100: data <= 32'h336239b6;
    11'b01001000101: data <= 32'h2e12a21c;
    11'b01001000110: data <= 32'hae9d3a18;
    11'b01001000111: data <= 32'hb8613cdb;
    11'b01001001000: data <= 32'hb311af18;
    11'b01001001001: data <= 32'h3cefbfb4;
    11'b01001001010: data <= 32'h4090c022;
    11'b01001001011: data <= 32'h3defb8e1;
    11'b01001001100: data <= 32'hb1ff37fc;
    11'b01001001101: data <= 32'hb92335a3;
    11'b01001001110: data <= 32'h312aafcb;
    11'b01001001111: data <= 32'h31fdb316;
    11'b01001010000: data <= 32'hbd73b842;
    11'b01001010001: data <= 32'hc125bd4e;
    11'b01001010010: data <= 32'hbe6ebe00;
    11'b01001010011: data <= 32'h37f9b473;
    11'b01001010100: data <= 32'h3d373ca3;
    11'b01001010101: data <= 32'h355f3ceb;
    11'b01001010110: data <= 32'hb993370e;
    11'b01001010111: data <= 32'hb9a538f5;
    11'b01001011000: data <= 32'hb6c13f64;
    11'b01001011001: data <= 32'hb82d401c;
    11'b01001011010: data <= 32'hb51632fa;
    11'b01001011011: data <= 32'h3a0dbf0c;
    11'b01001011100: data <= 32'h3ee3be5e;
    11'b01001011101: data <= 32'h3dd83291;
    11'b01001011110: data <= 32'h39283cd0;
    11'b01001011111: data <= 32'h39833832;
    11'b01001100000: data <= 32'h3d0cb69f;
    11'b01001100001: data <= 32'h3920b816;
    11'b01001100010: data <= 32'hbd41b7a9;
    11'b01001100011: data <= 32'hc0c6bc73;
    11'b01001100100: data <= 32'hbc5bbeb4;
    11'b01001100101: data <= 32'h3bdabcc3;
    11'b01001100110: data <= 32'h3d16b32f;
    11'b01001100111: data <= 32'hb3c32cb4;
    11'b01001101000: data <= 32'hbd6e2498;
    11'b01001101001: data <= 32'hbc0a3a68;
    11'b01001101010: data <= 32'hb7064024;
    11'b01001101011: data <= 32'hba0d3fdb;
    11'b01001101100: data <= 32'hbc9f27d4;
    11'b01001101101: data <= 32'hb7f3be30;
    11'b01001101110: data <= 32'h39a3ba91;
    11'b01001101111: data <= 32'h3ce03c82;
    11'b01001110000: data <= 32'h3c813efd;
    11'b01001110001: data <= 32'h3d6138fb;
    11'b01001110010: data <= 32'h3e75b4ce;
    11'b01001110011: data <= 32'h39fb2ce1;
    11'b01001110100: data <= 32'hbbfa37ef;
    11'b01001110101: data <= 32'hbe5db5af;
    11'b01001110110: data <= 32'hae80beca;
    11'b01001110111: data <= 32'h3e69bff3;
    11'b01001111000: data <= 32'h3d44bd01;
    11'b01001111001: data <= 32'hb646b904;
    11'b01001111010: data <= 32'hbcaab498;
    11'b01001111011: data <= 32'hb6a237ff;
    11'b01001111100: data <= 32'h271d3db8;
    11'b01001111101: data <= 32'hbc0f3c81;
    11'b01001111110: data <= 32'hc065b7d9;
    11'b01001111111: data <= 32'hbf1abdc3;
    11'b01010000000: data <= 32'hb1e0b5a8;
    11'b01010000001: data <= 32'h3b103d89;
    11'b01010000010: data <= 32'h3bec3e41;
    11'b01010000011: data <= 32'h3c063681;
    11'b01010000100: data <= 32'h3c5e2cc3;
    11'b01010000101: data <= 32'h377a3ccf;
    11'b01010000110: data <= 32'hb9793f74;
    11'b01010000111: data <= 32'hbabb386f;
    11'b01010001000: data <= 32'h3849bdff;
    11'b01010001001: data <= 32'h3f16c053;
    11'b01010001010: data <= 32'h3d0dbd47;
    11'b01010001011: data <= 32'habfcb7d2;
    11'b01010001100: data <= 32'hb157b4a4;
    11'b01010001101: data <= 32'h3aca9e31;
    11'b01010001110: data <= 32'h3a8f37f9;
    11'b01010001111: data <= 32'hbc3b3440;
    11'b01010010000: data <= 32'hc189bada;
    11'b01010010001: data <= 32'hc097bdaf;
    11'b01010010010: data <= 32'hb69cb7e6;
    11'b01010010011: data <= 32'h39513995;
    11'b01010010100: data <= 32'h365138ab;
    11'b01010010101: data <= 32'h2883b162;
    11'b01010010110: data <= 32'h323e35e6;
    11'b01010010111: data <= 32'h2e274047;
    11'b01010011000: data <= 32'hb8644196;
    11'b01010011001: data <= 32'hb97f3c4c;
    11'b01010011010: data <= 32'h3439bcd0;
    11'b01010011011: data <= 32'h3cb3be9d;
    11'b01010011100: data <= 32'h3b98b7cb;
    11'b01010011101: data <= 32'h36c4346e;
    11'b01010011110: data <= 32'h3c02ac6d;
    11'b01010011111: data <= 32'h4019b601;
    11'b01010100000: data <= 32'h3e079e5b;
    11'b01010100001: data <= 32'hbaa32fb2;
    11'b01010100010: data <= 32'hc10fb907;
    11'b01010100011: data <= 32'hbf23bd50;
    11'b01010100100: data <= 32'h2dd6bc3e;
    11'b01010100101: data <= 32'h3952b81d;
    11'b01010100110: data <= 32'hb39fb972;
    11'b01010100111: data <= 32'hba72bae5;
    11'b01010101000: data <= 32'hb4c53538;
    11'b01010101001: data <= 32'h2c644097;
    11'b01010101010: data <= 32'hb8604178;
    11'b01010101011: data <= 32'hbcc23b4b;
    11'b01010101100: data <= 32'hba78bbf7;
    11'b01010101101: data <= 32'h2a67bab9;
    11'b01010101110: data <= 32'h368b38a9;
    11'b01010101111: data <= 32'h39223bf6;
    11'b01010110000: data <= 32'h3e4d2bcc;
    11'b01010110001: data <= 32'h40edb75f;
    11'b01010110010: data <= 32'h3ec23441;
    11'b01010110011: data <= 32'hb7c13b42;
    11'b01010110100: data <= 32'hbec9333e;
    11'b01010110101: data <= 32'hb96cbc27;
    11'b01010110110: data <= 32'h3af4be41;
    11'b01010110111: data <= 32'h3a0ebdc7;
    11'b01010111000: data <= 32'hb869bde1;
    11'b01010111001: data <= 32'hbb3ebd30;
    11'b01010111010: data <= 32'h2ea4a9aa;
    11'b01010111011: data <= 32'h38eb3e77;
    11'b01010111100: data <= 32'hb7f23f3d;
    11'b01010111101: data <= 32'hbfac3424;
    11'b01010111110: data <= 32'hbfe9bb8b;
    11'b01010111111: data <= 32'hbb9ab3af;
    11'b01011000000: data <= 32'haf283c6e;
    11'b01011000001: data <= 32'h36413c0b;
    11'b01011000010: data <= 32'h3cc9b2c1;
    11'b01011000011: data <= 32'h3f8cb61b;
    11'b01011000100: data <= 32'h3d3f3c48;
    11'b01011000101: data <= 32'hb321404e;
    11'b01011000110: data <= 32'hbab73d0e;
    11'b01011000111: data <= 32'h3293b8dd;
    11'b01011001000: data <= 32'h3cf6be50;
    11'b01011001001: data <= 32'h3964bddd;
    11'b01011001010: data <= 32'hb7ecbd44;
    11'b01011001011: data <= 32'hb34ebcfe;
    11'b01011001100: data <= 32'h3cf1b81b;
    11'b01011001101: data <= 32'h3e2b38c6;
    11'b01011001110: data <= 32'hb45739d1;
    11'b01011001111: data <= 32'hc093b4ff;
    11'b01011010000: data <= 32'hc0e3bb5e;
    11'b01011010001: data <= 32'hbcd0b03e;
    11'b01011010010: data <= 32'hb55139eb;
    11'b01011010011: data <= 32'hb239318e;
    11'b01011010100: data <= 32'h30e3bb5a;
    11'b01011010101: data <= 32'h3a5eb60c;
    11'b01011010110: data <= 32'h39eb3f19;
    11'b01011010111: data <= 32'haf17420d;
    11'b01011011000: data <= 32'hb7733f61;
    11'b01011011001: data <= 32'h33e2b407;
    11'b01011011010: data <= 32'h3a6dbc2d;
    11'b01011011011: data <= 32'h339cb891;
    11'b01011011100: data <= 32'hb500b63e;
    11'b01011011101: data <= 32'h397ababe;
    11'b01011011110: data <= 32'h40bfbabd;
    11'b01011011111: data <= 32'h40a6ae4c;
    11'b01011100000: data <= 32'h2cb2346b;
    11'b01011100001: data <= 32'hbff2b436;
    11'b01011100010: data <= 32'hbf82b9d0;
    11'b01011100011: data <= 32'hb89bb655;
    11'b01011100100: data <= 32'hb1a6b256;
    11'b01011100101: data <= 32'hba40bc18;
    11'b01011100110: data <= 32'hbad3bef4;
    11'b01011100111: data <= 32'h2092b8b7;
    11'b01011101000: data <= 32'h381e3f52;
    11'b01011101001: data <= 32'ha8ab41d5;
    11'b01011101010: data <= 32'hb9633e66;
    11'b01011101011: data <= 32'hb84cb120;
    11'b01011101100: data <= 32'hb3d3b450;
    11'b01011101101: data <= 32'hb72d3924;
    11'b01011101110: data <= 32'hb4eb38da;
    11'b01011101111: data <= 32'h3c7fb803;
    11'b01011110000: data <= 32'h417dbbc1;
    11'b01011110001: data <= 32'h40f1aeb8;
    11'b01011110010: data <= 32'h35983a1a;
    11'b01011110011: data <= 32'hbcb437f5;
    11'b01011110100: data <= 32'hb925b484;
    11'b01011110101: data <= 32'h3761b930;
    11'b01011110110: data <= 32'h3035bbb6;
    11'b01011110111: data <= 32'hbc6fbf1e;
    11'b01011111000: data <= 32'hbcd8c05f;
    11'b01011111001: data <= 32'h2e96bb8e;
    11'b01011111010: data <= 32'h3b8d3c9d;
    11'b01011111011: data <= 32'h31363f84;
    11'b01011111100: data <= 32'hbc8239b5;
    11'b01011111101: data <= 32'hbe0fb518;
    11'b01011111110: data <= 32'hbcdf3537;
    11'b01011111111: data <= 32'hbc1e3da1;
    11'b01100000000: data <= 32'hb8cd3b7b;
    11'b01100000001: data <= 32'h39c6b90e;
    11'b01100000010: data <= 32'h4026bc17;
    11'b01100000011: data <= 32'h3f92369f;
    11'b01100000100: data <= 32'h36a73f2c;
    11'b01100000101: data <= 32'hb55d3e07;
    11'b01100000110: data <= 32'h376c33fb;
    11'b01100000111: data <= 32'h3c99b885;
    11'b01100001000: data <= 32'h32e3bb7c;
    11'b01100001001: data <= 32'hbca7be36;
    11'b01100001010: data <= 32'hba94bfed;
    11'b01100001011: data <= 32'h3bfcbcfb;
    11'b01100001100: data <= 32'h3f5930ec;
    11'b01100001101: data <= 32'h382738b5;
    11'b01100001110: data <= 32'hbd65b19f;
    11'b01100001111: data <= 32'hbf9cb7cb;
    11'b01100010000: data <= 32'hbdad3828;
    11'b01100010001: data <= 32'hbc963d4e;
    11'b01100010010: data <= 32'hbc3a35ab;
    11'b01100010011: data <= 32'hb4dfbd2c;
    11'b01100010100: data <= 32'h3a5dbcab;
    11'b01100010101: data <= 32'h3c093b72;
    11'b01100010110: data <= 32'h351a411f;
    11'b01100010111: data <= 32'h2e6f401d;
    11'b01100011000: data <= 32'h3a4f3875;
    11'b01100011001: data <= 32'h3beaaf0a;
    11'b01100011010: data <= 32'hb0efaa08;
    11'b01100011011: data <= 32'hbc8ab758;
    11'b01100011100: data <= 32'hb010bd20;
    11'b01100011101: data <= 32'h4005bd6d;
    11'b01100011110: data <= 32'h4135b8a7;
    11'b01100011111: data <= 32'h3af1b085;
    11'b01100100000: data <= 32'hbc4cb6cf;
    11'b01100100001: data <= 32'hbd4fb62f;
    11'b01100100010: data <= 32'hb92e3686;
    11'b01100100011: data <= 32'hb9d23908;
    11'b01100100100: data <= 32'hbdbab991;
    11'b01100100101: data <= 32'hbd56c037;
    11'b01100100110: data <= 32'hb435bdb8;
    11'b01100100111: data <= 32'h37703bb4;
    11'b01100101000: data <= 32'h344640db;
    11'b01100101001: data <= 32'h28253ec6;
    11'b01100101010: data <= 32'h343a36ce;
    11'b01100101011: data <= 32'h2f2c3788;
    11'b01100101100: data <= 32'hbaba3cba;
    11'b01100101101: data <= 32'hbce23a63;
    11'b01100101110: data <= 32'h33c6b8dc;
    11'b01100101111: data <= 32'h40b0bd4d;
    11'b01100110000: data <= 32'h4152b9ad;
    11'b01100110001: data <= 32'h3bc02c94;
    11'b01100110010: data <= 32'hb6d93056;
    11'b01100110011: data <= 32'had252a9e;
    11'b01100110100: data <= 32'h3918346c;
    11'b01100110101: data <= 32'had45a699;
    11'b01100110110: data <= 32'hbe4ebd9b;
    11'b01100110111: data <= 32'hbf2dc0ff;
    11'b01100111000: data <= 32'hb740bea6;
    11'b01100111001: data <= 32'h394d369d;
    11'b01100111010: data <= 32'h37143d81;
    11'b01100111011: data <= 32'hb482389e;
    11'b01100111100: data <= 32'hb884ac0f;
    11'b01100111101: data <= 32'hba5f3af4;
    11'b01100111110: data <= 32'hbd964010;
    11'b01100111111: data <= 32'hbdca3dac;
    11'b01101000000: data <= 32'hac8bb797;
    11'b01101000001: data <= 32'h3ea3bd4f;
    11'b01101000010: data <= 32'h3f82b564;
    11'b01101000011: data <= 32'h39c63b5f;
    11'b01101000100: data <= 32'h32c83c3f;
    11'b01101000101: data <= 32'h3c6638a7;
    11'b01101000110: data <= 32'h3e7d3591;
    11'b01101000111: data <= 32'h34b6a987;
    11'b01101001000: data <= 32'hbe32bca3;
    11'b01101001001: data <= 32'hbe32c03d;
    11'b01101001010: data <= 32'h3380beb8;
    11'b01101001011: data <= 32'h3dcab63f;
    11'b01101001100: data <= 32'h3a7a2539;
    11'b01101001101: data <= 32'hb77db8e9;
    11'b01101001110: data <= 32'hbba6b869;
    11'b01101001111: data <= 32'hbbda3b9c;
    11'b01101010000: data <= 32'hbd84402d;
    11'b01101010001: data <= 32'hbea73c47;
    11'b01101010010: data <= 32'hbb55bbfd;
    11'b01101010011: data <= 32'h3522bdef;
    11'b01101010100: data <= 32'h398e2ef8;
    11'b01101010101: data <= 32'h34933e9d;
    11'b01101010110: data <= 32'h38133e5d;
    11'b01101010111: data <= 32'h3e3a3a5c;
    11'b01101011000: data <= 32'h3ee038e7;
    11'b01101011001: data <= 32'h2e1e3981;
    11'b01101011010: data <= 32'hbe18a426;
    11'b01101011011: data <= 32'hbb99bc89;
    11'b01101011100: data <= 32'h3cb4bdc6;
    11'b01101011101: data <= 32'h4060bbba;
    11'b01101011110: data <= 32'h3c67bab0;
    11'b01101011111: data <= 32'hb547bc95;
    11'b01101100000: data <= 32'hb810b946;
    11'b01101100001: data <= 32'hb16c3a99;
    11'b01101100010: data <= 32'hb9903e06;
    11'b01101100011: data <= 32'hbec92fd9;
    11'b01101100100: data <= 32'hbf17bf1d;
    11'b01101100101: data <= 32'hbaddbee1;
    11'b01101100110: data <= 32'hb0f83339;
    11'b01101100111: data <= 32'ha3bd3e76;
    11'b01101101000: data <= 32'h36723cc9;
    11'b01101101001: data <= 32'h3ca436e9;
    11'b01101101010: data <= 32'h3bd43afe;
    11'b01101101011: data <= 32'hb8543ef6;
    11'b01101101100: data <= 32'hbe6d3d6b;
    11'b01101101101: data <= 32'hb854b06d;
    11'b01101101110: data <= 32'h3e4cbc80;
    11'b01101101111: data <= 32'h4073bc1c;
    11'b01101110000: data <= 32'h3c08ba16;
    11'b01101110001: data <= 32'h27a9ba0f;
    11'b01101110010: data <= 32'h388db4ba;
    11'b01101110011: data <= 32'h3ce239a3;
    11'b01101110100: data <= 32'h34733ad1;
    11'b01101110101: data <= 32'hbe19b8f6;
    11'b01101110110: data <= 32'hc047c051;
    11'b01101110111: data <= 32'hbcc4bf34;
    11'b01101111000: data <= 32'hb167ace5;
    11'b01101111001: data <= 32'h2a7339c4;
    11'b01101111010: data <= 32'h2e82a46d;
    11'b01101111011: data <= 32'h35e5b61f;
    11'b01101111100: data <= 32'h2c003b81;
    11'b01101111101: data <= 32'hbc6140f3;
    11'b01101111110: data <= 32'hbee6403e;
    11'b01101111111: data <= 32'hb93533ce;
    11'b01110000000: data <= 32'h3c21bbcd;
    11'b01110000001: data <= 32'h3d6cb945;
    11'b01110000010: data <= 32'h372f2609;
    11'b01110000011: data <= 32'h354b3092;
    11'b01110000100: data <= 32'h3e7c3382;
    11'b01110000101: data <= 32'h40b739ab;
    11'b01110000110: data <= 32'h3b813969;
    11'b01110000111: data <= 32'hbd35b80d;
    11'b01110001000: data <= 32'hbf85beda;
    11'b01110001001: data <= 32'hb8bdbe1f;
    11'b01110001010: data <= 32'h386db862;
    11'b01110001011: data <= 32'h368ab7fe;
    11'b01110001100: data <= 32'hafa8bd74;
    11'b01110001101: data <= 32'hb063bcbb;
    11'b01110001110: data <= 32'hb3813a46;
    11'b01110001111: data <= 32'hbc2140ff;
    11'b01110010000: data <= 32'hbec13f86;
    11'b01110010001: data <= 32'hbcbab1b0;
    11'b01110010010: data <= 32'hb159bc68;
    11'b01110010011: data <= 32'h2439b25a;
    11'b01110010100: data <= 32'hb5263aa0;
    11'b01110010101: data <= 32'h35b53a1f;
    11'b01110010110: data <= 32'h400e36d1;
    11'b01110010111: data <= 32'h412a3a1d;
    11'b01110011000: data <= 32'h3b143c7a;
    11'b01110011001: data <= 32'hbcdf37f7;
    11'b01110011010: data <= 32'hbd1bb8a1;
    11'b01110011011: data <= 32'h362fbb95;
    11'b01110011100: data <= 32'h3d75ba98;
    11'b01110011101: data <= 32'h3991bd2a;
    11'b01110011110: data <= 32'hb0a9c017;
    11'b01110011111: data <= 32'h2b5dbdee;
    11'b01110100000: data <= 32'h37083882;
    11'b01110100001: data <= 32'hb2f43fa8;
    11'b01110100010: data <= 32'hbd833b6e;
    11'b01110100011: data <= 32'hbee2bc02;
    11'b01110100100: data <= 32'hbd12bd61;
    11'b01110100101: data <= 32'hbc02295b;
    11'b01110100110: data <= 32'hbae63c07;
    11'b01110100111: data <= 32'h2f63380b;
    11'b01110101000: data <= 32'h3e81a9f7;
    11'b01110101001: data <= 32'h3f793998;
    11'b01110101010: data <= 32'h337b3f66;
    11'b01110101011: data <= 32'hbd3c3f1f;
    11'b01110101100: data <= 32'hba3a38cd;
    11'b01110101101: data <= 32'h3bbeb586;
    11'b01110101110: data <= 32'h3e20b9a9;
    11'b01110101111: data <= 32'h3829bcd1;
    11'b01110110000: data <= 32'had54bedd;
    11'b01110110001: data <= 32'h3a8fbc93;
    11'b01110110010: data <= 32'h3eef371a;
    11'b01110110011: data <= 32'h3b913cca;
    11'b01110110100: data <= 32'hbb192885;
    11'b01110110101: data <= 32'hbf7abe09;
    11'b01110110110: data <= 32'hbe54bd7b;
    11'b01110110111: data <= 32'hbc7018ca;
    11'b01110111000: data <= 32'hbaf5369c;
    11'b01110111001: data <= 32'hb289b8db;
    11'b01110111010: data <= 32'h3a56bc31;
    11'b01110111011: data <= 32'h3aac36c9;
    11'b01110111100: data <= 32'hb70540ab;
    11'b01110111101: data <= 32'hbd98410a;
    11'b01110111110: data <= 32'hb94d3c71;
    11'b01110111111: data <= 32'h39a8ac6f;
    11'b01111000000: data <= 32'h3a28b4a5;
    11'b01111000001: data <= 32'hb2eeb646;
    11'b01111000010: data <= 32'hb024b9dc;
    11'b01111000011: data <= 32'h3e67b813;
    11'b01111000100: data <= 32'h41ac3710;
    11'b01111000101: data <= 32'h3f0e3aac;
    11'b01111000110: data <= 32'hb7bfaf37;
    11'b01111000111: data <= 32'hbe19bcb8;
    11'b01111001000: data <= 32'hbbb4bb87;
    11'b01111001001: data <= 32'hb578b007;
    11'b01111001010: data <= 32'hb6edb831;
    11'b01111001011: data <= 32'hb6b3bfa9;
    11'b01111001100: data <= 32'h3052c011;
    11'b01111001101: data <= 32'h34be2922;
    11'b01111001110: data <= 32'hb80b4078;
    11'b01111001111: data <= 32'hbcec4086;
    11'b01111010000: data <= 32'hbaeb3976;
    11'b01111010001: data <= 32'hb27db3a0;
    11'b01111010010: data <= 32'hb8343134;
    11'b01111010011: data <= 32'hbcc53843;
    11'b01111010100: data <= 32'hb6042ec9;
    11'b01111010101: data <= 32'h3f65b1be;
    11'b01111010110: data <= 32'h42193664;
    11'b01111010111: data <= 32'h3efc3bc8;
    11'b01111011000: data <= 32'hb65a38cd;
    11'b01111011001: data <= 32'hbb55ae4a;
    11'b01111011010: data <= 32'h2f32b08f;
    11'b01111011011: data <= 32'h3944ae1b;
    11'b01111011100: data <= 32'h9b3abc82;
    11'b01111011101: data <= 32'hb814c12e;
    11'b01111011110: data <= 32'h2b0ec0d3;
    11'b01111011111: data <= 32'h3975b37c;
    11'b01111100000: data <= 32'h33c13e80;
    11'b01111100001: data <= 32'hb9a83cee;
    11'b01111100010: data <= 32'hbc4cb4d0;
    11'b01111100011: data <= 32'hbc5db8f0;
    11'b01111100100: data <= 32'hbe2d3711;
    11'b01111100101: data <= 32'hbf6e3ba3;
    11'b01111100110: data <= 32'hb9cd3015;
    11'b01111100111: data <= 32'h3d97b886;
    11'b01111101000: data <= 32'h408c3064;
    11'b01111101001: data <= 32'h3bc33d75;
    11'b01111101010: data <= 32'hb8e23e99;
    11'b01111101011: data <= 32'hb6593c55;
    11'b01111101100: data <= 32'h3b423902;
    11'b01111101101: data <= 32'h3c6331e0;
    11'b01111101110: data <= 32'hacb1bbb7;
    11'b01111101111: data <= 32'hb8f5c070;
    11'b01111110000: data <= 32'h37bcbff6;
    11'b01111110001: data <= 32'h3eeab41b;
    11'b01111110010: data <= 32'h3d9f3b2c;
    11'b01111110011: data <= 32'ha4b930cf;
    11'b01111110100: data <= 32'hbc09bc47;
    11'b01111110101: data <= 32'hbd33ba22;
    11'b01111110110: data <= 32'hbe85385d;
    11'b01111110111: data <= 32'hbf523975;
    11'b01111111000: data <= 32'hbbe0b9d1;
    11'b01111111001: data <= 32'h386bbe3d;
    11'b01111111010: data <= 32'h3c4cb5b0;
    11'b01111111011: data <= 32'h2a353e60;
    11'b01111111100: data <= 32'hbab64083;
    11'b01111111101: data <= 32'hb15b3e5c;
    11'b01111111110: data <= 32'h3b9e3b5f;
    11'b01111111111: data <= 32'h38cf38b3;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    