
module memory_rom_32(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbb8ebd16;
    11'b00000000001: data <= 32'hb88cb96e;
    11'b00000000010: data <= 32'h383c3a40;
    11'b00000000011: data <= 32'h34d13f66;
    11'b00000000100: data <= 32'hbd373c88;
    11'b00000000101: data <= 32'hc09ab80a;
    11'b00000000110: data <= 32'hbe7fbad7;
    11'b00000000111: data <= 32'hb58a36e3;
    11'b00000001000: data <= 32'h35b53d3a;
    11'b00000001001: data <= 32'h3a573806;
    11'b00000001010: data <= 32'h3ddcb7ef;
    11'b00000001011: data <= 32'h3e8d3239;
    11'b00000001100: data <= 32'h38ab3f52;
    11'b00000001101: data <= 32'hb956401b;
    11'b00000001110: data <= 32'hb7bf3553;
    11'b00000001111: data <= 32'h3a56bdb7;
    11'b00000010000: data <= 32'h3cbdbf03;
    11'b00000010001: data <= 32'h3055bd25;
    11'b00000010010: data <= 32'hb855bc64;
    11'b00000010011: data <= 32'h3742bb11;
    11'b00000010100: data <= 32'h3e97a80d;
    11'b00000010101: data <= 32'h3ae639d3;
    11'b00000010110: data <= 32'hbdd53500;
    11'b00000010111: data <= 32'hc187b995;
    11'b00000011000: data <= 32'hbfc5b9bb;
    11'b00000011001: data <= 32'hb80f3480;
    11'b00000011010: data <= 32'ha75a38c4;
    11'b00000011011: data <= 32'had93b5f2;
    11'b00000011100: data <= 32'h3512bad3;
    11'b00000011101: data <= 32'h3a5e390d;
    11'b00000011110: data <= 32'h36c84161;
    11'b00000011111: data <= 32'hb5934187;
    11'b00000100000: data <= 32'hb48239d3;
    11'b00000100001: data <= 32'h37fdbc12;
    11'b00000100010: data <= 32'h3928bbdd;
    11'b00000100011: data <= 32'ha132b492;
    11'b00000100100: data <= 32'h2d5eb671;
    11'b00000100101: data <= 32'h3e48bb40;
    11'b00000100110: data <= 32'h413fb903;
    11'b00000100111: data <= 32'h3d74309f;
    11'b00000101000: data <= 32'hbcbf3232;
    11'b00000101001: data <= 32'hc098b798;
    11'b00000101010: data <= 32'hbd04b9cc;
    11'b00000101011: data <= 32'hac48b645;
    11'b00000101100: data <= 32'hb4aeb896;
    11'b00000101101: data <= 32'hbbcebdab;
    11'b00000101110: data <= 32'hb8e5bd47;
    11'b00000101111: data <= 32'h35b538ed;
    11'b00000110000: data <= 32'h3732414f;
    11'b00000110001: data <= 32'hb61b4104;
    11'b00000110010: data <= 32'hbac538b6;
    11'b00000110011: data <= 32'hb832b871;
    11'b00000110100: data <= 32'hb4672ed1;
    11'b00000110101: data <= 32'hb5073b04;
    11'b00000110110: data <= 32'h35ff330e;
    11'b00000110111: data <= 32'h3ff7bb34;
    11'b00000111000: data <= 32'h41a5b9ec;
    11'b00000111001: data <= 32'h3e0a3720;
    11'b00000111010: data <= 32'hb90d3b73;
    11'b00000111011: data <= 32'hbcbe3227;
    11'b00000111100: data <= 32'ha95eb947;
    11'b00000111101: data <= 32'h38b0bbd3;
    11'b00000111110: data <= 32'hb65fbd7a;
    11'b00000111111: data <= 32'hbd89bfeb;
    11'b00001000000: data <= 32'hb99cbea4;
    11'b00001000001: data <= 32'h39df2e82;
    11'b00001000010: data <= 32'h3abc3ee3;
    11'b00001000011: data <= 32'hb8473dd9;
    11'b00001000100: data <= 32'hbe9a2c0b;
    11'b00001000101: data <= 32'hbe39b40b;
    11'b00001000110: data <= 32'hbc1d3af0;
    11'b00001000111: data <= 32'hb9893da1;
    11'b00001001000: data <= 32'h292f32d7;
    11'b00001001001: data <= 32'h3d92bc55;
    11'b00001001010: data <= 32'h403bb7ea;
    11'b00001001011: data <= 32'h3cf13d45;
    11'b00001001100: data <= 32'haede4010;
    11'b00001001101: data <= 32'hafe53ba7;
    11'b00001001110: data <= 32'h3aecb6a1;
    11'b00001001111: data <= 32'h3b15bb9b;
    11'b00001010000: data <= 32'hb7b1bcc6;
    11'b00001010001: data <= 32'hbce3bebd;
    11'b00001010010: data <= 32'h2897bebb;
    11'b00001010011: data <= 32'h3eeab8e2;
    11'b00001010100: data <= 32'h3ded37c3;
    11'b00001010101: data <= 32'hb83f357e;
    11'b00001010110: data <= 32'hc003b665;
    11'b00001010111: data <= 32'hbf4ab0a1;
    11'b00001011000: data <= 32'hbc723b92;
    11'b00001011001: data <= 32'hbb903bf5;
    11'b00001011010: data <= 32'hba0eb825;
    11'b00001011011: data <= 32'h3091be17;
    11'b00001011100: data <= 32'h3becb3f7;
    11'b00001011101: data <= 32'h3a5f4011;
    11'b00001011110: data <= 32'h30f14161;
    11'b00001011111: data <= 32'h34b13d44;
    11'b00001100000: data <= 32'h3b11ad0e;
    11'b00001100001: data <= 32'h3817b388;
    11'b00001100010: data <= 32'hb9a0ae84;
    11'b00001100011: data <= 32'hba7db9d4;
    11'b00001100100: data <= 32'h3bd4bdb7;
    11'b00001100101: data <= 32'h414cbc83;
    11'b00001100110: data <= 32'h3ff3b4c2;
    11'b00001100111: data <= 32'hb470ae51;
    11'b00001101000: data <= 32'hbe3db5f4;
    11'b00001101001: data <= 32'hbc36add4;
    11'b00001101010: data <= 32'hb7163807;
    11'b00001101011: data <= 32'hbb9726d7;
    11'b00001101100: data <= 32'hbe3abe06;
    11'b00001101101: data <= 32'hbbc1c00f;
    11'b00001101110: data <= 32'h330bb4d2;
    11'b00001101111: data <= 32'h38c43ff2;
    11'b00001110000: data <= 32'h311b40ba;
    11'b00001110001: data <= 32'ha8513be8;
    11'b00001110010: data <= 32'h2d9730eb;
    11'b00001110011: data <= 32'hb5713a22;
    11'b00001110100: data <= 32'hbc4e3ceb;
    11'b00001110101: data <= 32'hb8d93348;
    11'b00001110110: data <= 32'h3d6dbcad;
    11'b00001110111: data <= 32'h4195bd02;
    11'b00001111000: data <= 32'h3ff4b380;
    11'b00001111001: data <= 32'h2d963626;
    11'b00001111010: data <= 32'hb83432a4;
    11'b00001111011: data <= 32'h350d2b97;
    11'b00001111100: data <= 32'h384e29e0;
    11'b00001111101: data <= 32'hba43b995;
    11'b00001111110: data <= 32'hbfcdc00d;
    11'b00001111111: data <= 32'hbd2bc08c;
    11'b00010000000: data <= 32'h3512b95f;
    11'b00010000001: data <= 32'h3afc3c76;
    11'b00010000010: data <= 32'h2e1f3cb2;
    11'b00010000011: data <= 32'hb96630b4;
    11'b00010000100: data <= 32'hbabe31a8;
    11'b00010000101: data <= 32'hbc403df8;
    11'b00010000110: data <= 32'hbda23ff5;
    11'b00010000111: data <= 32'hbac93832;
    11'b00010001000: data <= 32'h3a6cbcd1;
    11'b00010001001: data <= 32'h3fd5bc58;
    11'b00010001010: data <= 32'h3db13730;
    11'b00010001011: data <= 32'h35603d6a;
    11'b00010001100: data <= 32'h37d73b90;
    11'b00010001101: data <= 32'h3dcc34e4;
    11'b00010001110: data <= 32'h3ca62864;
    11'b00010001111: data <= 32'hb977b861;
    11'b00010010000: data <= 32'hbf69be81;
    11'b00010010001: data <= 32'hba16c014;
    11'b00010010010: data <= 32'h3c9abc7e;
    11'b00010010011: data <= 32'h3dedac5d;
    11'b00010010100: data <= 32'h305bb15f;
    11'b00010010101: data <= 32'hbc13b946;
    11'b00010010110: data <= 32'hbc742c8f;
    11'b00010010111: data <= 32'hbc443e79;
    11'b00010011000: data <= 32'hbdcd3f2f;
    11'b00010011001: data <= 32'hbda7a407;
    11'b00010011010: data <= 32'hb646be65;
    11'b00010011011: data <= 32'h38f1bb37;
    11'b00010011100: data <= 32'h39073c71;
    11'b00010011101: data <= 32'h35b23ffb;
    11'b00010011110: data <= 32'h3b7c3d00;
    11'b00010011111: data <= 32'h3ecc37b4;
    11'b00010100000: data <= 32'h3c0e3871;
    11'b00010100001: data <= 32'hbab837df;
    11'b00010100010: data <= 32'hbe10b788;
    11'b00010100011: data <= 32'h2dcfbdba;
    11'b00010100100: data <= 32'h4011bd84;
    11'b00010100101: data <= 32'h3fd0bae8;
    11'b00010100110: data <= 32'h3483bad6;
    11'b00010100111: data <= 32'hb9c7bb27;
    11'b00010101000: data <= 32'hb63e27ad;
    11'b00010101001: data <= 32'hb3063d04;
    11'b00010101010: data <= 32'hbc763b9b;
    11'b00010101011: data <= 32'hbfc6bb8a;
    11'b00010101100: data <= 32'hbe03c02d;
    11'b00010101101: data <= 32'hb682bb27;
    11'b00010101110: data <= 32'h30183cad;
    11'b00010101111: data <= 32'h33643ed3;
    11'b00010110000: data <= 32'h397c3a28;
    11'b00010110001: data <= 32'h3c39367b;
    11'b00010110010: data <= 32'h34003d2d;
    11'b00010110011: data <= 32'hbccf3f40;
    11'b00010110100: data <= 32'hbd2b39f5;
    11'b00010110101: data <= 32'h3845baba;
    11'b00010110110: data <= 32'h4069bd58;
    11'b00010110111: data <= 32'h3f53baf5;
    11'b00010111000: data <= 32'h3602b86b;
    11'b00010111001: data <= 32'h2c30b6fc;
    11'b00010111010: data <= 32'h3bb53156;
    11'b00010111011: data <= 32'h3c133a80;
    11'b00010111100: data <= 32'hb8c53260;
    11'b00010111101: data <= 32'hc046bdf2;
    11'b00010111110: data <= 32'hbf8ac07b;
    11'b00010111111: data <= 32'hb825bc26;
    11'b00011000000: data <= 32'h33be382a;
    11'b00011000001: data <= 32'h306d3845;
    11'b00011000010: data <= 32'h2d76b526;
    11'b00011000011: data <= 32'h305c2c2d;
    11'b00011000100: data <= 32'hb7cd3f2f;
    11'b00011000101: data <= 32'hbde8413e;
    11'b00011000110: data <= 32'hbd6c3d19;
    11'b00011000111: data <= 32'h3193b958;
    11'b00011001000: data <= 32'h3d93bc77;
    11'b00011001001: data <= 32'h3c1fb3c0;
    11'b00011001010: data <= 32'h343835e6;
    11'b00011001011: data <= 32'h3ac234ce;
    11'b00011001100: data <= 32'h40483621;
    11'b00011001101: data <= 32'h3f983960;
    11'b00011001110: data <= 32'hb3de31f6;
    11'b00011001111: data <= 32'hbfd0bc75;
    11'b00011010000: data <= 32'hbdabbf31;
    11'b00011010001: data <= 32'h336dbc93;
    11'b00011010010: data <= 32'h3a99b6c2;
    11'b00011010011: data <= 32'h314cbac8;
    11'b00011010100: data <= 32'hb57abd9c;
    11'b00011010101: data <= 32'hb440b54e;
    11'b00011010110: data <= 32'hb8373f38;
    11'b00011010111: data <= 32'hbd6040fe;
    11'b00011011000: data <= 32'hbe683ad4;
    11'b00011011001: data <= 32'hba43bc05;
    11'b00011011010: data <= 32'h24a2bb61;
    11'b00011011011: data <= 32'haa943770;
    11'b00011011100: data <= 32'ha94f3c6e;
    11'b00011011101: data <= 32'h3c93392c;
    11'b00011011110: data <= 32'h40ed36c7;
    11'b00011011111: data <= 32'h3fa13b4b;
    11'b00011100000: data <= 32'hb4e73bfb;
    11'b00011100001: data <= 32'hbe682c4a;
    11'b00011100010: data <= 32'hb862bb32;
    11'b00011100011: data <= 32'h3cb8bc32;
    11'b00011100100: data <= 32'h3d5abc2f;
    11'b00011100101: data <= 32'h32d7be72;
    11'b00011100110: data <= 32'hb48bbf56;
    11'b00011100111: data <= 32'h33dab81b;
    11'b00011101000: data <= 32'h355a3da5;
    11'b00011101001: data <= 32'hb9d83ea0;
    11'b00011101010: data <= 32'hbf16aecb;
    11'b00011101011: data <= 32'hbecfbe1f;
    11'b00011101100: data <= 32'hbc59bac9;
    11'b00011101101: data <= 32'hba4c39c1;
    11'b00011101110: data <= 32'hb5b23c0d;
    11'b00011101111: data <= 32'h3ac0314b;
    11'b00011110000: data <= 32'h3f612dd3;
    11'b00011110001: data <= 32'h3c953d2c;
    11'b00011110010: data <= 32'hb988403b;
    11'b00011110011: data <= 32'hbd573d74;
    11'b00011110100: data <= 32'h2a99a914;
    11'b00011110101: data <= 32'h3e1cba25;
    11'b00011110110: data <= 32'h3cedbbd3;
    11'b00011110111: data <= 32'h2d42bd6c;
    11'b00011111000: data <= 32'h313fbdaf;
    11'b00011111001: data <= 32'h3d91b605;
    11'b00011111010: data <= 32'h3e9c3b8b;
    11'b00011111011: data <= 32'h2d303a46;
    11'b00011111100: data <= 32'hbebcba73;
    11'b00011111101: data <= 32'hbff0bedd;
    11'b00011111110: data <= 32'hbd0dba6b;
    11'b00011111111: data <= 32'hba20362c;
    11'b00100000000: data <= 32'hb7ba2a06;
    11'b00100000001: data <= 32'h332abbfd;
    11'b00100000010: data <= 32'h3ab4b86c;
    11'b00100000011: data <= 32'h345b3def;
    11'b00100000100: data <= 32'hbc0d419a;
    11'b00100000101: data <= 32'hbcfc3fe5;
    11'b00100000110: data <= 32'ha5683469;
    11'b00100000111: data <= 32'h3b5ab780;
    11'b00100001000: data <= 32'h35e9b53b;
    11'b00100001001: data <= 32'hb559b60d;
    11'b00100001010: data <= 32'h38e5b89b;
    11'b00100001011: data <= 32'h40dcaebb;
    11'b00100001100: data <= 32'h4141397e;
    11'b00100001101: data <= 32'h38fa381e;
    11'b00100001110: data <= 32'hbd7db919;
    11'b00100001111: data <= 32'hbdecbcea;
    11'b00100010000: data <= 32'hb7c6b8eb;
    11'b00100010001: data <= 32'haf0bb2f5;
    11'b00100010010: data <= 32'hb677bcbd;
    11'b00100010011: data <= 32'hb49cc060;
    11'b00100010100: data <= 32'h32cabcbc;
    11'b00100010101: data <= 32'h28213d44;
    11'b00100010110: data <= 32'hbae54140;
    11'b00100010111: data <= 32'hbce33e37;
    11'b00100011000: data <= 32'hb91dade3;
    11'b00100011001: data <= 32'hb4c0b4f8;
    11'b00100011010: data <= 32'hbaa23713;
    11'b00100011011: data <= 32'hbb47386b;
    11'b00100011100: data <= 32'h398aa871;
    11'b00100011101: data <= 32'h415fab3a;
    11'b00100011110: data <= 32'h4154397e;
    11'b00100011111: data <= 32'h38a23bf7;
    11'b00100100000: data <= 32'hbc1d35ff;
    11'b00100100001: data <= 32'hb87eb2d7;
    11'b00100100010: data <= 32'h38fab323;
    11'b00100100011: data <= 32'h38b0b8b0;
    11'b00100100100: data <= 32'hb531bf7d;
    11'b00100100101: data <= 32'hb6eec15b;
    11'b00100100110: data <= 32'h368abdbe;
    11'b00100100111: data <= 32'h39b63b2b;
    11'b00100101000: data <= 32'hb08d3ef5;
    11'b00100101001: data <= 32'hbc523769;
    11'b00100101010: data <= 32'hbd19ba41;
    11'b00100101011: data <= 32'hbd43b487;
    11'b00100101100: data <= 32'hbea03aef;
    11'b00100101101: data <= 32'hbd673a04;
    11'b00100101110: data <= 32'h3537b538;
    11'b00100101111: data <= 32'h400db798;
    11'b00100110000: data <= 32'h3f363a13;
    11'b00100110001: data <= 32'h2ae83f3d;
    11'b00100110010: data <= 32'hba843e4c;
    11'b00100110011: data <= 32'h31bb3a1c;
    11'b00100110100: data <= 32'h3cfa33a9;
    11'b00100110101: data <= 32'h396cb686;
    11'b00100110110: data <= 32'hb820be4a;
    11'b00100110111: data <= 32'hb47dc068;
    11'b00100111000: data <= 32'h3cf7bcc6;
    11'b00100111001: data <= 32'h3fb1379f;
    11'b00100111010: data <= 32'h3a6f39fe;
    11'b00100111011: data <= 32'hba1cb7e0;
    11'b00100111100: data <= 32'hbd9cbcb1;
    11'b00100111101: data <= 32'hbdcab28d;
    11'b00100111110: data <= 32'hbe743a74;
    11'b00100111111: data <= 32'hbdad2e7d;
    11'b00101000000: data <= 32'hb428bd7a;
    11'b00101000001: data <= 32'h3b5bbd0a;
    11'b00101000010: data <= 32'h3992397b;
    11'b00101000011: data <= 32'hb7a1409c;
    11'b00101000100: data <= 32'hb9c44046;
    11'b00101000101: data <= 32'h35b33c66;
    11'b00101000110: data <= 32'h3b9b3849;
    11'b00101000111: data <= 32'haa4d337f;
    11'b00101001000: data <= 32'hbc48b818;
    11'b00101001001: data <= 32'hafa6bc9a;
    11'b00101001010: data <= 32'h401db9bc;
    11'b00101001011: data <= 32'h41b233a4;
    11'b00101001100: data <= 32'h3da13414;
    11'b00101001101: data <= 32'hb655b915;
    11'b00101001110: data <= 32'hbb00bab7;
    11'b00101001111: data <= 32'hb8c92ef2;
    11'b00101010000: data <= 32'hba463802;
    11'b00101010001: data <= 32'hbc99bb15;
    11'b00101010010: data <= 32'hb9e4c103;
    11'b00101010011: data <= 32'h2dffbff4;
    11'b00101010100: data <= 32'h30b3367b;
    11'b00101010101: data <= 32'hb8014022;
    11'b00101010110: data <= 32'hb8bb3e9f;
    11'b00101010111: data <= 32'h28d938cc;
    11'b00101011000: data <= 32'h99ad3843;
    11'b00101011001: data <= 32'hbcc43bb4;
    11'b00101011010: data <= 32'hbf1838c3;
    11'b00101011011: data <= 32'hb278b4ed;
    11'b00101011100: data <= 32'h4070b78a;
    11'b00101011101: data <= 32'h41aa3135;
    11'b00101011110: data <= 32'h3d1a3715;
    11'b00101011111: data <= 32'hb1832e40;
    11'b00101100000: data <= 32'h213b2efe;
    11'b00101100001: data <= 32'h39533930;
    11'b00101100010: data <= 32'h326a356f;
    11'b00101100011: data <= 32'hbaddbdca;
    11'b00101100100: data <= 32'hbb6bc1ea;
    11'b00101100101: data <= 32'h2127c066;
    11'b00101100110: data <= 32'h38472b3e;
    11'b00101100111: data <= 32'h30483ccc;
    11'b00101101000: data <= 32'hb4b336d0;
    11'b00101101001: data <= 32'hb5b2b5c2;
    11'b00101101010: data <= 32'hbaf4357a;
    11'b00101101011: data <= 32'hbff63da0;
    11'b00101101100: data <= 32'hc0723c3b;
    11'b00101101101: data <= 32'hb866b4b2;
    11'b00101101110: data <= 32'h3e3aba3b;
    11'b00101101111: data <= 32'h3f662d6a;
    11'b00101110000: data <= 32'h380e3bed;
    11'b00101110001: data <= 32'hb17c3c79;
    11'b00101110010: data <= 32'h3a063c45;
    11'b00101110011: data <= 32'h3e243cae;
    11'b00101110100: data <= 32'h38db386f;
    11'b00101110101: data <= 32'hbb4abc80;
    11'b00101110110: data <= 32'hbb46c0c2;
    11'b00101110111: data <= 32'h3883beff;
    11'b00101111000: data <= 32'h3e29b156;
    11'b00101111001: data <= 32'h3c4032f2;
    11'b00101111010: data <= 32'h2febba1b;
    11'b00101111011: data <= 32'hb64cbc4a;
    11'b00101111100: data <= 32'hbba13416;
    11'b00101111101: data <= 32'hbf7b3dd6;
    11'b00101111110: data <= 32'hc0423987;
    11'b00101111111: data <= 32'hbbbdbc71;
    11'b00110000000: data <= 32'h3762be28;
    11'b00110000001: data <= 32'h382fafac;
    11'b00110000010: data <= 32'hb5903d63;
    11'b00110000011: data <= 32'hb4433e72;
    11'b00110000100: data <= 32'h3c143d68;
    11'b00110000101: data <= 32'h3e1b3d6d;
    11'b00110000110: data <= 32'h301a3c44;
    11'b00110000111: data <= 32'hbdb4aca4;
    11'b00110001000: data <= 32'hbb28bc80;
    11'b00110001001: data <= 32'h3ccfbba1;
    11'b00110001010: data <= 32'h40beb252;
    11'b00110001011: data <= 32'h3e8bb586;
    11'b00110001100: data <= 32'h3705bcc4;
    11'b00110001101: data <= 32'h2abebc0a;
    11'b00110001110: data <= 32'haece380e;
    11'b00110001111: data <= 32'hbae43d39;
    11'b00110010000: data <= 32'hbe3cadad;
    11'b00110010001: data <= 32'hbceac044;
    11'b00110010010: data <= 32'hb69ec083;
    11'b00110010011: data <= 32'hb4f8b669;
    11'b00110010100: data <= 32'hb9593c8f;
    11'b00110010101: data <= 32'hb33f3c7a;
    11'b00110010110: data <= 32'h3acd3997;
    11'b00110010111: data <= 32'h3a6d3c55;
    11'b00110011000: data <= 32'hbb083e57;
    11'b00110011001: data <= 32'hc0423c46;
    11'b00110011010: data <= 32'hbc1994ef;
    11'b00110011011: data <= 32'h3d64b634;
    11'b00110011100: data <= 32'h40abb0da;
    11'b00110011101: data <= 32'h3d87b4c0;
    11'b00110011110: data <= 32'h36f1b9ac;
    11'b00110011111: data <= 32'h39f9b316;
    11'b00110100000: data <= 32'h3cbc3c35;
    11'b00110100001: data <= 32'h36543ceb;
    11'b00110100010: data <= 32'hbb71b8ba;
    11'b00110100011: data <= 32'hbd10c11a;
    11'b00110100100: data <= 32'hb8f8c0c1;
    11'b00110100101: data <= 32'hb221b88f;
    11'b00110100110: data <= 32'hb32d36f5;
    11'b00110100111: data <= 32'h2c71b045;
    11'b00110101000: data <= 32'h3892b828;
    11'b00110101001: data <= 32'h289c3869;
    11'b00110101010: data <= 32'hbe8a3f67;
    11'b00110101011: data <= 32'hc10c3e8f;
    11'b00110101100: data <= 32'hbcfc34bf;
    11'b00110101101: data <= 32'h3a7eb788;
    11'b00110101110: data <= 32'h3d51b2b5;
    11'b00110101111: data <= 32'h35f72f84;
    11'b00110110000: data <= 32'h2e6b31a6;
    11'b00110110001: data <= 32'h3d303975;
    11'b00110110010: data <= 32'h404b3e32;
    11'b00110110011: data <= 32'h3c643d7e;
    11'b00110110100: data <= 32'hb9c9b5ba;
    11'b00110110101: data <= 32'hbccdbfcf;
    11'b00110110110: data <= 32'hb2afbed9;
    11'b00110110111: data <= 32'h392bb7a4;
    11'b00110111000: data <= 32'h390eb5a6;
    11'b00110111001: data <= 32'h37cbbda0;
    11'b00110111010: data <= 32'h381ebe25;
    11'b00110111011: data <= 32'hae6c3181;
    11'b00110111100: data <= 32'hbdfd3f4d;
    11'b00110111101: data <= 32'hc07f3da8;
    11'b00110111110: data <= 32'hbd83b529;
    11'b00110111111: data <= 32'hae18bc88;
    11'b00111000000: data <= 32'haccab6d5;
    11'b00111000001: data <= 32'hba553722;
    11'b00111000010: data <= 32'hb5073976;
    11'b00111000011: data <= 32'h3dd33b9f;
    11'b00111000100: data <= 32'h408d3e62;
    11'b00111000101: data <= 32'h3ac13e91;
    11'b00111000110: data <= 32'hbc6f3829;
    11'b00111000111: data <= 32'hbccbb905;
    11'b00111001000: data <= 32'h35dfb8dc;
    11'b00111001001: data <= 32'h3dd1b16e;
    11'b00111001010: data <= 32'h3cc4ba44;
    11'b00111001011: data <= 32'h39a4bfe2;
    11'b00111001100: data <= 32'h3a23bee9;
    11'b00111001101: data <= 32'h38bf3424;
    11'b00111001110: data <= 32'hb6dc3eb3;
    11'b00111001111: data <= 32'hbd8639c7;
    11'b00111010000: data <= 32'hbd2bbd26;
    11'b00111010001: data <= 32'hba8dbf55;
    11'b00111010010: data <= 32'hbc2bb932;
    11'b00111010011: data <= 32'hbd943616;
    11'b00111010100: data <= 32'hb7a73516;
    11'b00111010101: data <= 32'h3d173407;
    11'b00111010110: data <= 32'h3ea33c34;
    11'b00111010111: data <= 32'hac9e3f47;
    11'b00111011000: data <= 32'hbf253dfe;
    11'b00111011001: data <= 32'hbd343904;
    11'b00111011010: data <= 32'h38d43443;
    11'b00111011011: data <= 32'h3e102fcf;
    11'b00111011100: data <= 32'h3b39b996;
    11'b00111011101: data <= 32'h3767be70;
    11'b00111011110: data <= 32'h3c91bc41;
    11'b00111011111: data <= 32'h3ede3a17;
    11'b00111100000: data <= 32'h3ba23e5f;
    11'b00111100001: data <= 32'hb6cd3182;
    11'b00111100010: data <= 32'hbc2ebf1c;
    11'b00111100011: data <= 32'hbbb7bfba;
    11'b00111100100: data <= 32'hbc3bb8f8;
    11'b00111100101: data <= 32'hbc74a8d3;
    11'b00111100110: data <= 32'hb402ba2f;
    11'b00111100111: data <= 32'h3c01bc56;
    11'b00111101000: data <= 32'h3b0f31dd;
    11'b00111101001: data <= 32'hbb013f15;
    11'b00111101010: data <= 32'hc0573fed;
    11'b00111101011: data <= 32'hbd793c47;
    11'b00111101100: data <= 32'h350d363a;
    11'b00111101101: data <= 32'h394a3160;
    11'b00111101110: data <= 32'hb2d7b4b2;
    11'b00111101111: data <= 32'hb27cb9fc;
    11'b00111110000: data <= 32'h3d72b07d;
    11'b00111110001: data <= 32'h41263d0a;
    11'b00111110010: data <= 32'h3f3c3e7f;
    11'b00111110011: data <= 32'h27613254;
    11'b00111110100: data <= 32'hbaa8bd45;
    11'b00111110101: data <= 32'hb86ebcb2;
    11'b00111110110: data <= 32'hb465b2c8;
    11'b00111110111: data <= 32'hb453b7da;
    11'b00111111000: data <= 32'h3180bfb7;
    11'b00111111001: data <= 32'h3af9c086;
    11'b00111111010: data <= 32'h38a4b7ae;
    11'b00111111011: data <= 32'hbaed3e36;
    11'b00111111100: data <= 32'hbf4b3ef9;
    11'b00111111101: data <= 32'hbcd5383f;
    11'b00111111110: data <= 32'hb439b31e;
    11'b00111111111: data <= 32'hb8f4a9d3;
    11'b01000000000: data <= 32'hbe2d2cdd;
    11'b01000000001: data <= 32'hbb74af88;
    11'b01000000010: data <= 32'h3d2633e7;
    11'b01000000011: data <= 32'h41583d09;
    11'b01000000100: data <= 32'h3ea33e8c;
    11'b01000000101: data <= 32'hb4353a1e;
    11'b01000000110: data <= 32'hba72afb3;
    11'b01000000111: data <= 32'h29672e35;
    11'b01000001000: data <= 32'h38f236ee;
    11'b01000001001: data <= 32'h3640b93d;
    11'b01000001010: data <= 32'h35e2c0e5;
    11'b01000001011: data <= 32'h3b49c128;
    11'b01000001100: data <= 32'h3be6b843;
    11'b01000001101: data <= 32'h2ca13d63;
    11'b01000001110: data <= 32'hba623c29;
    11'b01000001111: data <= 32'hba31b7bb;
    11'b01000010000: data <= 32'hb990bc02;
    11'b01000010001: data <= 32'hbe1fb43e;
    11'b01000010010: data <= 32'hc09831c1;
    11'b01000010011: data <= 32'hbd22b33e;
    11'b01000010100: data <= 32'h3c0cb525;
    11'b01000010101: data <= 32'h40183896;
    11'b01000010110: data <= 32'h39ce3de0;
    11'b01000010111: data <= 32'hbbf63dbc;
    11'b01000011000: data <= 32'hbb543c45;
    11'b01000011001: data <= 32'h36893c94;
    11'b01000011010: data <= 32'h3b3a3bb1;
    11'b01000011011: data <= 32'h3385b702;
    11'b01000011100: data <= 32'h20f8c027;
    11'b01000011101: data <= 32'h3ba8bfb9;
    11'b01000011110: data <= 32'h3f309f47;
    11'b01000011111: data <= 32'h3d853d19;
    11'b01000100000: data <= 32'h35953649;
    11'b01000100001: data <= 32'hb3d7bca8;
    11'b01000100010: data <= 32'hb959bcf0;
    11'b01000100011: data <= 32'hbe22b0d0;
    11'b01000100100: data <= 32'hc0232bcf;
    11'b01000100101: data <= 32'hbc4abc09;
    11'b01000100110: data <= 32'h39eebe4c;
    11'b01000100111: data <= 32'h3ccbb7e0;
    11'b01000101000: data <= 32'hb3a93c69;
    11'b01000101001: data <= 32'hbe0b3ed4;
    11'b01000101010: data <= 32'hbb673dfb;
    11'b01000101011: data <= 32'h362c3d6e;
    11'b01000101100: data <= 32'h35843c4b;
    11'b01000101101: data <= 32'hba51a371;
    11'b01000101110: data <= 32'hbacebca7;
    11'b01000101111: data <= 32'h3ab5bb03;
    11'b01000110000: data <= 32'h40d338ed;
    11'b01000110001: data <= 32'h406d3d19;
    11'b01000110010: data <= 32'h3b72320a;
    11'b01000110011: data <= 32'h2db8bbe3;
    11'b01000110100: data <= 32'hb2b9b89e;
    11'b01000110101: data <= 32'hb9b63714;
    11'b01000110110: data <= 32'hbc83aa03;
    11'b01000110111: data <= 32'hb850bf9c;
    11'b01000111000: data <= 32'h38d2c174;
    11'b01000111001: data <= 32'h399cbd44;
    11'b01000111010: data <= 32'hb7e939aa;
    11'b01000111011: data <= 32'hbd1b3d8a;
    11'b01000111100: data <= 32'hb8d13b71;
    11'b01000111101: data <= 32'h30b33983;
    11'b01000111110: data <= 32'hb94d3a31;
    11'b01000111111: data <= 32'hc02f359f;
    11'b01001000000: data <= 32'hbf13b5f0;
    11'b01001000001: data <= 32'h384eb3bb;
    11'b01001000010: data <= 32'h40c839f2;
    11'b01001000011: data <= 32'h40173c9b;
    11'b01001000100: data <= 32'h38ff36db;
    11'b01001000101: data <= 32'h2c51ac5b;
    11'b01001000110: data <= 32'h361d3949;
    11'b01001000111: data <= 32'h34fa3d2f;
    11'b01001001000: data <= 32'hb3b22b5f;
    11'b01001001001: data <= 32'hb27dc08a;
    11'b01001001010: data <= 32'h3850c211;
    11'b01001001011: data <= 32'h3a6cbd9a;
    11'b01001001100: data <= 32'h31213808;
    11'b01001001101: data <= 32'hb4b03965;
    11'b01001001110: data <= 32'h2a90b223;
    11'b01001001111: data <= 32'h242cb4ac;
    11'b01001010000: data <= 32'hbd943689;
    11'b01001010001: data <= 32'hc1b03832;
    11'b01001010010: data <= 32'hc065b272;
    11'b01001010011: data <= 32'h32cfb834;
    11'b01001010100: data <= 32'h3ef42f79;
    11'b01001010101: data <= 32'h3c193a23;
    11'b01001010110: data <= 32'hb4743a34;
    11'b01001010111: data <= 32'hb1e23b5b;
    11'b01001011000: data <= 32'h3a553ede;
    11'b01001011001: data <= 32'h3ac43fcc;
    11'b01001011010: data <= 32'haf4b360c;
    11'b01001011011: data <= 32'hb7acbf65;
    11'b01001011100: data <= 32'h3629c0a1;
    11'b01001011101: data <= 32'h3d1eb9ea;
    11'b01001011110: data <= 32'h3cfd3874;
    11'b01001011111: data <= 32'h3aef065c;
    11'b01001100000: data <= 32'h39fabc62;
    11'b01001100001: data <= 32'h3267ba68;
    11'b01001100010: data <= 32'hbd4c36b6;
    11'b01001100011: data <= 32'hc12238a6;
    11'b01001100100: data <= 32'hbf94b93b;
    11'b01001100101: data <= 32'h293bbe2b;
    11'b01001100110: data <= 32'h3af6bbae;
    11'b01001100111: data <= 32'hb07e3275;
    11'b01001101000: data <= 32'hbc403abd;
    11'b01001101001: data <= 32'hb5103cfe;
    11'b01001101010: data <= 32'h3b523f9f;
    11'b01001101011: data <= 32'h38db4009;
    11'b01001101100: data <= 32'hbb1e39e9;
    11'b01001101101: data <= 32'hbd5ebb54;
    11'b01001101110: data <= 32'h2a0ebc56;
    11'b01001101111: data <= 32'h3e983086;
    11'b01001110000: data <= 32'h3fd83991;
    11'b01001110001: data <= 32'h3dcab528;
    11'b01001110010: data <= 32'h3c62bce5;
    11'b01001110011: data <= 32'h3923b676;
    11'b01001110100: data <= 32'hb7ae3bfb;
    11'b01001110101: data <= 32'hbde53995;
    11'b01001110110: data <= 32'hbc7dbd16;
    11'b01001110111: data <= 32'h2a65c11a;
    11'b01001111000: data <= 32'h347cbf35;
    11'b01001111001: data <= 32'hb982b435;
    11'b01001111010: data <= 32'hbc6637bd;
    11'b01001111011: data <= 32'ha792392f;
    11'b01001111100: data <= 32'h3b2a3c73;
    11'b01001111101: data <= 32'haece3e0c;
    11'b01001111110: data <= 32'hc0103bac;
    11'b01001111111: data <= 32'hc095aaa9;
    11'b01010000000: data <= 32'hb5f6b170;
    11'b01010000001: data <= 32'h3e28386c;
    11'b01010000010: data <= 32'h3ef83915;
    11'b01010000011: data <= 32'h3c30b49e;
    11'b01010000100: data <= 32'h3b45b8e3;
    11'b01010000101: data <= 32'h3c6b3943;
    11'b01010000110: data <= 32'h38d03f91;
    11'b01010000111: data <= 32'hb5303bb4;
    11'b01010001000: data <= 32'hb7e6be03;
    11'b01010001001: data <= 32'h2cfac196;
    11'b01010001010: data <= 32'h323ebf4b;
    11'b01010001011: data <= 32'hb588b5a7;
    11'b01010001100: data <= 32'hb4ffb007;
    11'b01010001101: data <= 32'h394fb82f;
    11'b01010001110: data <= 32'h3ba7af17;
    11'b01010001111: data <= 32'hb94f3ad3;
    11'b01010010000: data <= 32'hc16a3c10;
    11'b01010010001: data <= 32'hc1623480;
    11'b01010010010: data <= 32'hb91eb06d;
    11'b01010010011: data <= 32'h3b99309f;
    11'b01010010100: data <= 32'h3963331b;
    11'b01010010101: data <= 32'hacb7b0e9;
    11'b01010010110: data <= 32'h35ff315f;
    11'b01010010111: data <= 32'h3d853e82;
    11'b01010011000: data <= 32'h3d1b4118;
    11'b01010011001: data <= 32'h2f923d20;
    11'b01010011010: data <= 32'hb835bc6b;
    11'b01010011011: data <= 32'had5ac00e;
    11'b01010011100: data <= 32'h373dbbc7;
    11'b01010011101: data <= 32'h3808a921;
    11'b01010011110: data <= 32'h39fdb94b;
    11'b01010011111: data <= 32'h3d90be31;
    11'b01010100000: data <= 32'h3cc7bb76;
    11'b01010100001: data <= 32'hb89538c5;
    11'b01010100010: data <= 32'hc0c33c33;
    11'b01010100011: data <= 32'hc07629d2;
    11'b01010100100: data <= 32'hb8abbb25;
    11'b01010100101: data <= 32'h32cfba86;
    11'b01010100110: data <= 32'hb8cbb651;
    11'b01010100111: data <= 32'hbca9b21c;
    11'b01010101000: data <= 32'ha9bf36f7;
    11'b01010101001: data <= 32'h3dd03f13;
    11'b01010101010: data <= 32'h3cfa4100;
    11'b01010101011: data <= 32'hb6093dd4;
    11'b01010101100: data <= 32'hbcfeb49a;
    11'b01010101101: data <= 32'hb7aeb996;
    11'b01010101110: data <= 32'h396832a1;
    11'b01010101111: data <= 32'h3c763661;
    11'b01010110000: data <= 32'h3d21bb41;
    11'b01010110001: data <= 32'h3eaabf7b;
    11'b01010110010: data <= 32'h3e03baa5;
    11'b01010110011: data <= 32'h31b63c08;
    11'b01010110100: data <= 32'hbccd3ce1;
    11'b01010110101: data <= 32'hbcb3b660;
    11'b01010110110: data <= 32'hb454bf10;
    11'b01010110111: data <= 32'hb47abe70;
    11'b01010111000: data <= 32'hbd52baa3;
    11'b01010111001: data <= 32'hbe0db797;
    11'b01010111010: data <= 32'h29dcae83;
    11'b01010111011: data <= 32'h3de33b2f;
    11'b01010111100: data <= 32'h39c53ef0;
    11'b01010111101: data <= 32'hbd683d86;
    11'b01010111110: data <= 32'hc0493773;
    11'b01010111111: data <= 32'hbb423637;
    11'b01011000000: data <= 32'h38ab3b8c;
    11'b01011000001: data <= 32'h3b6b3888;
    11'b01011000010: data <= 32'h3a8abb22;
    11'b01011000011: data <= 32'h3d07bdd4;
    11'b01011000100: data <= 32'h3ec4288c;
    11'b01011000101: data <= 32'h3c943f58;
    11'b01011000110: data <= 32'h2f253e15;
    11'b01011000111: data <= 32'hb2b5b8c5;
    11'b01011001000: data <= 32'h245fc002;
    11'b01011001001: data <= 32'hb5bebe4f;
    11'b01011001010: data <= 32'hbcc6b9ef;
    11'b01011001011: data <= 32'hbb97bac5;
    11'b01011001100: data <= 32'h3940bca6;
    11'b01011001101: data <= 32'h3e58b79b;
    11'b01011001110: data <= 32'h33b039e4;
    11'b01011001111: data <= 32'hbff93c9b;
    11'b01011010000: data <= 32'hc1003a22;
    11'b01011010001: data <= 32'hbc2b390a;
    11'b01011010010: data <= 32'h31fa3a50;
    11'b01011010011: data <= 32'ha9b7342d;
    11'b01011010100: data <= 32'hb711ba89;
    11'b01011010101: data <= 32'h3649ba53;
    11'b01011010110: data <= 32'h3eaa3b8b;
    11'b01011010111: data <= 32'h3f0e40eb;
    11'b01011011000: data <= 32'h3a1d3f04;
    11'b01011011001: data <= 32'h2974b574;
    11'b01011011010: data <= 32'h9897bd45;
    11'b01011011011: data <= 32'hb117b8d1;
    11'b01011011100: data <= 32'hb7c4af75;
    11'b01011011101: data <= 32'h258cbc50;
    11'b01011011110: data <= 32'h3d6fc03b;
    11'b01011011111: data <= 32'h3f22be05;
    11'b01011100000: data <= 32'h33973154;
    11'b01011100001: data <= 32'hbee93c05;
    11'b01011100010: data <= 32'hbfbc389a;
    11'b01011100011: data <= 32'hb9a02919;
    11'b01011100100: data <= 32'hb423aa37;
    11'b01011100101: data <= 32'hbcf4b548;
    11'b01011100110: data <= 32'hbef5bad3;
    11'b01011100111: data <= 32'hb5ceb7a3;
    11'b01011101000: data <= 32'h3e143c81;
    11'b01011101001: data <= 32'h3f0740a8;
    11'b01011101010: data <= 32'h373a3ebd;
    11'b01011101011: data <= 32'hb82c329e;
    11'b01011101100: data <= 32'hb5c5ac45;
    11'b01011101101: data <= 32'h28b03a3c;
    11'b01011101110: data <= 32'h300e3963;
    11'b01011101111: data <= 32'h38a2bc4c;
    11'b01011110000: data <= 32'h3e4ec0e3;
    11'b01011110001: data <= 32'h3f93be68;
    11'b01011110010: data <= 32'h3a01361d;
    11'b01011110011: data <= 32'hb8fc3c74;
    11'b01011110100: data <= 32'hb979319e;
    11'b01011110101: data <= 32'ha833ba57;
    11'b01011110110: data <= 32'hb7aabac1;
    11'b01011110111: data <= 32'hbfd6b9d8;
    11'b01011111000: data <= 32'hc099bbe9;
    11'b01011111001: data <= 32'hb80eba82;
    11'b01011111010: data <= 32'h3dc93545;
    11'b01011111011: data <= 32'h3d223d8a;
    11'b01011111100: data <= 32'hb72c3d07;
    11'b01011111101: data <= 32'hbd933965;
    11'b01011111110: data <= 32'hba283bfc;
    11'b01011111111: data <= 32'h29773ef7;
    11'b01100000000: data <= 32'h2e363c75;
    11'b01100000001: data <= 32'h31dcbb74;
    11'b01100000010: data <= 32'h3c0dc028;
    11'b01100000011: data <= 32'h3f00bab6;
    11'b01100000100: data <= 32'h3db73ca2;
    11'b01100000101: data <= 32'h39443d9c;
    11'b01100000110: data <= 32'h3826ad04;
    11'b01100000111: data <= 32'h3887bc97;
    11'b01100001000: data <= 32'hb64ebaff;
    11'b01100001001: data <= 32'hbf76b825;
    11'b01100001010: data <= 32'hbf78bc3f;
    11'b01100001011: data <= 32'h24c8be62;
    11'b01100001100: data <= 32'h3e2fbc06;
    11'b01100001101: data <= 32'h3a3c309b;
    11'b01100001110: data <= 32'hbcab3979;
    11'b01100001111: data <= 32'hbf393a36;
    11'b01100010000: data <= 32'hba7e3d19;
    11'b01100010001: data <= 32'hae403f01;
    11'b01100010010: data <= 32'hb8ef3b79;
    11'b01100010011: data <= 32'hbc21baa4;
    11'b01100010100: data <= 32'hadccbda6;
    11'b01100010101: data <= 32'h3d732f0a;
    11'b01100010110: data <= 32'h3f463f50;
    11'b01100010111: data <= 32'h3d5b3e4a;
    11'b01100011000: data <= 32'h3bb9a856;
    11'b01100011001: data <= 32'h39beb98a;
    11'b01100011010: data <= 32'hb0a62ac0;
    11'b01100011011: data <= 32'hbcb43553;
    11'b01100011100: data <= 32'hbb1ebb6e;
    11'b01100011101: data <= 32'h3a0ac099;
    11'b01100011110: data <= 32'h3ed3c01d;
    11'b01100011111: data <= 32'h38e0b931;
    11'b01100100000: data <= 32'hbc6b3514;
    11'b01100100001: data <= 32'hbd29380a;
    11'b01100100010: data <= 32'hb44939bc;
    11'b01100100011: data <= 32'hb1ff3b8b;
    11'b01100100100: data <= 32'hbe343545;
    11'b01100100101: data <= 32'hc0b0baca;
    11'b01100100110: data <= 32'hbc5dbbcc;
    11'b01100100111: data <= 32'h3b973783;
    11'b01100101000: data <= 32'h3ec83f06;
    11'b01100101001: data <= 32'h3c423d4e;
    11'b01100101010: data <= 32'h378631b8;
    11'b01100101011: data <= 32'h360734cb;
    11'b01100101100: data <= 32'h2b943dc7;
    11'b01100101101: data <= 32'hb7a33d89;
    11'b01100101110: data <= 32'hb1dfb8f2;
    11'b01100101111: data <= 32'h3c28c0f4;
    11'b01100110000: data <= 32'h3eb2c063;
    11'b01100110001: data <= 32'h3a89b857;
    11'b01100110010: data <= 32'hb40e35e3;
    11'b01100110011: data <= 32'ha8972de9;
    11'b01100110100: data <= 32'h3960b174;
    11'b01100110101: data <= 32'hacaa2774;
    11'b01100110110: data <= 32'hc031b096;
    11'b01100110111: data <= 32'hc1e6bb08;
    11'b01100111000: data <= 32'hbd8bbc2a;
    11'b01100111001: data <= 32'h3a29ad59;
    11'b01100111010: data <= 32'h3cc63a8a;
    11'b01100111011: data <= 32'h3052390e;
    11'b01100111100: data <= 32'hb7c534b4;
    11'b01100111101: data <= 32'hae823cac;
    11'b01100111110: data <= 32'h305c40ea;
    11'b01100111111: data <= 32'hb46e4008;
    11'b01101000000: data <= 32'hb592b51f;
    11'b01101000001: data <= 32'h37f3c01f;
    11'b01101000010: data <= 32'h3d1dbdb0;
    11'b01101000011: data <= 32'h3c8c3482;
    11'b01101000100: data <= 32'h3a8839b4;
    11'b01101000101: data <= 32'h3ce5b2a0;
    11'b01101000110: data <= 32'h3dfeb9bb;
    11'b01101000111: data <= 32'h32eeb2f3;
    11'b01101001000: data <= 32'hbfb527bd;
    11'b01101001001: data <= 32'hc10cb9d1;
    11'b01101001010: data <= 32'hbad0bde3;
    11'b01101001011: data <= 32'h3b39bcc9;
    11'b01101001100: data <= 32'h3946b7b3;
    11'b01101001101: data <= 32'hb9ebb268;
    11'b01101001110: data <= 32'hbc6230a0;
    11'b01101001111: data <= 32'hb2673d62;
    11'b01101010000: data <= 32'h31f540fc;
    11'b01101010001: data <= 32'hb9433f7c;
    11'b01101010010: data <= 32'hbd58b30f;
    11'b01101010011: data <= 32'hb945bd7b;
    11'b01101010100: data <= 32'h38e3b58a;
    11'b01101010101: data <= 32'h3cf13c85;
    11'b01101010110: data <= 32'h3d7f3ba0;
    11'b01101010111: data <= 32'h3eddb512;
    11'b01101011000: data <= 32'h3ef3b88b;
    11'b01101011001: data <= 32'h380937b2;
    11'b01101011010: data <= 32'hbcd73b5d;
    11'b01101011011: data <= 32'hbdcbb4f0;
    11'b01101011100: data <= 32'h2938bf6d;
    11'b01101011101: data <= 32'h3c91c035;
    11'b01101011110: data <= 32'h35e1bd5a;
    11'b01101011111: data <= 32'hbba9b9a8;
    11'b01101100000: data <= 32'hba7ab2de;
    11'b01101100001: data <= 32'h35da3a02;
    11'b01101100010: data <= 32'h35fe3e76;
    11'b01101100011: data <= 32'hbd093c8f;
    11'b01101100100: data <= 32'hc0fab517;
    11'b01101100101: data <= 32'hbef3bab7;
    11'b01101100110: data <= 32'h1fdc3444;
    11'b01101100111: data <= 32'h3bc93d25;
    11'b01101101000: data <= 32'h3c3339a8;
    11'b01101101001: data <= 32'h3cbab5d7;
    11'b01101101010: data <= 32'h3d3d2d99;
    11'b01101101011: data <= 32'h391f3ece;
    11'b01101101100: data <= 32'hb70c401e;
    11'b01101101101: data <= 32'hb8203371;
    11'b01101101110: data <= 32'h386ebf62;
    11'b01101101111: data <= 32'h3c89c05a;
    11'b01101110000: data <= 32'h356cbce4;
    11'b01101110001: data <= 32'hb705b8f3;
    11'b01101110010: data <= 32'h3438b8a8;
    11'b01101110011: data <= 32'h3d94b220;
    11'b01101110100: data <= 32'h39ff3805;
    11'b01101110101: data <= 32'hbe4c3718;
    11'b01101110110: data <= 32'hc206b660;
    11'b01101110111: data <= 32'hc01bb998;
    11'b01101111000: data <= 32'hb1ff28e8;
    11'b01101111001: data <= 32'h37b23852;
    11'b01101111010: data <= 32'h2c9aac95;
    11'b01101111011: data <= 32'h2b25b83c;
    11'b01101111100: data <= 32'h38f7398f;
    11'b01101111101: data <= 32'h392e413e;
    11'b01101111110: data <= 32'hac2e417b;
    11'b01101111111: data <= 32'hb5e038d3;
    11'b01110000000: data <= 32'h32f8bd97;
    11'b01110000001: data <= 32'h395cbd6a;
    11'b01110000010: data <= 32'h35f3b428;
    11'b01110000011: data <= 32'h358bad8d;
    11'b01110000100: data <= 32'h3daeba6b;
    11'b01110000101: data <= 32'h4099bb10;
    11'b01110000110: data <= 32'h3caaa967;
    11'b01110000111: data <= 32'hbd513653;
    11'b01110001000: data <= 32'hc112b281;
    11'b01110001001: data <= 32'hbda7bac9;
    11'b01110001010: data <= 32'h2e59ba30;
    11'b01110001011: data <= 32'h25b7b928;
    11'b01110001100: data <= 32'hbb66bc04;
    11'b01110001101: data <= 32'hbaafbada;
    11'b01110001110: data <= 32'h349d3a08;
    11'b01110001111: data <= 32'h39b04135;
    11'b01110010000: data <= 32'hb1cb410e;
    11'b01110010001: data <= 32'hbc2b38bb;
    11'b01110010010: data <= 32'hba79ba26;
    11'b01110010011: data <= 32'haf19b18a;
    11'b01110010100: data <= 32'h34003acd;
    11'b01110010101: data <= 32'h39f8364b;
    11'b01110010110: data <= 32'h3f70bb2e;
    11'b01110010111: data <= 32'h4106bbd1;
    11'b01110011000: data <= 32'h3d93356c;
    11'b01110011001: data <= 32'hb9363c8d;
    11'b01110011010: data <= 32'hbd773543;
    11'b01110011011: data <= 32'hb479bbda;
    11'b01110011100: data <= 32'h389dbdf2;
    11'b01110011101: data <= 32'hb367bdca;
    11'b01110011110: data <= 32'hbd73be1e;
    11'b01110011111: data <= 32'hbaefbcda;
    11'b01110100000: data <= 32'h397d316a;
    11'b01110100001: data <= 32'h3c013e93;
    11'b01110100010: data <= 32'hb81c3e54;
    11'b01110100011: data <= 32'hbfe2343a;
    11'b01110100100: data <= 32'hbf52b4a8;
    11'b01110100101: data <= 32'hba2d391e;
    11'b01110100110: data <= 32'hac6e3d4d;
    11'b01110100111: data <= 32'h365b3564;
    11'b01110101000: data <= 32'h3d04bc1c;
    11'b01110101001: data <= 32'h3f9fb8c3;
    11'b01110101010: data <= 32'h3d493d40;
    11'b01110101011: data <= 32'h2b33406b;
    11'b01110101100: data <= 32'hb4063bae;
    11'b01110101101: data <= 32'h3869bade;
    11'b01110101110: data <= 32'h3a41bdfc;
    11'b01110101111: data <= 32'hb515bd16;
    11'b01110110000: data <= 32'hbc76bd3a;
    11'b01110110001: data <= 32'hab7bbda1;
    11'b01110110010: data <= 32'h3e8eb9b4;
    11'b01110110011: data <= 32'h3df335dd;
    11'b01110110100: data <= 32'hb95b3893;
    11'b01110110101: data <= 32'hc0ccaa5b;
    11'b01110110110: data <= 32'hc030afb4;
    11'b01110110111: data <= 32'hbb0d3969;
    11'b01110111000: data <= 32'hb6f83ae3;
    11'b01110111001: data <= 32'hb843b594;
    11'b01110111010: data <= 32'ha4a4bd41;
    11'b01110111011: data <= 32'h3b54b1e4;
    11'b01110111100: data <= 32'h3c534036;
    11'b01110111101: data <= 32'h36f841b4;
    11'b01110111110: data <= 32'h30e53d2d;
    11'b01110111111: data <= 32'h3820b7b5;
    11'b01111000000: data <= 32'h36f4b99e;
    11'b01111000001: data <= 32'hb684b1bc;
    11'b01111000010: data <= 32'hb86db7f3;
    11'b01111000011: data <= 32'h3b92bd83;
    11'b01111000100: data <= 32'h4106bd8c;
    11'b01111000101: data <= 32'h3fa8b6c2;
    11'b01111000110: data <= 32'hb70d3296;
    11'b01111000111: data <= 32'hbfb49455;
    11'b01111001000: data <= 32'hbd5fb107;
    11'b01111001001: data <= 32'hb5982eef;
    11'b01111001010: data <= 32'hb944b0af;
    11'b01111001011: data <= 32'hbdffbd04;
    11'b01111001100: data <= 32'hbc90bec7;
    11'b01111001101: data <= 32'h340bb122;
    11'b01111001110: data <= 32'h3bb94023;
    11'b01111001111: data <= 32'h36994117;
    11'b01111010000: data <= 32'hb4403c4f;
    11'b01111010001: data <= 32'hb4e8ac0d;
    11'b01111010010: data <= 32'hb50d371f;
    11'b01111010011: data <= 32'hb8f03c99;
    11'b01111010100: data <= 32'hb39d3523;
    11'b01111010101: data <= 32'h3d61bd10;
    11'b01111010110: data <= 32'h414fbe33;
    11'b01111010111: data <= 32'h3ff0b4de;
    11'b01111011000: data <= 32'h2bc639ba;
    11'b01111011001: data <= 32'hba4a37c4;
    11'b01111011010: data <= 32'h9a0fb1bb;
    11'b01111011011: data <= 32'h376fb7a2;
    11'b01111011100: data <= 32'hb978bb18;
    11'b01111011101: data <= 32'hbfefbef0;
    11'b01111011110: data <= 32'hbdc1bfc9;
    11'b01111011111: data <= 32'h363ab8e3;
    11'b01111100000: data <= 32'h3cbe3c87;
    11'b01111100001: data <= 32'h32683da4;
    11'b01111100010: data <= 32'hbc1f36c4;
    11'b01111100011: data <= 32'hbcf7319c;
    11'b01111100100: data <= 32'hbba03d26;
    11'b01111100101: data <= 32'hbb193f92;
    11'b01111100110: data <= 32'hb800386e;
    11'b01111100111: data <= 32'h3a08bd2f;
    11'b01111101000: data <= 32'h3f86bd25;
    11'b01111101001: data <= 32'h3e6d37a7;
    11'b01111101010: data <= 32'h383b3eb5;
    11'b01111101011: data <= 32'h35883c6c;
    11'b01111101100: data <= 32'h3c64aafe;
    11'b01111101101: data <= 32'h3be2b832;
    11'b01111101110: data <= 32'hb91bb9bb;
    11'b01111101111: data <= 32'hbf62bd7f;
    11'b01111110000: data <= 32'hbabebf7b;
    11'b01111110001: data <= 32'h3cd0bd0f;
    11'b01111110010: data <= 32'h3ea8b0e9;
    11'b01111110011: data <= 32'h2d8b3034;
    11'b01111110100: data <= 32'hbdcbb357;
    11'b01111110101: data <= 32'hbe0031d9;
    11'b01111110110: data <= 32'hbbaa3db0;
    11'b01111110111: data <= 32'hbc1e3ea6;
    11'b01111111000: data <= 32'hbce52897;
    11'b01111111001: data <= 32'hb82bbe46;
    11'b01111111010: data <= 32'h3908bb93;
    11'b01111111011: data <= 32'h3c0d3ce3;
    11'b01111111100: data <= 32'h39bb4099;
    11'b01111111101: data <= 32'h3ab13d78;
    11'b01111111110: data <= 32'h3d4330d2;
    11'b01111111111: data <= 32'h3ab92e24;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    