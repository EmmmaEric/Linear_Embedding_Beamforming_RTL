
    module interp_rom_2(
    CLK, rst,
    Addr, CEB, Q
    );

    input CLK, rst;
    input [9:0] Addr;
    input CEB;		
    output [20:0] Q;

    (*rom_style = "block" *) reg [20:0] data;

    always @(posedge CLK) begin
    if (rst) begin
        data <= 20'd0;
    end else begin
    if (CEB)
    case(Addr)
            10'b00000000: data <= 20'b00101001110010001010;
        10'b00000001: data <= 20'b10101101010010110111;
        10'b00000010: data <= 20'b00011100011010110000;
        10'b00000011: data <= 20'b00101101011010001011;
        10'b00000100: data <= 20'b00100110100001110110;
        10'b00000101: data <= 20'b10101000110011000101;
        10'b00000110: data <= 20'b00101000100010001110;
        10'b00000111: data <= 20'b10101001010010100000;
        10'b00001000: data <= 20'b00110011110011011010;
        10'b00001001: data <= 20'b00101000010001110100;
        10'b00001010: data <= 20'b00100011010010100011;
        10'b00001011: data <= 20'b10110011000011000000;
        10'b00001100: data <= 20'b00101110100010110010;
        10'b00001101: data <= 20'b10100000011010011000;
        10'b00001110: data <= 20'b10101101111010011001;
        10'b00001111: data <= 20'b00100100101010000101;
        10'b00010000: data <= 20'b10101001010010110111;
        10'b00010001: data <= 20'b10100101011010110000;
        10'b00010010: data <= 20'b10101101000010100100;
        10'b00010011: data <= 20'b10100111110010100001;
        10'b00010100: data <= 20'b10100100111010100110;
        10'b00010101: data <= 20'b00100101110010100010;
        10'b00010110: data <= 20'b10101000000010010101;
        10'b00010111: data <= 20'b00101111001010000100;
        10'b00011000: data <= 20'b10100010001010101100;
        10'b00011001: data <= 20'b00110110000011001100;
        10'b00011010: data <= 20'b00110000100011010001;
        10'b00011011: data <= 20'b10101000001010110111;
        10'b00011100: data <= 20'b00101100001010100010;
        10'b00011101: data <= 20'b00101000111010011001;
        10'b00011110: data <= 20'b00101101010001110110;
        10'b00011111: data <= 20'b00101100101001111101;
        10'b00100000: data <= 20'b10100011100010011101;
        10'b00100001: data <= 20'b10100111110010010010;
        10'b00100010: data <= 20'b10101100110010110001;
        10'b00100011: data <= 20'b10100100110010100110;
        10'b00100100: data <= 20'b00101011000010010000;
        10'b00100101: data <= 20'b10011101010010100001;
        10'b00100110: data <= 20'b10101001101010100001;
        10'b00100111: data <= 20'b10101011100011000001;
        10'b00101000: data <= 20'b00100100100010000100;
        10'b00101001: data <= 20'b10101111101010111110;
        10'b00101010: data <= 20'b00101000100010000011;
        10'b00101011: data <= 20'b00110000010011000010;
        10'b00101100: data <= 20'b00101111001010010000;
        10'b00101101: data <= 20'b00101010011010101011;
        10'b00101110: data <= 20'b10101010101010000110;
        10'b00101111: data <= 20'b10011110110010100000;
        10'b00110000: data <= 20'b00101111010010100110;
        10'b00110001: data <= 20'b10100111101010000101;
        10'b00110010: data <= 20'b10101100111011001010;
        10'b00110011: data <= 20'b10011111110001111011;
        10'b00110100: data <= 20'b00100101100011000111;
        10'b00110101: data <= 20'b00011110011010110001;
        10'b00110110: data <= 20'b00101100100010100100;
        10'b00110111: data <= 20'b10100001001010011111;
        10'b00111000: data <= 20'b10100100110010110000;
        10'b00111001: data <= 20'b00011110010010000111;
        10'b00111010: data <= 20'b10101000110010110000;
        10'b00111011: data <= 20'b00101010000010101010;
        10'b00111100: data <= 20'b00101100000010100110;
        10'b00111101: data <= 20'b10101011101010101001;
        10'b00111110: data <= 20'b00101001010010011001;
        10'b00111111: data <= 20'b00101001100010000101;
        10'b01000000: data <= 20'b00101000100010011011;
        10'b01000001: data <= 20'b10101101110010111101;
        10'b01000010: data <= 20'b10100001000010010101;
        10'b01000011: data <= 20'b10100000010010110010;
        10'b01000100: data <= 20'b10101100110010100111;
        10'b01000101: data <= 20'b00100111100001110000;
        10'b01000110: data <= 20'b10101101101010101011;
        10'b01000111: data <= 20'b00100111101010010011;
        10'b01001000: data <= 20'b00111000001011011100;
        10'b01001001: data <= 20'b10110010110011000000;
        10'b01001010: data <= 20'b10101010001001111100;
        10'b01001011: data <= 20'b10110010101010101000;
        10'b01001100: data <= 20'b10110000001011000000;
        10'b01001101: data <= 20'b10110000100010010111;
        10'b01001110: data <= 20'b10100010001010001101;
        10'b01001111: data <= 20'b10101111010010101101;
        10'b01010000: data <= 20'b00101001000010101010;
        10'b01010001: data <= 20'b10100110000010110001;
        10'b01010010: data <= 20'b10101100110001100010;
        10'b01010011: data <= 20'b10110000111001111111;
        10'b01010100: data <= 20'b00100001111001010110;
        10'b01010101: data <= 20'b00101011010010110001;
        10'b01010110: data <= 20'b10101111101010101111;
        10'b01010111: data <= 20'b00101111101010100001;
        10'b01011000: data <= 20'b00101000000010000001;
        10'b01011001: data <= 20'b00100100100010100001;
        10'b01011010: data <= 20'b10100111001001101101;
        10'b01011011: data <= 20'b00101000100010011110;
        10'b01011100: data <= 20'b10101000100011001010;
        10'b01011101: data <= 20'b10101101110010111000;
        10'b01011110: data <= 20'b10101100101010100000;
        10'b01011111: data <= 20'b00011111101010111001;
        10'b01100000: data <= 20'b10100110101010101011;
        10'b01100001: data <= 20'b10101010100010101101;
        10'b01100010: data <= 20'b00101000101010010011;
        10'b01100011: data <= 20'b10100011011011000101;
        10'b01100100: data <= 20'b00101101000000110000;
        10'b01100101: data <= 20'b00100000100010110001;
        10'b01100110: data <= 20'b10010000111001110000;
        10'b01100111: data <= 20'b10101100100010100010;
        10'b01101000: data <= 20'b00110000000010111011;
        10'b01101001: data <= 20'b00011100110010011011;
        10'b01101010: data <= 20'b00101000110010010010;
        10'b01101011: data <= 20'b00100101001010011001;
        10'b01101100: data <= 20'b00100001000010110110;
        10'b01101101: data <= 20'b10101000011010001011;
        10'b01101110: data <= 20'b10010000111010010010;
        10'b01101111: data <= 20'b10100110111010000100;
        10'b01110000: data <= 20'b10101100000001110110;
        10'b01110001: data <= 20'b00101000100010101001;
        10'b01110010: data <= 20'b10101010100010011101;
        10'b01110011: data <= 20'b10010000110001011000;
        10'b01110100: data <= 20'b00101010110010111001;
        10'b01110101: data <= 20'b10101110010010111001;
        10'b01110110: data <= 20'b10000001001010100011;
        10'b01110111: data <= 20'b10101001000010101101;
        10'b01111000: data <= 20'b00101001011010110011;
        10'b01111001: data <= 20'b00100100000010011101;
        10'b01111010: data <= 20'b10100110001010010100;
        10'b01111011: data <= 20'b10100100110010011110;
        10'b01111100: data <= 20'b00100101000010101110;
        10'b01111101: data <= 20'b10101001111010100110;
        10'b01111110: data <= 20'b00110000100011001011;
        10'b01111111: data <= 20'b10110000001010000101;
        10'b10000000: data <= 20'b00100100111010110010;
        10'b10000001: data <= 20'b10101010101010010001;
        10'b10000010: data <= 20'b00101000011011000101;
        10'b10000011: data <= 20'b00100101111010011111;
        10'b10000100: data <= 20'b00101001100010011110;
        10'b10000101: data <= 20'b00110100011010100000;
        10'b10000110: data <= 20'b10110001101001011100;
        10'b10000111: data <= 20'b10101110011011010100;
        10'b10001000: data <= 20'b10101101011011000101;
        10'b10001001: data <= 20'b00101110000010010010;
        10'b10001010: data <= 20'b10100101101010001010;
        10'b10001011: data <= 20'b10100011000010000011;
        10'b10001100: data <= 20'b00101010100010100000;
        10'b10001101: data <= 20'b10100110111011001100;
        10'b10001110: data <= 20'b00100101010010100111;
        10'b10001111: data <= 20'b10101110010010110011;
        10'b10010000: data <= 20'b00101100101010011110;
        10'b10010001: data <= 20'b10101010010010100101;
        10'b10010010: data <= 20'b10101101011011011001;
        10'b10010011: data <= 20'b10101100110010101101;
        10'b10010100: data <= 20'b10100010011010111100;
        10'b10010101: data <= 20'b10100111011010010101;
        10'b10010110: data <= 20'b10100111110010110001;
        10'b10010111: data <= 20'b10100100011011000111;
        10'b10011000: data <= 20'b10100001111010101110;
        10'b10011001: data <= 20'b10101101111010101111;
        10'b10011010: data <= 20'b00101111010010001111;
        10'b10011011: data <= 20'b00101101101010100110;
        10'b10011100: data <= 20'b00100111100010010111;
        10'b10011101: data <= 20'b10101100101010000010;
        10'b10011110: data <= 20'b10101100000010001011;
        10'b10011111: data <= 20'b00110000010010001000;
        10'b10100000: data <= 20'b00101001001001100100;
        10'b10100001: data <= 20'b00100101110010101100;
        10'b10100010: data <= 20'b00100000101010110110;
        10'b10100011: data <= 20'b00101010100010101001;
        10'b10100100: data <= 20'b10101100101010011001;
        10'b10100101: data <= 20'b10101101100011000001;
        10'b10100110: data <= 20'b10101000101010111010;
        10'b10100111: data <= 20'b10101001101001010111;
        10'b10101000: data <= 20'b10101111000011000011;
        10'b10101001: data <= 20'b10101011110010010000;
        10'b10101010: data <= 20'b10011100001010001010;
        10'b10101011: data <= 20'b00101100001010011000;
        10'b10101100: data <= 20'b00101011010010001010;
        10'b10101101: data <= 20'b10101101100010110111;
        10'b10101110: data <= 20'b00101110101011000100;
        10'b10101111: data <= 20'b00101100001010110000;
        10'b10110000: data <= 20'b10101101111010110101;
        10'b10110001: data <= 20'b00100100001010010001;
        10'b10110010: data <= 20'b10100110110010110001;
        10'b10110011: data <= 20'b10101100111011000011;
        10'b10110100: data <= 20'b00100111101011000001;
        10'b10110101: data <= 20'b10101011111010011100;
        10'b10110110: data <= 20'b00101010001001010000;
        10'b10110111: data <= 20'b00110011011011010011;
        10'b10111000: data <= 20'b10100010000010100011;
        10'b10111001: data <= 20'b00110000111011000001;
        10'b10111010: data <= 20'b00100101111010101111;
        10'b10111011: data <= 20'b10101111010010110111;
        10'b10111100: data <= 20'b10101001001010101011;
        10'b10111101: data <= 20'b00101010011010110011;
        10'b10111110: data <= 20'b10101011001010001010;
        10'b10111111: data <= 20'b10101010100010110110;
        10'b11000000: data <= 20'b10100011110010010101;
        10'b11000001: data <= 20'b00101100001010011101;
        10'b11000010: data <= 20'b00101100110010110011;
        10'b11000011: data <= 20'b10100100011011100110;
        10'b11000100: data <= 20'b10101101010011010011;
        10'b11000101: data <= 20'b10100111000010010000;
        10'b11000110: data <= 20'b10101100000010111001;
        10'b11000111: data <= 20'b10101010010010101001;
        10'b11001000: data <= 20'b10101010111010100010;
        10'b11001001: data <= 20'b10011110001010100000;
        10'b11001010: data <= 20'b00100001110010100100;
        10'b11001011: data <= 20'b00100111110010011011;
        10'b11001100: data <= 20'b10100101000010011100;
        10'b11001101: data <= 20'b00101101010010111010;
        10'b11001110: data <= 20'b00100100110010101001;
        10'b11001111: data <= 20'b00110000111010100011;
        10'b11010000: data <= 20'b00110010001011010001;
        10'b11010001: data <= 20'b00100000111010110001;
        10'b11010010: data <= 20'b00100101000010100110;
        10'b11010011: data <= 20'b00110011011010110010;
        10'b11010100: data <= 20'b00101010100010110001;
        10'b11010101: data <= 20'b00110001001011000000;
        10'b11010110: data <= 20'b10100100110010010010;
        10'b11010111: data <= 20'b00101111010011000100;
        10'b11011000: data <= 20'b00100001010010110111;
        10'b11011001: data <= 20'b00101100011010000000;
        10'b11011010: data <= 20'b00110000111010111110;
        10'b11011011: data <= 20'b10100100110010110100;
        10'b11011100: data <= 20'b00100001011010110110;
        10'b11011101: data <= 20'b10101110001010110010;
        10'b11011110: data <= 20'b10101101001010000001;
        10'b11011111: data <= 20'b10110001100010111100;
        10'b11100000: data <= 20'b10101001111010111100;
        10'b11100001: data <= 20'b00101011001010100001;
        10'b11100010: data <= 20'b00100100010001110100;
        10'b11100011: data <= 20'b10100011000010111100;
        10'b11100100: data <= 20'b10011110000010011000;
        10'b11100101: data <= 20'b00010101100010110000;
        10'b11100110: data <= 20'b00101000001010001110;
        10'b11100111: data <= 20'b10100100110010101001;
        10'b11101000: data <= 20'b00100010101010110001;
        10'b11101001: data <= 20'b00100100110010111011;
        10'b11101010: data <= 20'b10100110111010100001;
        10'b11101011: data <= 20'b00100001110010010001;
        10'b11101100: data <= 20'b00011010000010100011;
        10'b11101101: data <= 20'b10100010100010011011;
        10'b11101110: data <= 20'b10101101000010100110;
        10'b11101111: data <= 20'b10011001000001110110;
        10'b11110000: data <= 20'b10101000110010100010;
        10'b11110001: data <= 20'b10101101010011000111;
        10'b11110010: data <= 20'b10101001010010100000;
        10'b11110011: data <= 20'b00110100001010110101;
        10'b11110100: data <= 20'b00101001111010110011;
        10'b11110101: data <= 20'b10101101011010110111;
        10'b11110110: data <= 20'b00100111000010011110;
        10'b11110111: data <= 20'b10101010111010111101;
        10'b11111000: data <= 20'b00101100110010000111;
        10'b11111001: data <= 20'b00101110011010010111;
        10'b11111010: data <= 20'b10100100000001111010;
        10'b11111011: data <= 20'b00100101000010110100;
        10'b11111100: data <= 20'b10100101000011010010;
        10'b11111101: data <= 20'b10100111001010010101;
        10'b11111110: data <= 20'b00100110000010011010;
        10'b11111111: data <= 20'b10110101000011010111;
        10'b100000000: data <= 20'b00101011000001110111;
        10'b100000001: data <= 20'b10101100101010101011;
        10'b100000010: data <= 20'b00101000101010101010;
        10'b100000011: data <= 20'b10101100011011000000;
        10'b100000100: data <= 20'b00100111100010011010;
        10'b100000101: data <= 20'b10100110100011000000;
        10'b100000110: data <= 20'b00101100000010100000;
        10'b100000111: data <= 20'b00101001001010011001;
        10'b100001000: data <= 20'b00100010000010010011;
        10'b100001001: data <= 20'b10101000000011001011;
        10'b100001010: data <= 20'b00110000000010111101;
        10'b100001011: data <= 20'b10101111001010111100;
        10'b100001100: data <= 20'b10101100010010110001;
        10'b100001101: data <= 20'b00101010001010001001;
        10'b100001110: data <= 20'b00010011100010010111;
        10'b100001111: data <= 20'b10101111100010111101;
        10'b100010000: data <= 20'b10101100101010110100;
        10'b100010001: data <= 20'b10100011001010010010;
        10'b100010010: data <= 20'b00101101000010011001;
        10'b100010011: data <= 20'b10100001010010100100;
        10'b100010100: data <= 20'b10101000000010101101;
        10'b100010101: data <= 20'b00100111000010011011;
        10'b100010110: data <= 20'b10101010100011000001;
        10'b100010111: data <= 20'b00101001101010101011;
        10'b100011000: data <= 20'b00101111101010110101;
        10'b100011001: data <= 20'b10101000110010000001;
        10'b100011010: data <= 20'b10100111001010011110;
        10'b100011011: data <= 20'b10111001000011111011;
        10'b100011100: data <= 20'b00011100110011000010;
        10'b100011101: data <= 20'b10101000111010011001;
        10'b100011110: data <= 20'b10101100110010011100;
        10'b100011111: data <= 20'b10100101010010001001;
        10'b100100000: data <= 20'b10100001100010110011;
        10'b100100001: data <= 20'b00011010111010100111;
        10'b100100010: data <= 20'b10101100000010111111;
        10'b100100011: data <= 20'b10101010111001011010;
        10'b100100100: data <= 20'b10100000000010000110;
        10'b100100101: data <= 20'b00101111110010101000;
        10'b100100110: data <= 20'b00101101111010101011;
        10'b100100111: data <= 20'b10100010011010101110;
        10'b100101000: data <= 20'b00100011000001011011;
        10'b100101001: data <= 20'b10101001100001001000;
        10'b100101010: data <= 20'b00101110100011000010;
        10'b100101011: data <= 20'b00110000110010011110;
        10'b100101100: data <= 20'b00101011001010110101;
        10'b100101101: data <= 20'b00011101111010100010;
        10'b100101110: data <= 20'b10101001100001101110;
        10'b100101111: data <= 20'b00101110100011000010;
        10'b100110000: data <= 20'b00100001011010100001;
        10'b100110001: data <= 20'b00110100000011101001;
        10'b100110010: data <= 20'b00101110011010110011;
        10'b100110011: data <= 20'b10101000111010100111;
        10'b100110100: data <= 20'b00011010001000001111;
        10'b100110101: data <= 20'b00101001000010011111;
        10'b100110110: data <= 20'b10100010000010100111;
        10'b100110111: data <= 20'b00100001110010010100;
        10'b100111000: data <= 20'b00101101010010101011;
        10'b100111001: data <= 20'b00101000010010011101;
        10'b100111010: data <= 20'b10101100000010110101;
        10'b100111011: data <= 20'b00100011001010110000;
        10'b100111100: data <= 20'b00101111011011000100;
        10'b100111101: data <= 20'b10111001001011001011;
        10'b100111110: data <= 20'b10101000111010110010;
        10'b100111111: data <= 20'b10101011101010100011;
        10'b101000000: data <= 20'b10100010000001000010;
        10'b101000001: data <= 20'b00100111010010101101;
        10'b101000010: data <= 20'b10100010100001101100;
        10'b101000011: data <= 20'b10100101000010000010;
        10'b101000100: data <= 20'b00101010000010101110;
        10'b101000101: data <= 20'b00111000101011011011;
        10'b101000110: data <= 20'b00101011001010000011;
        10'b101000111: data <= 20'b00100001011010100010;
        10'b101001000: data <= 20'b00101101000010110010;
        10'b101001001: data <= 20'b00101001111010100100;
        10'b101001010: data <= 20'b00101000100010101110;
        10'b101001011: data <= 20'b00101010011010000100;
        10'b101001100: data <= 20'b00100000010010110100;
        10'b101001101: data <= 20'b00110010001011000110;
        10'b101001110: data <= 20'b00011100110010011000;
        10'b101001111: data <= 20'b00101001000010111100;
        10'b101010000: data <= 20'b00100010100010111110;
        10'b101010001: data <= 20'b10100010101001111101;
        10'b101010010: data <= 20'b00010000110010110101;
        10'b101010011: data <= 20'b10101000111001100110;
        10'b101010100: data <= 20'b10100100001011000111;
        10'b101010101: data <= 20'b10101011011011000011;
        10'b101010110: data <= 20'b10110100101010111111;
        10'b101010111: data <= 20'b00100101111010101000;
        10'b101011000: data <= 20'b00110000111010101001;
        10'b101011001: data <= 20'b00100100010010000011;
        10'b101011010: data <= 20'b00101101000010101011;
        10'b101011011: data <= 20'b00101111110010110101;
        10'b101011100: data <= 20'b10101011001011000100;
        10'b101011101: data <= 20'b10101000111010110110;
        10'b101011110: data <= 20'b10101011000010110001;
        10'b101011111: data <= 20'b10101000100010011000;
        10'b101100000: data <= 20'b10101101011010100010;
        10'b101100001: data <= 20'b10011101100001011011;
        10'b101100010: data <= 20'b10101010000010111011;
        10'b101100011: data <= 20'b10100101111010110001;
        10'b101100100: data <= 20'b10011000011010100000;
        10'b101100101: data <= 20'b10100101010010100000;
        10'b101100110: data <= 20'b00100111010010100100;
        10'b101100111: data <= 20'b10101011111001011100;
        10'b101101000: data <= 20'b00101000000010010011;
        10'b101101001: data <= 20'b10100100000010001111;
        10'b101101010: data <= 20'b10110101100010100100;
        10'b101101011: data <= 20'b00110011011011000001;
        10'b101101100: data <= 20'b00101001111010101100;
        10'b101101101: data <= 20'b10100100001010011000;
        10'b101101110: data <= 20'b10101000110010110110;
        10'b101101111: data <= 20'b00101001011010100010;
        10'b101110000: data <= 20'b10100110110010011111;
        10'b101110001: data <= 20'b10101101000001010100;
        10'b101110010: data <= 20'b00110100000011100001;
        10'b101110011: data <= 20'b10101010101010010101;
        10'b101110100: data <= 20'b10101110000010111101;
        10'b101110101: data <= 20'b00100100101010011101;
        10'b101110110: data <= 20'b00011101000010011110;
        10'b101110111: data <= 20'b10101001100010101111;
        10'b101111000: data <= 20'b00110111111011100000;
        10'b101111001: data <= 20'b10100101011001101000;
        10'b101111010: data <= 20'b10101011000001111000;
        10'b101111011: data <= 20'b00101001001001111111;
        10'b101111100: data <= 20'b00101010110010111110;
        10'b101111101: data <= 20'b10101000001010001110;
        10'b101111110: data <= 20'b00110010000011000110;
        10'b101111111: data <= 20'b00101101111010101010;
        10'b110000000: data <= 20'b10110000100010011101;
        10'b110000001: data <= 20'b00100000011010101100;
        10'b110000010: data <= 20'b00100010000010010010;
        10'b110000011: data <= 20'b00100110010010001001;
        10'b110000100: data <= 20'b00010001100010000101;
        10'b110000101: data <= 20'b10100101010010011000;
        10'b110000110: data <= 20'b00110111001011011001;
        10'b110000111: data <= 20'b00011010101010101011;
        10'b110001000: data <= 20'b10101110110010110011;
        10'b110001001: data <= 20'b00101011010001111101;
        10'b110001010: data <= 20'b00100000011010001011;
        10'b110001011: data <= 20'b10101010111001101110;
        10'b110001100: data <= 20'b00101100110010101101;
        10'b110001101: data <= 20'b10110001100010111000;
        10'b110001110: data <= 20'b10101101010001111010;
        10'b110001111: data <= 20'b00101110100011001010;
        10'b110010000: data <= 20'b10101000101010110010;
        10'b110010001: data <= 20'b00100010111010110010;
        10'b110010010: data <= 20'b00101000111010100101;
        10'b110010011: data <= 20'b00110001010010100111;
        10'b110010100: data <= 20'b10100001100001110000;
        10'b110010101: data <= 20'b10101011100010110010;
        10'b110010110: data <= 20'b00101010110001111111;
        10'b110010111: data <= 20'b10101011010010101111;
        10'b110011000: data <= 20'b10110000011010011000;
        10'b110011001: data <= 20'b00101001001010100100;
        10'b110011010: data <= 20'b00101101001010100110;
        10'b110011011: data <= 20'b00101010100010011011;
        10'b110011100: data <= 20'b00100011010010100100;
        10'b110011101: data <= 20'b10100101100010100001;
        10'b110011110: data <= 20'b10101010100010110011;
        10'b110011111: data <= 20'b10101010101010101000;
        10'b110100000: data <= 20'b00100110001010011101;
        10'b110100001: data <= 20'b10110001010011000011;
        10'b110100010: data <= 20'b00100011101010001000;
        10'b110100011: data <= 20'b00101101000010110101;
        10'b110100100: data <= 20'b10110000000010110101;
        10'b110100101: data <= 20'b10100011101001111000;
        10'b110100110: data <= 20'b10101000100010110111;
        10'b110100111: data <= 20'b00100110101010101110;
        10'b110101000: data <= 20'b00110110111011010000;
        10'b110101001: data <= 20'b00110010011010111100;
        10'b110101010: data <= 20'b10101001001010001010;
        10'b110101011: data <= 20'b10110100101011001110;
        10'b110101100: data <= 20'b10100111111010111010;
        10'b110101101: data <= 20'b00101101111010000011;
        10'b110101110: data <= 20'b10101100000000000011;
        10'b110101111: data <= 20'b10101101010011000010;
        10'b110110000: data <= 20'b00101000011010011100;
        10'b110110001: data <= 20'b00100110010010010111;
        10'b110110010: data <= 20'b00100110110010100001;
        10'b110110011: data <= 20'b10100111000010100110;
        10'b110110100: data <= 20'b10100101111010001011;
        10'b110110101: data <= 20'b00101111010010111110;
        10'b110110110: data <= 20'b00100111101010010011;
        10'b110110111: data <= 20'b00101011000011000001;
        10'b110111000: data <= 20'b10111100011011010011;
        10'b110111001: data <= 20'b10101110101010110101;
        10'b110111010: data <= 20'b00101011001010101011;
        10'b110111011: data <= 20'b00100001001010100110;
        10'b110111100: data <= 20'b10010000111010010011;
        10'b110111101: data <= 20'b10110010010011000101;
        10'b110111110: data <= 20'b00101010100010110110;
        10'b110111111: data <= 20'b10101101110010110101;
        10'b111000000: data <= 20'b10110000001011001011;
        10'b111000001: data <= 20'b10101010010001111110;
        10'b111000010: data <= 20'b10110001010011011110;
        10'b111000011: data <= 20'b00101011011010110101;
        10'b111000100: data <= 20'b00100111010010100000;
        10'b111000101: data <= 20'b10110110010011010001;
        10'b111000110: data <= 20'b10010010110010010001;
        10'b111000111: data <= 20'b00100110100001111101;
        10'b111001000: data <= 20'b00011111000010101101;
        10'b111001001: data <= 20'b10101001000001100001;
        10'b111001010: data <= 20'b00011010110001100001;
        10'b111001011: data <= 20'b00100111000010110111;
        10'b111001100: data <= 20'b10100100100001010010;
        10'b111001101: data <= 20'b00110011100010011010;
        10'b111001110: data <= 20'b10101111111010110011;
        10'b111001111: data <= 20'b00110110001010110001;
        10'b111010000: data <= 20'b00100100101010110000;
        10'b111010001: data <= 20'b10101001100010110111;
        10'b111010010: data <= 20'b10100110001010010011;
        10'b111010011: data <= 20'b00100111100010000001;
        10'b111010100: data <= 20'b00110101000011010011;
        10'b111010101: data <= 20'b00011010101010000001;
        10'b111010110: data <= 20'b10100110000010011010;
        10'b111010111: data <= 20'b10011001010010011011;
        10'b111011000: data <= 20'b00101110101001110010;
        10'b111011001: data <= 20'b00100111100010000111;
        10'b111011010: data <= 20'b00100101000011000011;
        10'b111011011: data <= 20'b00100000100010101110;
        10'b111011100: data <= 20'b00100001000010010011;
        10'b111011101: data <= 20'b10100010000010101001;
        10'b111011110: data <= 20'b00110000101010101110;
        10'b111011111: data <= 20'b10101100001010110001;
        10'b111100000: data <= 20'b00110011111011001100;
        10'b111100001: data <= 20'b00100001011010010000;
        10'b111100010: data <= 20'b10101101100010101011;
        10'b111100011: data <= 20'b00101001011001110001;
        10'b111100100: data <= 20'b00101010110011000010;
        10'b111100101: data <= 20'b10101000100010100111;
        10'b111100110: data <= 20'b10011000100011010010;
        10'b111100111: data <= 20'b10011001011010001001;
        10'b111101000: data <= 20'b10100101010010111110;
        10'b111101001: data <= 20'b10100111111010101101;
        10'b111101010: data <= 20'b10011110011011000000;
        10'b111101011: data <= 20'b00101011100001110101;
        10'b111101100: data <= 20'b10101010111010000001;
        10'b111101101: data <= 20'b00100001111010001010;
        10'b111101110: data <= 20'b00100100000010110000;
        10'b111101111: data <= 20'b10100111101010101010;
        10'b111110000: data <= 20'b00101001101010101001;
        10'b111110001: data <= 20'b10011100001010100101;
        10'b111110010: data <= 20'b10101100011011010110;
        10'b111110011: data <= 20'b10101100100001100011;
        10'b111110100: data <= 20'b00010111000010011010;
        10'b111110101: data <= 20'b00101101010010100101;
        10'b111110110: data <= 20'b00101011000010010100;
        10'b111110111: data <= 20'b10101001101010011011;
        10'b111111000: data <= 20'b00100110111010100101;
        10'b111111001: data <= 20'b00110001001010110110;
        10'b111111010: data <= 20'b10110000000010110111;
        10'b111111011: data <= 20'b10100010111010111010;
        10'b111111100: data <= 20'b00101110011010110010;
        10'b111111101: data <= 20'b10101110110011000100;
        10'b111111110: data <= 20'b00011101101001111101;
        10'b111111111: data <= 20'b00100000000010101111;
        10'b1000000000: data <= 20'b10100110111010001100;
        10'b1000000001: data <= 20'b10101010101010011101;
        10'b1000000010: data <= 20'b00101011100001010010;
        10'b1000000011: data <= 20'b10101011010010100111;
        10'b1000000100: data <= 20'b00101001101001111000;
        10'b1000000101: data <= 20'b10100110110010110000;
        10'b1000000110: data <= 20'b10101000001001101011;
        10'b1000000111: data <= 20'b10100110111010111111;
        10'b1000001000: data <= 20'b00101000001010101011;
        10'b1000001001: data <= 20'b10101000110010101010;
        10'b1000001010: data <= 20'b10011111101010100111;
        10'b1000001011: data <= 20'b10101101110001110001;
        10'b1000001100: data <= 20'b10101101100010110101;
        10'b1000001101: data <= 20'b10100011100010010000;
        10'b1000001110: data <= 20'b00101010110011000000;
        10'b1000001111: data <= 20'b00101001001010011011;
        10'b1000010000: data <= 20'b00100010011011100011;
        10'b1000010001: data <= 20'b00011100100010001010;
        10'b1000010010: data <= 20'b00100100000010111001;
        10'b1000010011: data <= 20'b10100011111011000100;
        10'b1000010100: data <= 20'b00110000101011001000;
        10'b1000010101: data <= 20'b10011010001010100111;
        10'b1000010110: data <= 20'b10110100110010000010;
        10'b1000010111: data <= 20'b00100110001010110010;
        10'b1000011000: data <= 20'b00010011000010010000;
        10'b1000011001: data <= 20'b10101000011001011010;
        10'b1000011010: data <= 20'b10010001010011000011;
        10'b1000011011: data <= 20'b00011010101010101110;
        10'b1000011100: data <= 20'b00011111000011000100;
        10'b1000011101: data <= 20'b10011110111010001000;
        10'b1000011110: data <= 20'b10100000000010110101;
        10'b1000011111: data <= 20'b10101011000001001110;
        10'b1000100000: data <= 20'b10110001011001100101;
        10'b1000100001: data <= 20'b10101010011011010100;
        10'b1000100010: data <= 20'b10011111001010110001;
        10'b1000100011: data <= 20'b00100010110001111100;
        10'b1000100100: data <= 20'b10100000010010110000;
        10'b1000100101: data <= 20'b00101100011010101111;
        10'b1000100110: data <= 20'b10110001100010100100;
        10'b1000100111: data <= 20'b00101100111010110100;
        10'b1000101000: data <= 20'b10110000010011000101;
        10'b1000101001: data <= 20'b10101111111010110010;
        10'b1000101010: data <= 20'b10100101001010000101;
        10'b1000101011: data <= 20'b10100100110010011101;
        10'b1000101100: data <= 20'b00110001010010110001;
        10'b1000101101: data <= 20'b10101010010010000010;
        10'b1000101110: data <= 20'b00100010010010010101;
        10'b1000101111: data <= 20'b10101011110010000000;
        10'b1000110000: data <= 20'b10100100000010001011;
        10'b1000110001: data <= 20'b10101011110010111111;
        10'b1000110010: data <= 20'b00101100111010000101;
        10'b1000110011: data <= 20'b00110000000010011001;
        10'b1000110100: data <= 20'b10101011001010101000;
        10'b1000110101: data <= 20'b10101100011010010110;
        10'b1000110110: data <= 20'b00101100010001111111;
        10'b1000110111: data <= 20'b00101110011010110010;
        10'b1000111000: data <= 20'b10101010011010100111;
        10'b1000111001: data <= 20'b10101011110010110010;
        10'b1000111010: data <= 20'b10100100101010101101;
        10'b1000111011: data <= 20'b00101000000010100110;
        10'b1000111100: data <= 20'b00100100000010111101;
        10'b1000111101: data <= 20'b10100000011010100110;
        10'b1000111110: data <= 20'b00100011111010100111;
        10'b1000111111: data <= 20'b00110001011011011011;
        10'b1001000000: data <= 20'b10101100010010101101;
        10'b1001000001: data <= 20'b10101110100010011000;
        10'b1001000010: data <= 20'b10011111101010110011;
        10'b1001000011: data <= 20'b10101011101010010101;
        10'b1001000100: data <= 20'b10100101000010111110;
        10'b1001000101: data <= 20'b10101000001010011111;
        10'b1001000110: data <= 20'b10110000010011000000;
        10'b1001000111: data <= 20'b10110000001011001110;
        10'b1001001000: data <= 20'b00011000101010101010;
        10'b1001001001: data <= 20'b10101101011010010101;
        10'b1001001010: data <= 20'b10110101111011000000;
        10'b1001001011: data <= 20'b10011101011010010110;
        10'b1001001100: data <= 20'b10101001100010011110;
        10'b1001001101: data <= 20'b00110000100011000010;
        10'b1001001110: data <= 20'b00110010101011001001;
        10'b1001001111: data <= 20'b10101111101010100101;
        10'b1001010000: data <= 20'b00101111011001110011;
        10'b1001010001: data <= 20'b00100010111010100001;
        10'b1001010010: data <= 20'b00100000010010101010;
        10'b1001010011: data <= 20'b00101001000010000011;
        10'b1001010100: data <= 20'b10101010010010001011;
        10'b1001010101: data <= 20'b00011011000010010000;
        10'b1001010110: data <= 20'b00001011010010110001;
        10'b1001010111: data <= 20'b00100110111010100011;
        10'b1001011000: data <= 20'b00110001000011001011;
        10'b1001011001: data <= 20'b10110000000010111000;
        10'b1001011010: data <= 20'b10110110101001110001;
        10'b1001011011: data <= 20'b10101110011010010011;
        10'b1001011100: data <= 20'b10101111111010010111;
        10'b1001011101: data <= 20'b10101110000010010111;
        10'b1001011110: data <= 20'b10101011011010110011;
        10'b1001011111: data <= 20'b00100001101010110001;
        10'b1001100000: data <= 20'b10100000011010111001;
        10'b1001100001: data <= 20'b00100111011010110010;
        10'b1001100010: data <= 20'b10101101011010100010;
        10'b1001100011: data <= 20'b00101101000010010001;
        10'b1001100100: data <= 20'b00010010110010100011;
        10'b1001100101: data <= 20'b00101000001010110001;
        10'b1001100110: data <= 20'b10101100001011000100;
        10'b1001100111: data <= 20'b00110100011011001100;
        10'b1001101000: data <= 20'b00100011011010110101;
        10'b1001101001: data <= 20'b10101100011010000100;
        10'b1001101010: data <= 20'b10101100001010010001;
        10'b1001101011: data <= 20'b00011111111001100000;
        10'b1001101100: data <= 20'b10110010110011000010;
        10'b1001101101: data <= 20'b00101010110010001111;
        10'b1001101110: data <= 20'b00100001011010010001;
        10'b1001101111: data <= 20'b00101101010010111110;
        10'b1001110000: data <= 20'b00110100000011010010;
        10'b1001110001: data <= 20'b00101000011010000000;
        10'b1001110010: data <= 20'b00100110010010011001;
        10'b1001110011: data <= 20'b10101100101000110010;
        10'b1001110100: data <= 20'b10110000100010100111;
        10'b1001110101: data <= 20'b00101100000010011110;
        10'b1001110110: data <= 20'b00101000111010011001;
        10'b1001110111: data <= 20'b00101011010010110111;
        10'b1001111000: data <= 20'b10100110000010011011;
        10'b1001111001: data <= 20'b10011100010010110011;
        10'b1001111010: data <= 20'b00110011011011000100;
        10'b1001111011: data <= 20'b10100011000010010000;
        10'b1001111100: data <= 20'b00100111000010100111;
        10'b1001111101: data <= 20'b10101100010010011011;
        10'b1001111110: data <= 20'b00110010100011001000;
        10'b1001111111: data <= 20'b10101101111010111001;
        10'b1010000000: data <= 20'b00101010011010100011;
        10'b1010000001: data <= 20'b00100100011010011111;
        10'b1010000010: data <= 20'b10101000101010010010;
        10'b1010000011: data <= 20'b00101000000010010010;
        10'b1010000100: data <= 20'b10101110101011010010;
        10'b1010000101: data <= 20'b00110001101011011000;
        10'b1010000110: data <= 20'b00101100111001111000;
        10'b1010000111: data <= 20'b00100111001010000111;
        10'b1010001000: data <= 20'b10101000101010000100;
        10'b1010001001: data <= 20'b00101100110010011010;
        10'b1010001010: data <= 20'b00101101000010000010;
        10'b1010001011: data <= 20'b10101011100010011010;
        10'b1010001100: data <= 20'b00101011101010110101;
        10'b1010001101: data <= 20'b00100000011010000111;
        10'b1010001110: data <= 20'b00011111110010011010;
        10'b1010001111: data <= 20'b00101100100010110101;
        10'b1010010000: data <= 20'b00110010110010100000;
        10'b1010010001: data <= 20'b00100100111010100001;
        10'b1010010010: data <= 20'b00011110100010101010;
        10'b1010010011: data <= 20'b10100100110010110100;
        10'b1010010100: data <= 20'b00100101000010000111;
        10'b1010010101: data <= 20'b00101011110010110101;
        10'b1010010110: data <= 20'b00010100111010011000;
        10'b1010010111: data <= 20'b00101010010010001101;
        10'b1010011000: data <= 20'b00101111000010100110;
        10'b1010011001: data <= 20'b00101110011011011001;
        10'b1010011010: data <= 20'b00101010001010110001;
        10'b1010011011: data <= 20'b00101000111001111010;
        10'b1010011100: data <= 20'b00101001110010001011;
        10'b1010011101: data <= 20'b00100110100010010111;
        10'b1010011110: data <= 20'b00100110100010100010;
        10'b1010011111: data <= 20'b10101100000010101110;
        10'b1010100000: data <= 20'b10011101001010100001;
        10'b1010100001: data <= 20'b00010111000001100101;
        10'b1010100010: data <= 20'b10100011110011000001;
        10'b1010100011: data <= 20'b00101101111011000000;
        10'b1010100100: data <= 20'b10100101101010110001;
        10'b1010100101: data <= 20'b10100000010010011001;
        10'b1010100110: data <= 20'b00101100000010110001;
        10'b1010100111: data <= 20'b00101010101011000101;
        10'b1010101000: data <= 20'b10011001101010110001;
        10'b1010101001: data <= 20'b10110000110010010001;
        10'b1010101010: data <= 20'b10100001101011110001;
        10'b1010101011: data <= 20'b00010100101010111111;
        10'b1010101100: data <= 20'b10101100111011001010;
        10'b1010101101: data <= 20'b00011101011010001011;
        10'b1010101110: data <= 20'b10101001001010011110;
        10'b1010101111: data <= 20'b10101000010010011110;
        10'b1010110000: data <= 20'b10100010110010101110;
        10'b1010110001: data <= 20'b00101101101010100110;
        10'b1010110010: data <= 20'b00101011010010110100;
        10'b1010110011: data <= 20'b00100000110010101000;
        10'b1010110100: data <= 20'b00100100100010111011;
        10'b1010110101: data <= 20'b00101000101010010111;
        10'b1010110110: data <= 20'b00101000111010000011;
        10'b1010110111: data <= 20'b10110000100010110100;
        10'b1010111000: data <= 20'b00101110111010110010;
        10'b1010111001: data <= 20'b00100001101010010100;
        10'b1010111010: data <= 20'b10101100000010011001;
        10'b1010111011: data <= 20'b10101011101010111111;
        10'b1010111100: data <= 20'b00101011011010001011;
        10'b1010111101: data <= 20'b10101000011010001111;
        10'b1010111110: data <= 20'b10101101100011000110;
        10'b1010111111: data <= 20'b00101001000010011001;
        10'b1011000000: data <= 20'b00110001000010110100;
        10'b1011000001: data <= 20'b00101100011010011101;
        10'b1011000010: data <= 20'b00101000101010100100;
        10'b1011000011: data <= 20'b10110111111011010111;
        10'b1011000100: data <= 20'b10101001101010111011;
        10'b1011000101: data <= 20'b10101010111010110011;
        10'b1011000110: data <= 20'b10100010011010100001;
        10'b1011000111: data <= 20'b10110001011011010001;
        10'b1011001000: data <= 20'b00101000100010011111;
        10'b1011001001: data <= 20'b00101010000001110101;
        10'b1011001010: data <= 20'b00011111110011001100;
        10'b1011001011: data <= 20'b00101100011010110100;
        10'b1011001100: data <= 20'b00100011101010000110;
        10'b1011001101: data <= 20'b10110000110011010000;
        10'b1011001110: data <= 20'b10100001111010101110;
        10'b1011001111: data <= 20'b00101011111010001001;
        10'b1011010000: data <= 20'b00101110100010101001;
        10'b1011010001: data <= 20'b00101110101010110010;
        10'b1011010010: data <= 20'b00101011111010011100;
        10'b1011010011: data <= 20'b00011111010010110011;
        10'b1011010100: data <= 20'b00110001100010110000;
        10'b1011010101: data <= 20'b00101001000010010110;
        10'b1011010110: data <= 20'b00101001100010000010;
        10'b1011010111: data <= 20'b10100110100010100001;
        10'b1011011000: data <= 20'b00100010110010001001;
        10'b1011011001: data <= 20'b10011111000010011010;
        10'b1011011010: data <= 20'b10100000000010010001;
        10'b1011011011: data <= 20'b10011001100010011011;
        10'b1011011100: data <= 20'b10100011011010100111;
        10'b1011011101: data <= 20'b00101010010010011001;
        10'b1011011110: data <= 20'b10110011100010100001;
        10'b1011011111: data <= 20'b10101111001010110101;
        10'b1011100000: data <= 20'b10100100011010000110;
        10'b1011100001: data <= 20'b10101001000010011110;
        10'b1011100010: data <= 20'b00011110100010011101;
        10'b1011100011: data <= 20'b10100101110010101111;
        10'b1011100100: data <= 20'b00101011011001100101;
        10'b1011100101: data <= 20'b10101100111010110100;
        10'b1011100110: data <= 20'b00110010111010100001;
        10'b1011100111: data <= 20'b10100111001001010100;
        10'b1011101000: data <= 20'b00101001100011000100;
        10'b1011101001: data <= 20'b10011110101010011111;
        10'b1011101010: data <= 20'b10101000010010110001;
        10'b1011101011: data <= 20'b00011110000001100111;
        10'b1011101100: data <= 20'b10101100011010111010;
        10'b1011101101: data <= 20'b10100000000010100001;
        10'b1011101110: data <= 20'b10011101010010110001;
        10'b1011101111: data <= 20'b00100101010010100110;
        10'b1011110000: data <= 20'b00101000010010010101;
        10'b1011110001: data <= 20'b10101011110010100000;
        10'b1011110010: data <= 20'b00100111101010100010;
        10'b1011110011: data <= 20'b10101100100010110100;
        10'b1011110100: data <= 20'b10100001111010111100;
        10'b1011110101: data <= 20'b00101000001010101011;
        10'b1011110110: data <= 20'b00101001011010001011;
        10'b1011110111: data <= 20'b00110000110010101001;
        10'b1011111000: data <= 20'b10100101000010100000;
        10'b1011111001: data <= 20'b00101001101010010101;
        10'b1011111010: data <= 20'b10100110110001111100;
        10'b1011111011: data <= 20'b00100011000010110101;
        10'b1011111100: data <= 20'b00100101000010001100;
        10'b1011111101: data <= 20'b10101100010010101001;
        10'b1011111110: data <= 20'b10100000001010011000;
        10'b1011111111: data <= 20'b00100110101010001101;
        10'b1100000000: data <= 20'b10101100110011010001;
        10'b1100000001: data <= 20'b10101000001011001000;
        10'b1100000010: data <= 20'b00100100111010000100;
        10'b1100000011: data <= 20'b00100100100010100001;
        10'b1100000100: data <= 20'b00100110110001110111;
        10'b1100000101: data <= 20'b10001110101010100110;
        10'b1100000110: data <= 20'b10110111111010110000;
        10'b1100000111: data <= 20'b00101010100001111001;
        10'b1100001000: data <= 20'b00100011011001000101;
        10'b1100001001: data <= 20'b00110001010010110110;
        10'b1100001010: data <= 20'b10100011111011011010;
        10'b1100001011: data <= 20'b00100100001010101000;
        10'b1100001100: data <= 20'b00100101111001111001;
        10'b1100001101: data <= 20'b10100000110010101001;
        10'b1100001110: data <= 20'b00101100101010110010;
        10'b1100001111: data <= 20'b00101000001010101010;
        10'b1100010000: data <= 20'b10110100101011010101;
        10'b1100010001: data <= 20'b00101000001010101000;
        10'b1100010010: data <= 20'b00100111001010101010;
        10'b1100010011: data <= 20'b10101011110010101100;
        10'b1100010100: data <= 20'b00101110100010111011;
        10'b1100010101: data <= 20'b00110000001010111001;
        10'b1100010110: data <= 20'b00100100001010000101;
        10'b1100010111: data <= 20'b10101111110011000000;
        10'b1100011000: data <= 20'b00100011101010100100;
        10'b1100011001: data <= 20'b00110111011011001011;
        10'b1100011010: data <= 20'b00101101000010010001;
        10'b1100011011: data <= 20'b10101000000001100110;
        10'b1100011100: data <= 20'b00101100100010100011;
        10'b1100011101: data <= 20'b10101001001010111110;
        10'b1100011110: data <= 20'b00101000111001111100;
        10'b1100011111: data <= 20'b00101101011010001000;
        10'b1100100000: data <= 20'b10101001110010001010;
        10'b1100100001: data <= 20'b00100100010010000110;
        10'b1100100010: data <= 20'b10100010000010000010;
        10'b1100100011: data <= 20'b10100100000010100110;
        10'b1100100100: data <= 20'b00011101111010000110;
        10'b1100100101: data <= 20'b00011101010010100010;
        10'b1100100110: data <= 20'b10101100101010111010;
        10'b1100100111: data <= 20'b10101110011000101101;
        10'b1100101000: data <= 20'b00101001111010101011;
        10'b1100101001: data <= 20'b00101100010010001111;
        10'b1100101010: data <= 20'b10101000001010101100;
        10'b1100101011: data <= 20'b10101101011010110011;
        10'b1100101100: data <= 20'b10011100010010010001;
        10'b1100101101: data <= 20'b00110000000011000010;
        10'b1100101110: data <= 20'b10101110000010110001;
        10'b1100101111: data <= 20'b00101101111010110100;
        10'b1100110000: data <= 20'b00101000001010000011;
        10'b1100110001: data <= 20'b00110001111010111101;
        10'b1100110010: data <= 20'b00101010110010011101;
        10'b1100110011: data <= 20'b10101000001010101001;
        10'b1100110100: data <= 20'b10011011000010111100;
        10'b1100110101: data <= 20'b10101001011010110110;
        10'b1100110110: data <= 20'b10110001101010100100;
        10'b1100110111: data <= 20'b10100000101010011001;
        10'b1100111000: data <= 20'b10101100100010110100;
        10'b1100111001: data <= 20'b00100101010010000100;
        10'b1100111010: data <= 20'b00101011110001101001;
        10'b1100111011: data <= 20'b10101000000001110101;
        10'b1100111100: data <= 20'b00100001010010100000;
        10'b1100111101: data <= 20'b00100010110010010011;
        10'b1100111110: data <= 20'b10101000110011001010;
        10'b1100111111: data <= 20'b10101100001001110001;
        10'b1101000000: data <= 20'b00110000011010101011;
        10'b1101000001: data <= 20'b10101100111010101101;
        10'b1101000010: data <= 20'b00101010010001111111;
        10'b1101000011: data <= 20'b00100110110010100011;
        10'b1101000100: data <= 20'b00011010110010110000;
        10'b1101000101: data <= 20'b00101100101011110100;
        10'b1101000110: data <= 20'b10100001111010111101;
        10'b1101000111: data <= 20'b00100101001010100100;
        10'b1101001000: data <= 20'b10101010110010111110;
        10'b1101001001: data <= 20'b00101101101010111111;
        10'b1101001010: data <= 20'b10101001010001110010;
        10'b1101001011: data <= 20'b00100000000010011000;
        10'b1101001100: data <= 20'b00101000110010100010;
        10'b1101001101: data <= 20'b10101100111010011101;
        10'b1101001110: data <= 20'b00111000010011010010;
        10'b1101001111: data <= 20'b00010000001010100100;
        10'b1101010000: data <= 20'b00100110111010000101;
        10'b1101010001: data <= 20'b00101110010010011011;
        10'b1101010010: data <= 20'b00100100100001010011;
        10'b1101010011: data <= 20'b00100101110010101011;
        10'b1101010100: data <= 20'b00101100001011001101;
        10'b1101010101: data <= 20'b10101101101001111000;
        10'b1101010110: data <= 20'b00100111111010000010;
        10'b1101010111: data <= 20'b10100010000010010000;
        10'b1101011000: data <= 20'b10011010001010100110;
        10'b1101011001: data <= 20'b00110101100011001100;
        10'b1101011010: data <= 20'b10110100010010100111;
        10'b1101011011: data <= 20'b00100100110010000100;
        10'b1101011100: data <= 20'b10100100000010110100;
        10'b1101011101: data <= 20'b00101001011001101010;
        10'b1101011110: data <= 20'b00101001100010100100;
        10'b1101011111: data <= 20'b10110011001011000001;
        10'b1101100000: data <= 20'b00100100111010100001;
        10'b1101100001: data <= 20'b00101001010001010111;
        10'b1101100010: data <= 20'b10100111110010100011;
        10'b1101100011: data <= 20'b00101010001010100000;
        10'b1101100100: data <= 20'b10101011010010010100;
        10'b1101100101: data <= 20'b00101101101010101101;
        10'b1101100110: data <= 20'b00110001111010101100;
        10'b1101100111: data <= 20'b00101100100001111100;
        10'b1101101000: data <= 20'b10101111110010111010;
        10'b1101101001: data <= 20'b10101000100001011001;
        10'b1101101010: data <= 20'b10101011101011001101;
        10'b1101101011: data <= 20'b00100100101010011111;
        10'b1101101100: data <= 20'b00011001110010010111;
        10'b1101101101: data <= 20'b00101111000010111101;
        10'b1101101110: data <= 20'b00011101111010101101;
        10'b1101101111: data <= 20'b10101100110010110110;
        10'b1101110000: data <= 20'b00101000001000110010;
        10'b1101110001: data <= 20'b00101010011010100011;
        10'b1101110010: data <= 20'b00101100010011000011;
        10'b1101110011: data <= 20'b00110000111010110110;
        10'b1101110100: data <= 20'b10100000001010110101;
        10'b1101110101: data <= 20'b10110001101011010010;
        10'b1101110110: data <= 20'b00101000111010010101;
        10'b1101110111: data <= 20'b10101101100010111000;
        10'b1101111000: data <= 20'b10100000001010010101;
        10'b1101111001: data <= 20'b10100100011010110011;
        10'b1101111010: data <= 20'b00101100000011000001;
        10'b1101111011: data <= 20'b00011101001010010001;
        10'b1101111100: data <= 20'b00101000001010110111;
        10'b1101111101: data <= 20'b00011110100010100001;
        10'b1101111110: data <= 20'b00010010110010010100;
        10'b1101111111: data <= 20'b00100001010010100011;
        10'b1110000000: data <= 20'b10110011001010010111;
        10'b1110000001: data <= 20'b10101001100010011000;
        10'b1110000010: data <= 20'b10100000011010011110;
        10'b1110000011: data <= 20'b00110100000011010111;
        10'b1110000100: data <= 20'b10001000011011001010;
        10'b1110000101: data <= 20'b00100001101010100000;
        10'b1110000110: data <= 20'b10101001010001110111;
        10'b1110000111: data <= 20'b00101011000010101110;
        10'b1110001000: data <= 20'b10110010000010100101;
        10'b1110001001: data <= 20'b10110000110010010001;
        10'b1110001010: data <= 20'b00011001100010010001;
        10'b1110001011: data <= 20'b10011100000010111101;
        10'b1110001100: data <= 20'b00101100011010100111;
        10'b1110001101: data <= 20'b00101100111010110110;
        10'b1110001110: data <= 20'b10101000111010001011;
        10'b1110001111: data <= 20'b00011110110010110100;
        10'b1110010000: data <= 20'b10101100010010101100;
        10'b1110010001: data <= 20'b10100110010010110010;
        10'b1110010010: data <= 20'b10100101111010000100;
        10'b1110010011: data <= 20'b00001110101010010001;
        10'b1110010100: data <= 20'b00101000100010111011;
        10'b1110010101: data <= 20'b00011100111010101110;
        10'b1110010110: data <= 20'b00110101110011000110;
        10'b1110010111: data <= 20'b10101100111010111000;
        10'b1110011000: data <= 20'b10100101101010100011;
        10'b1110011001: data <= 20'b00100000110001010000;
        10'b1110011010: data <= 20'b10100100101001111000;
        10'b1110011011: data <= 20'b10100010000010100001;
        10'b1110011100: data <= 20'b00110001010010100010;
        10'b1110011101: data <= 20'b00101101101010100110;
        10'b1110011110: data <= 20'b10100101001010100101;
        10'b1110011111: data <= 20'b10111000001011000001;
        10'b1110100000: data <= 20'b00100000100010110111;
        10'b1110100001: data <= 20'b10011111011010010010;
        10'b1110100010: data <= 20'b00101000110010100011;
        10'b1110100011: data <= 20'b00011101010010110010;
        10'b1110100100: data <= 20'b00101101010010100111;
        10'b1110100101: data <= 20'b10100011011001110000;
        10'b1110100110: data <= 20'b00100110110010110000;
        10'b1110100111: data <= 20'b10100110101010110001;
        10'b1110101000: data <= 20'b00101100000010101011;
        10'b1110101001: data <= 20'b00100100001001101001;
        10'b1110101010: data <= 20'b10101010101010110000;
        10'b1110101011: data <= 20'b00101000110001011000;
        10'b1110101100: data <= 20'b10101101100011000011;
        10'b1110101101: data <= 20'b00011000111001111111;
        10'b1110101110: data <= 20'b00101010010010110000;
        10'b1110101111: data <= 20'b10101100101011100001;
        10'b1110110000: data <= 20'b00101011011011000011;
        10'b1110110001: data <= 20'b00101010101010111001;
        10'b1110110010: data <= 20'b00100011111010100100;
        10'b1110110011: data <= 20'b00101011001010000111;
        10'b1110110100: data <= 20'b00101010100010011000;
        10'b1110110101: data <= 20'b10101011100001100101;
        10'b1110110110: data <= 20'b00101101011010101010;
        10'b1110110111: data <= 20'b10110011010010101011;
        10'b1110111000: data <= 20'b00101011101010101111;
        10'b1110111001: data <= 20'b10011110110010011100;
        10'b1110111010: data <= 20'b10101001000010100000;
        10'b1110111011: data <= 20'b10100101010010100110;
        10'b1110111100: data <= 20'b10101100111010011000;
        10'b1110111101: data <= 20'b10101011101010110010;
        10'b1110111110: data <= 20'b00011001100010000001;
        10'b1110111111: data <= 20'b10101010111010110010;
        10'b1111000000: data <= 20'b00101111010010101110;
        10'b1111000001: data <= 20'b00101001001010110110;
        10'b1111000010: data <= 20'b00110000011010010111;
        10'b1111000011: data <= 20'b10101110100001111110;
        10'b1111000100: data <= 20'b00100100111010100001;
        10'b1111000101: data <= 20'b00110000110011000100;
        10'b1111000110: data <= 20'b00100100111010100100;
        10'b1111000111: data <= 20'b10101011000011100100;
        10'b1111001000: data <= 20'b10101010010010001101;
        10'b1111001001: data <= 20'b10100010100010100011;
        10'b1111001010: data <= 20'b00100010100001010110;
        10'b1111001011: data <= 20'b00100010011010000000;
        10'b1111001100: data <= 20'b10101100010011000001;
        10'b1111001101: data <= 20'b00110010011011010000;
        10'b1111001110: data <= 20'b00101100001010100001;
        10'b1111001111: data <= 20'b00001001111010001111;
        10'b1111010000: data <= 20'b10101110100011000110;
        10'b1111010001: data <= 20'b10100100010010010001;
        10'b1111010010: data <= 20'b10010000011010101000;
        10'b1111010011: data <= 20'b00101101100011000100;
        10'b1111010100: data <= 20'b10111010100011100001;
        10'b1111010101: data <= 20'b00100100000010100111;
        10'b1111010110: data <= 20'b10011000011010110001;
        10'b1111010111: data <= 20'b00101001000011010100;
        10'b1111011000: data <= 20'b00101000101001001110;
        10'b1111011001: data <= 20'b00101001110010010010;
        10'b1111011010: data <= 20'b10110000001011010101;
        10'b1111011011: data <= 20'b10100100110010101010;
        10'b1111011100: data <= 20'b10101010000010000000;
        10'b1111011101: data <= 20'b00100110101010010100;
        10'b1111011110: data <= 20'b10101000000010100001;
        10'b1111011111: data <= 20'b00100111100010101000;
        10'b1111100000: data <= 20'b10101011110001011100;
        10'b1111100001: data <= 20'b10011010000011000101;
        10'b1111100010: data <= 20'b10100110111011000000;
        10'b1111100011: data <= 20'b00100100101001111111;
        10'b1111100100: data <= 20'b00100110111001010111;
        10'b1111100101: data <= 20'b00100010010010111101;
        10'b1111100110: data <= 20'b00101110101010111111;
        10'b1111100111: data <= 20'b10101011101010110011;
        10'b1111101000: data <= 20'b00011101101010011101;
        10'b1111101001: data <= 20'b00101101000011010011;
        10'b1111101010: data <= 20'b00100001010010010000;
        10'b1111101011: data <= 20'b10101100110010100010;
        10'b1111101100: data <= 20'b00101001001010011100;
        10'b1111101101: data <= 20'b10101001101010110001;
        10'b1111101110: data <= 20'b00100101010010010100;
        10'b1111101111: data <= 20'b00101010010010000101;
        10'b1111110000: data <= 20'b10110000001011000010;
        10'b1111110001: data <= 20'b00110011101010000111;
        10'b1111110010: data <= 20'b10100100010010010100;
        10'b1111110011: data <= 20'b00101001010010110010;
        10'b1111110100: data <= 20'b10011110111010100001;
        10'b1111110101: data <= 20'b10011100110010110111;
        10'b1111110110: data <= 20'b10011101001010000100;
        10'b1111110111: data <= 20'b10100111110010110011;
        10'b1111111000: data <= 20'b10011100111011000010;
        10'b1111111001: data <= 20'b00101001101011001011;
        10'b1111111010: data <= 20'b00100001000001111100;
        10'b1111111011: data <= 20'b10101000010010010001;
        10'b1111111100: data <= 20'b00011101100010100001;
    
    endcase
    end
    end

    assign Q = data;

    endmodule

        