
module memory_rom_58(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'habe1be4d;
    11'b00000000001: data <= 32'haf21bb87;
    11'b00000000010: data <= 32'h25583afb;
    11'b00000000011: data <= 32'hb9cd3ee4;
    11'b00000000100: data <= 32'hbec33507;
    11'b00000000101: data <= 32'hbea8be92;
    11'b00000000110: data <= 32'hbb47bea4;
    11'b00000000111: data <= 32'hb83c2dd9;
    11'b00000001000: data <= 32'hb7033d19;
    11'b00000001001: data <= 32'h35573b1e;
    11'b00000001010: data <= 32'h3ddc364b;
    11'b00000001011: data <= 32'h3d3a3c19;
    11'b00000001100: data <= 32'hb71d3f58;
    11'b00000001101: data <= 32'hbebd3d8f;
    11'b00000001110: data <= 32'hb95c2bcd;
    11'b00000001111: data <= 32'h3d88b9ed;
    11'b00000010000: data <= 32'h3fe9ba73;
    11'b00000010001: data <= 32'h3b03bbdd;
    11'b00000010010: data <= 32'h30ddbce0;
    11'b00000010011: data <= 32'h3a9ab84e;
    11'b00000010100: data <= 32'h3d983ab4;
    11'b00000010101: data <= 32'h36323c77;
    11'b00000010110: data <= 32'hbd54b75d;
    11'b00000010111: data <= 32'hbfb7c028;
    11'b00000011000: data <= 32'hbd09bee9;
    11'b00000011001: data <= 32'hb8c0aeac;
    11'b00000011010: data <= 32'hb5d037ec;
    11'b00000011011: data <= 32'h2ea6b521;
    11'b00000011100: data <= 32'h39cab884;
    11'b00000011101: data <= 32'h35c13b17;
    11'b00000011110: data <= 32'hbc4b40e4;
    11'b00000011111: data <= 32'hbf4f4054;
    11'b00000100000: data <= 32'hb9b13826;
    11'b00000100001: data <= 32'h3b79b875;
    11'b00000100010: data <= 32'h3c70b7a5;
    11'b00000100011: data <= 32'h31bcb3d5;
    11'b00000100100: data <= 32'h3402b4a8;
    11'b00000100101: data <= 32'h3efb2d39;
    11'b00000100110: data <= 32'h41173b35;
    11'b00000100111: data <= 32'h3c993b40;
    11'b00000101000: data <= 32'hbc1db6d6;
    11'b00000101001: data <= 32'hbeaebe94;
    11'b00000101010: data <= 32'hb98ebd59;
    11'b00000101011: data <= 32'h30b9b62c;
    11'b00000101100: data <= 32'h2d64b8cb;
    11'b00000101101: data <= 32'ha895bec1;
    11'b00000101110: data <= 32'h32c8bdfa;
    11'b00000101111: data <= 32'ha25338df;
    11'b00000110000: data <= 32'hbc3040dd;
    11'b00000110001: data <= 32'hbed13fc8;
    11'b00000110010: data <= 32'hbc4d2ddb;
    11'b00000110011: data <= 32'hb0ceba0d;
    11'b00000110100: data <= 32'hb435ae85;
    11'b00000110101: data <= 32'hb9fa3865;
    11'b00000110110: data <= 32'h2f993675;
    11'b00000110111: data <= 32'h402c3563;
    11'b00000111000: data <= 32'h41933b53;
    11'b00000111001: data <= 32'h3c723cdd;
    11'b00000111010: data <= 32'hbbe6378f;
    11'b00000111011: data <= 32'hbc8bb78c;
    11'b00000111100: data <= 32'h3459b8aa;
    11'b00000111101: data <= 32'h3c20b7ab;
    11'b00000111110: data <= 32'h3759bd3c;
    11'b00000111111: data <= 32'hab8bc0ca;
    11'b00001000000: data <= 32'h34f4bf5d;
    11'b00001000001: data <= 32'h3888364e;
    11'b00001000010: data <= 32'hb27a3f8f;
    11'b00001000011: data <= 32'hbce73bfe;
    11'b00001000100: data <= 32'hbdaeba73;
    11'b00001000101: data <= 32'hbca5bc68;
    11'b00001000110: data <= 32'hbd4b2e86;
    11'b00001000111: data <= 32'hbd803a59;
    11'b00001001000: data <= 32'hb1293373;
    11'b00001001001: data <= 32'h3eceb09f;
    11'b00001001010: data <= 32'h402539a4;
    11'b00001001011: data <= 32'h363c3f08;
    11'b00001001100: data <= 32'hbcbf3ea8;
    11'b00001001101: data <= 32'hb9893a1e;
    11'b00001001110: data <= 32'h3b3130c0;
    11'b00001001111: data <= 32'h3d25b46e;
    11'b00001010000: data <= 32'h34d1bcda;
    11'b00001010001: data <= 32'haec1c023;
    11'b00001010010: data <= 32'h3b3fbdc8;
    11'b00001010011: data <= 32'h3f193604;
    11'b00001010100: data <= 32'h3c1c3cef;
    11'b00001010101: data <= 32'hb8982c39;
    11'b00001010110: data <= 32'hbdc2bda5;
    11'b00001010111: data <= 32'hbdc6bcb3;
    11'b00001011000: data <= 32'hbdc8303b;
    11'b00001011001: data <= 32'hbd6d3562;
    11'b00001011010: data <= 32'hb66fba6c;
    11'b00001011011: data <= 32'h3b61bcdd;
    11'b00001011100: data <= 32'h3bfe3411;
    11'b00001011101: data <= 32'hb653402c;
    11'b00001011110: data <= 32'hbd6c40b5;
    11'b00001011111: data <= 32'hb8583d3a;
    11'b00001100000: data <= 32'h3a013716;
    11'b00001100001: data <= 32'h38c62e71;
    11'b00001100010: data <= 32'hb7fab718;
    11'b00001100011: data <= 32'hb535bc2e;
    11'b00001100100: data <= 32'h3e16b986;
    11'b00001100101: data <= 32'h41a637b0;
    11'b00001100110: data <= 32'h3f983af4;
    11'b00001100111: data <= 32'haec6b1b9;
    11'b00001101000: data <= 32'hbc59bca4;
    11'b00001101001: data <= 32'hbac2b99a;
    11'b00001101010: data <= 32'hb9263137;
    11'b00001101011: data <= 32'hba6eb70f;
    11'b00001101100: data <= 32'hb7ebc020;
    11'b00001101101: data <= 32'h349dc08c;
    11'b00001101110: data <= 32'h35f9b395;
    11'b00001101111: data <= 32'hb8763fba;
    11'b00001110000: data <= 32'hbcb24031;
    11'b00001110001: data <= 32'hb8e33ad7;
    11'b00001110010: data <= 32'ha24e31b5;
    11'b00001110011: data <= 32'hb9473700;
    11'b00001110100: data <= 32'hbe453727;
    11'b00001110101: data <= 32'hb9b3afe7;
    11'b00001110110: data <= 32'h3eb9b3bc;
    11'b00001110111: data <= 32'h42093774;
    11'b00001111000: data <= 32'h3f7c3b41;
    11'b00001111001: data <= 32'had383665;
    11'b00001111010: data <= 32'hb891af51;
    11'b00001111011: data <= 32'h32613277;
    11'b00001111100: data <= 32'h370635b8;
    11'b00001111101: data <= 32'hb398bb7a;
    11'b00001111110: data <= 32'hb825c170;
    11'b00001111111: data <= 32'h30a8c156;
    11'b00010000000: data <= 32'h3917b7d2;
    11'b00010000001: data <= 32'h30a33d84;
    11'b00010000010: data <= 32'hb86b3c54;
    11'b00010000011: data <= 32'hb92db2ca;
    11'b00010000100: data <= 32'hba3ab58d;
    11'b00010000101: data <= 32'hbeab38f5;
    11'b00010000110: data <= 32'hc0903b32;
    11'b00010000111: data <= 32'hbc5721a1;
    11'b00010001000: data <= 32'h3d00b883;
    11'b00010001001: data <= 32'h407d3029;
    11'b00010001010: data <= 32'h3c0d3c89;
    11'b00010001011: data <= 32'hb70c3d4a;
    11'b00010001100: data <= 32'hb11e3c42;
    11'b00010001101: data <= 32'h3c063c38;
    11'b00010001110: data <= 32'h3be539ab;
    11'b00010001111: data <= 32'hb30bba0e;
    11'b00010010000: data <= 32'hb951c0af;
    11'b00010010001: data <= 32'h36ecc059;
    11'b00010010010: data <= 32'h3e3eb60c;
    11'b00010010011: data <= 32'h3d3d3a10;
    11'b00010010100: data <= 32'h33e8a05f;
    11'b00010010101: data <= 32'hb775bc62;
    11'b00010010110: data <= 32'hbb89b8e0;
    11'b00010010111: data <= 32'hbefe39c5;
    11'b00010011000: data <= 32'hc06b39e5;
    11'b00010011001: data <= 32'hbcf4b9d8;
    11'b00010011010: data <= 32'h37fbbe3a;
    11'b00010011011: data <= 32'h3c22b7ba;
    11'b00010011100: data <= 32'ha8903ce0;
    11'b00010011101: data <= 32'hba783f71;
    11'b00010011110: data <= 32'h280d3e4c;
    11'b00010011111: data <= 32'h3c893d62;
    11'b00010100000: data <= 32'h38c63c33;
    11'b00010100001: data <= 32'hbb6618f4;
    11'b00010100010: data <= 32'hbc31bccc;
    11'b00010100011: data <= 32'h3a36bcb5;
    11'b00010100100: data <= 32'h40daac7b;
    11'b00010100101: data <= 32'h404e35fe;
    11'b00010100110: data <= 32'h3a16b815;
    11'b00010100111: data <= 32'hade4bc9a;
    11'b00010101000: data <= 32'hb549b401;
    11'b00010101001: data <= 32'hbac53b42;
    11'b00010101010: data <= 32'hbdc833e9;
    11'b00010101011: data <= 32'hbc8abf23;
    11'b00010101100: data <= 32'hb04bc12f;
    11'b00010101101: data <= 32'h316abc40;
    11'b00010101110: data <= 32'hb8133be4;
    11'b00010101111: data <= 32'hba233e3d;
    11'b00010110000: data <= 32'h2e8e3c29;
    11'b00010110001: data <= 32'h39563b48;
    11'b00010110010: data <= 32'hb6f23cd9;
    11'b00010110011: data <= 32'hbfe13b0b;
    11'b00010110100: data <= 32'hbe3dab95;
    11'b00010110101: data <= 32'h3a72b6a1;
    11'b00010110110: data <= 32'h411b2d3a;
    11'b00010110111: data <= 32'h402034c2;
    11'b00010111000: data <= 32'h394bb358;
    11'b00010111001: data <= 32'h348cb596;
    11'b00010111010: data <= 32'h399a38fc;
    11'b00010111011: data <= 32'h36f53d02;
    11'b00010111100: data <= 32'hb88eac8e;
    11'b00010111101: data <= 32'hbbc1c0b1;
    11'b00010111110: data <= 32'hb5d5c1e3;
    11'b00010111111: data <= 32'h3069bcf8;
    11'b00011000000: data <= 32'hac95383b;
    11'b00011000001: data <= 32'hb20e386a;
    11'b00011000010: data <= 32'h3372b28e;
    11'b00011000011: data <= 32'h2f352dba;
    11'b00011000100: data <= 32'hbd4d3cc4;
    11'b00011000101: data <= 32'hc1533d93;
    11'b00011000110: data <= 32'hbfa835cd;
    11'b00011000111: data <= 32'h36beb737;
    11'b00011001000: data <= 32'h3f15b1f2;
    11'b00011001001: data <= 32'h3c3035ad;
    11'b00011001010: data <= 32'h27b9373e;
    11'b00011001011: data <= 32'h37dd398a;
    11'b00011001100: data <= 32'h3e323de2;
    11'b00011001101: data <= 32'h3d0a3e8d;
    11'b00011001110: data <= 32'hb3ef2f0b;
    11'b00011001111: data <= 32'hbc11bfca;
    11'b00011010000: data <= 32'hb39ac0a1;
    11'b00011010001: data <= 32'h3a66bb22;
    11'b00011010010: data <= 32'h3b752e6e;
    11'b00011010011: data <= 32'h38edb88b;
    11'b00011010100: data <= 32'h37eebd6d;
    11'b00011010101: data <= 32'h19f2b7dd;
    11'b00011010110: data <= 32'hbd7d3ca7;
    11'b00011010111: data <= 32'hc0f93d7f;
    11'b00011011000: data <= 32'hbf7aaea3;
    11'b00011011001: data <= 32'hb113bd07;
    11'b00011011010: data <= 32'h3848ba6e;
    11'b00011011011: data <= 32'hb4263522;
    11'b00011011100: data <= 32'hb9533b1e;
    11'b00011011101: data <= 32'h38373c9d;
    11'b00011011110: data <= 32'h3f343ec4;
    11'b00011011111: data <= 32'h3c9e3f55;
    11'b00011100000: data <= 32'hb9ea39d4;
    11'b00011100001: data <= 32'hbd93ba47;
    11'b00011100010: data <= 32'ha8b3bc4c;
    11'b00011100011: data <= 32'h3e19b412;
    11'b00011100100: data <= 32'h3ed9aecf;
    11'b00011100101: data <= 32'h3c5dbcb5;
    11'b00011100110: data <= 32'h3a41bed0;
    11'b00011100111: data <= 32'h381ab5fc;
    11'b00011101000: data <= 32'hb7333d4b;
    11'b00011101001: data <= 32'hbe003c28;
    11'b00011101010: data <= 32'hbdc9bbdd;
    11'b00011101011: data <= 32'hb8d1c06c;
    11'b00011101100: data <= 32'hb6bbbd7d;
    11'b00011101101: data <= 32'hbc222fa2;
    11'b00011101110: data <= 32'hbb2a392d;
    11'b00011101111: data <= 32'h385e38cb;
    11'b00011110000: data <= 32'h3df73c42;
    11'b00011110001: data <= 32'h35353ecc;
    11'b00011110010: data <= 32'hbebf3da9;
    11'b00011110011: data <= 32'hbfa736f5;
    11'b00011110100: data <= 32'ha7039e6b;
    11'b00011110101: data <= 32'h3ea83259;
    11'b00011110110: data <= 32'h3e64ae85;
    11'b00011110111: data <= 32'h3ab0bc35;
    11'b00011111000: data <= 32'h3b34bc84;
    11'b00011111001: data <= 32'h3d73360e;
    11'b00011111010: data <= 32'h3b323ebe;
    11'b00011111011: data <= 32'hb51e3a43;
    11'b00011111100: data <= 32'hbba3be13;
    11'b00011111101: data <= 32'hb9c3c112;
    11'b00011111110: data <= 32'hb8d1bdbc;
    11'b00011111111: data <= 32'hbac7b017;
    11'b00100000000: data <= 32'hb77bb274;
    11'b00100000001: data <= 32'h398eb9a8;
    11'b00100000010: data <= 32'h3c20aaa1;
    11'b00100000011: data <= 32'hb8083d5c;
    11'b00100000100: data <= 32'hc0b33f28;
    11'b00100000101: data <= 32'hc0603bfc;
    11'b00100000110: data <= 32'hb40a337d;
    11'b00100000111: data <= 32'h3c0e2f7c;
    11'b00100001000: data <= 32'h3838aa9a;
    11'b00100001001: data <= 32'hacb0b7d6;
    11'b00100001010: data <= 32'h3a26b1d8;
    11'b00100001011: data <= 32'h401b3cc7;
    11'b00100001100: data <= 32'h3f6e400f;
    11'b00100001101: data <= 32'h34cf3adc;
    11'b00100001110: data <= 32'hba36bce3;
    11'b00100001111: data <= 32'hb8a1bf72;
    11'b00100010000: data <= 32'hacedbaa5;
    11'b00100010001: data <= 32'h26c0b364;
    11'b00100010010: data <= 32'h34b6bca1;
    11'b00100010011: data <= 32'h3b94bff0;
    11'b00100010100: data <= 32'h3aefbb96;
    11'b00100010101: data <= 32'hb8fc3c31;
    11'b00100010110: data <= 32'hc0463ee9;
    11'b00100010111: data <= 32'hbfb2396c;
    11'b00100011000: data <= 32'hb842b685;
    11'b00100011001: data <= 32'hab8bb701;
    11'b00100011010: data <= 32'hbb30ae38;
    11'b00100011011: data <= 32'hbc63a9b2;
    11'b00100011100: data <= 32'h38113522;
    11'b00100011101: data <= 32'h40783d90;
    11'b00100011110: data <= 32'h3f9c4018;
    11'b00100011111: data <= 32'h20413cd7;
    11'b00100100000: data <= 32'hbc3eb2d5;
    11'b00100100001: data <= 32'hb65db80e;
    11'b00100100010: data <= 32'h38ee3070;
    11'b00100100011: data <= 32'h3a8aaf93;
    11'b00100100100: data <= 32'h3a0fbeb2;
    11'b00100100101: data <= 32'h3c69c0f9;
    11'b00100100110: data <= 32'h3c9dbc42;
    11'b00100100111: data <= 32'h31033c51;
    11'b00100101000: data <= 32'hbc313da3;
    11'b00100101001: data <= 32'hbcb3b06b;
    11'b00100101010: data <= 32'hb924bd5d;
    11'b00100101011: data <= 32'hbb3fbbfd;
    11'b00100101100: data <= 32'hbf55b2cc;
    11'b00100101101: data <= 32'hbe61af37;
    11'b00100101110: data <= 32'h35c1aedd;
    11'b00100101111: data <= 32'h3fba396d;
    11'b00100110000: data <= 32'h3ca43e6e;
    11'b00100110001: data <= 32'hbb143e3f;
    11'b00100110010: data <= 32'hbe473b13;
    11'b00100110011: data <= 32'hb56d39d0;
    11'b00100110100: data <= 32'h3b0f3b26;
    11'b00100110101: data <= 32'h3a7e2e19;
    11'b00100110110: data <= 32'h3701be27;
    11'b00100110111: data <= 32'h3b93c00a;
    11'b00100111000: data <= 32'h3ebab668;
    11'b00100111001: data <= 32'h3d823daf;
    11'b00100111010: data <= 32'h34c43c85;
    11'b00100111011: data <= 32'hb5a9ba0f;
    11'b00100111100: data <= 32'hb816bf04;
    11'b00100111101: data <= 32'hbc3cbc11;
    11'b00100111110: data <= 32'hbf1db337;
    11'b00100111111: data <= 32'hbd2eb950;
    11'b00101000000: data <= 32'h3777bd21;
    11'b00101000001: data <= 32'h3ddfb8ca;
    11'b00101000010: data <= 32'h348f3b36;
    11'b00101000011: data <= 32'hbe783e9c;
    11'b00101000100: data <= 32'hbf493d9a;
    11'b00101000101: data <= 32'hb5fb3c79;
    11'b00101000110: data <= 32'h37f43be3;
    11'b00101000111: data <= 32'hb03632f3;
    11'b00101001000: data <= 32'hb8f9bbda;
    11'b00101001001: data <= 32'h3772bc3f;
    11'b00101001010: data <= 32'h4022376c;
    11'b00101001011: data <= 32'h408b3f08;
    11'b00101001100: data <= 32'h3c5a3c3b;
    11'b00101001101: data <= 32'h29e1b987;
    11'b00101001110: data <= 32'hb425bccf;
    11'b00101001111: data <= 32'hb853b47c;
    11'b00101010000: data <= 32'hbb68218c;
    11'b00101010001: data <= 32'hb816bd37;
    11'b00101010010: data <= 32'h39c9c0f8;
    11'b00101010011: data <= 32'h3cc8beb8;
    11'b00101010100: data <= 32'ha75e357d;
    11'b00101010101: data <= 32'hbe193dbf;
    11'b00101010110: data <= 32'hbdc93c54;
    11'b00101010111: data <= 32'hb55d3841;
    11'b00101011000: data <= 32'hb433371d;
    11'b00101011001: data <= 32'hbde7315d;
    11'b00101011010: data <= 32'hbf5bb76e;
    11'b00101011011: data <= 32'hae4fb662;
    11'b00101011100: data <= 32'h401b3a38;
    11'b00101011101: data <= 32'h409e3ec6;
    11'b00101011110: data <= 32'h3b103c7d;
    11'b00101011111: data <= 32'hb1d1232e;
    11'b00101100000: data <= 32'hac6a2c34;
    11'b00101100001: data <= 32'h32523b1c;
    11'b00101100010: data <= 32'ha1893749;
    11'b00101100011: data <= 32'h2c18be5d;
    11'b00101100100: data <= 32'h3a9dc1f1;
    11'b00101100101: data <= 32'h3ceebfa8;
    11'b00101100110: data <= 32'h3767344f;
    11'b00101100111: data <= 32'hb83b3c56;
    11'b00101101000: data <= 32'hb802339f;
    11'b00101101001: data <= 32'hae2cb7d8;
    11'b00101101010: data <= 32'hbad3b2eb;
    11'b00101101011: data <= 32'hc0c72ceb;
    11'b00101101100: data <= 32'hc0f9b531;
    11'b00101101101: data <= 32'hb674b87a;
    11'b00101101110: data <= 32'h3ebb3159;
    11'b00101101111: data <= 32'h3e323c49;
    11'b00101110000: data <= 32'hac193c7b;
    11'b00101110001: data <= 32'hba293ab2;
    11'b00101110010: data <= 32'h9c3f3d18;
    11'b00101110011: data <= 32'h390d3f4c;
    11'b00101110100: data <= 32'h33423b02;
    11'b00101110101: data <= 32'hb09bbd6b;
    11'b00101110110: data <= 32'h381dc0fc;
    11'b00101110111: data <= 32'h3daabcee;
    11'b00101111000: data <= 32'h3d97394c;
    11'b00101111001: data <= 32'h3a4b3a74;
    11'b00101111010: data <= 32'h3838b81e;
    11'b00101111011: data <= 32'h34a7bc7c;
    11'b00101111100: data <= 32'hbaf6b5ac;
    11'b00101111101: data <= 32'hc0a73210;
    11'b00101111110: data <= 32'hc06bb86e;
    11'b00101111111: data <= 32'hb484bdc9;
    11'b00110000000: data <= 32'h3cdebc48;
    11'b00110000001: data <= 32'h3888308e;
    11'b00110000010: data <= 32'hbbe93b50;
    11'b00110000011: data <= 32'hbc963cbb;
    11'b00110000100: data <= 32'h2af83eaa;
    11'b00110000101: data <= 32'h38503fef;
    11'b00110000110: data <= 32'hb6ea3c1e;
    11'b00110000111: data <= 32'hbc9cba46;
    11'b00110001000: data <= 32'hb22bbdcd;
    11'b00110001001: data <= 32'h3de6b275;
    11'b00110001010: data <= 32'h402f3c80;
    11'b00110001011: data <= 32'h3e54395c;
    11'b00110001100: data <= 32'h3c28b9ad;
    11'b00110001101: data <= 32'h3905bac5;
    11'b00110001110: data <= 32'hb5163517;
    11'b00110001111: data <= 32'hbda63923;
    11'b00110010000: data <= 32'hbd2abad5;
    11'b00110010001: data <= 32'h2e13c0da;
    11'b00110010010: data <= 32'h3b40c052;
    11'b00110010011: data <= 32'h258eb892;
    11'b00110010100: data <= 32'hbca83875;
    11'b00110010101: data <= 32'hbad23a6e;
    11'b00110010110: data <= 32'h34aa3c25;
    11'b00110010111: data <= 32'h2fb53d62;
    11'b00110011000: data <= 32'hbe283b03;
    11'b00110011001: data <= 32'hc0c2b3dd;
    11'b00110011010: data <= 32'hbb95b8af;
    11'b00110011011: data <= 32'h3d1235f3;
    11'b00110011100: data <= 32'h40143ca4;
    11'b00110011101: data <= 32'h3d68387e;
    11'b00110011110: data <= 32'h3a18b56a;
    11'b00110011111: data <= 32'h39f63199;
    11'b00110100000: data <= 32'h36ed3dfa;
    11'b00110100001: data <= 32'hb52f3d37;
    11'b00110100010: data <= 32'hb77bbb36;
    11'b00110100011: data <= 32'h3514c196;
    11'b00110100100: data <= 32'h3a67c0c6;
    11'b00110100101: data <= 32'h322ab92a;
    11'b00110100110: data <= 32'hb6cb3381;
    11'b00110100111: data <= 32'h2df0ab27;
    11'b00110101000: data <= 32'h3a1bb03d;
    11'b00110101001: data <= 32'hb2443748;
    11'b00110101010: data <= 32'hc09f3938;
    11'b00110101011: data <= 32'hc2131c89;
    11'b00110101100: data <= 32'hbd38b718;
    11'b00110101101: data <= 32'h3b0626aa;
    11'b00110101110: data <= 32'h3d00386f;
    11'b00110101111: data <= 32'h34873528;
    11'b00110110000: data <= 32'ha79531e9;
    11'b00110110001: data <= 32'h39633ce5;
    11'b00110110010: data <= 32'h3b9640e9;
    11'b00110110011: data <= 32'h323a3f4f;
    11'b00110110100: data <= 32'hb673b8c1;
    11'b00110110101: data <= 32'h29bcc08b;
    11'b00110110110: data <= 32'h3a0abe6d;
    11'b00110110111: data <= 32'h3a7cad5e;
    11'b00110111000: data <= 32'h39b62d5e;
    11'b00110111001: data <= 32'h3ca4baf5;
    11'b00110111010: data <= 32'h3d35bc17;
    11'b00110111011: data <= 32'hadd72911;
    11'b00110111100: data <= 32'hc0613995;
    11'b00110111101: data <= 32'hc160a416;
    11'b00110111110: data <= 32'hbc39bc07;
    11'b00110111111: data <= 32'h3827bc11;
    11'b00111000000: data <= 32'h3306b6b5;
    11'b00111000001: data <= 32'hbb09acd1;
    11'b00111000010: data <= 32'hb97735ca;
    11'b00111000011: data <= 32'h391c3e2a;
    11'b00111000100: data <= 32'h3c274126;
    11'b00111000101: data <= 32'hb08b3f9d;
    11'b00111000110: data <= 32'hbcccae6c;
    11'b00111000111: data <= 32'hb99cbcbe;
    11'b00111001000: data <= 32'h38c2b5c1;
    11'b00111001001: data <= 32'h3d2d3934;
    11'b00111001010: data <= 32'h3dae2bc0;
    11'b00111001011: data <= 32'h3ea9bce1;
    11'b00111001100: data <= 32'h3e79bc41;
    11'b00111001101: data <= 32'h36c337b6;
    11'b00111001110: data <= 32'hbcee3cb3;
    11'b00111001111: data <= 32'hbe4ead60;
    11'b00111010000: data <= 32'hb6bbbef8;
    11'b00111010001: data <= 32'h3557c001;
    11'b00111010010: data <= 32'hb756bc9e;
    11'b00111010011: data <= 32'hbd76b78c;
    11'b00111010100: data <= 32'hb919a653;
    11'b00111010101: data <= 32'h3b083af0;
    11'b00111010110: data <= 32'h3ad33f19;
    11'b00111010111: data <= 32'hbbdb3e11;
    11'b00111011000: data <= 32'hc09d34ed;
    11'b00111011001: data <= 32'hbe01b29e;
    11'b00111011010: data <= 32'h34af3824;
    11'b00111011011: data <= 32'h3cbf3b9e;
    11'b00111011100: data <= 32'h3c91a661;
    11'b00111011101: data <= 32'h3d0bbc4d;
    11'b00111011110: data <= 32'h3e28b538;
    11'b00111011111: data <= 32'h3c343e16;
    11'b00111100000: data <= 32'ha9ea3f94;
    11'b00111100001: data <= 32'hb75620af;
    11'b00111100010: data <= 32'h2d71c005;
    11'b00111100011: data <= 32'h3479c059;
    11'b00111100100: data <= 32'hb801bc91;
    11'b00111100101: data <= 32'hbb61b92c;
    11'b00111100110: data <= 32'h30e5ba41;
    11'b00111100111: data <= 32'h3da8b62e;
    11'b00111101000: data <= 32'h39b338d5;
    11'b00111101001: data <= 32'hbe763c00;
    11'b00111101010: data <= 32'hc1cf37a9;
    11'b00111101011: data <= 32'hbf3e303e;
    11'b00111101100: data <= 32'h9ce837b4;
    11'b00111101101: data <= 32'h37883834;
    11'b00111101110: data <= 32'h99bdb52b;
    11'b00111101111: data <= 32'h32c6ba06;
    11'b00111110000: data <= 32'h3cb5386a;
    11'b00111110001: data <= 32'h3ddd40d8;
    11'b00111110010: data <= 32'h393740d2;
    11'b00111110011: data <= 32'hacbb3481;
    11'b00111110100: data <= 32'h2569be1a;
    11'b00111110101: data <= 32'h321fbd4d;
    11'b00111110110: data <= 32'hae63b59f;
    11'b00111110111: data <= 32'h244db82e;
    11'b00111111000: data <= 32'h3c9dbdf0;
    11'b00111111001: data <= 32'h3feabdc2;
    11'b00111111010: data <= 32'h3ab3b06b;
    11'b00111111011: data <= 32'hbdfc3a72;
    11'b00111111100: data <= 32'hc0fd379f;
    11'b00111111101: data <= 32'hbd79b2a2;
    11'b00111111110: data <= 32'haf81b559;
    11'b00111111111: data <= 32'hb734b5e8;
    11'b01000000000: data <= 32'hbd43ba32;
    11'b01000000001: data <= 32'hba29b92e;
    11'b01000000010: data <= 32'h3b033ab3;
    11'b01000000011: data <= 32'h3e2e40f9;
    11'b01000000100: data <= 32'h384d40ab;
    11'b01000000101: data <= 32'hb8ee3889;
    11'b01000000110: data <= 32'hb902b852;
    11'b01000000111: data <= 32'ha8f22bd8;
    11'b01000001000: data <= 32'h344839a9;
    11'b01000001001: data <= 32'h3943b42e;
    11'b01000001010: data <= 32'h3e77bf31;
    11'b01000001011: data <= 32'h4062beca;
    11'b01000001100: data <= 32'h3cc226e1;
    11'b01000001101: data <= 32'hb8fc3ca0;
    11'b01000001110: data <= 32'hbd0337b0;
    11'b01000001111: data <= 32'hb6b2ba55;
    11'b01000010000: data <= 32'ha02fbce3;
    11'b01000010001: data <= 32'hbc48bc48;
    11'b01000010010: data <= 32'hc006bc76;
    11'b01000010011: data <= 32'hbc18bb67;
    11'b01000010100: data <= 32'h3ba9334d;
    11'b01000010101: data <= 32'h3db03e4b;
    11'b01000010110: data <= 32'hb00d3e9e;
    11'b01000010111: data <= 32'hbe613975;
    11'b01000011000: data <= 32'hbd9235e0;
    11'b01000011001: data <= 32'hb5483c95;
    11'b01000011010: data <= 32'h32d33d53;
    11'b01000011011: data <= 32'h36beb0ee;
    11'b01000011100: data <= 32'h3c78becc;
    11'b01000011101: data <= 32'h3f69bc9b;
    11'b01000011110: data <= 32'h3e283b45;
    11'b01000011111: data <= 32'h37bd3f5a;
    11'b01000100000: data <= 32'h2c5238c8;
    11'b01000100001: data <= 32'h36d8bc3f;
    11'b01000100010: data <= 32'h313fbda5;
    11'b01000100011: data <= 32'hbc8fbbe0;
    11'b01000100100: data <= 32'hbf19bc4c;
    11'b01000100101: data <= 32'hb6c2bdba;
    11'b01000100110: data <= 32'h3dc4bb8e;
    11'b01000100111: data <= 32'h3d5132b0;
    11'b01000101000: data <= 32'hb9be3a47;
    11'b01000101001: data <= 32'hc05f38c6;
    11'b01000101010: data <= 32'hbe9939b6;
    11'b01000101011: data <= 32'hb7603d4e;
    11'b01000101100: data <= 32'hb4a63c81;
    11'b01000101101: data <= 32'hb92fb60f;
    11'b01000101110: data <= 32'haf35bdc1;
    11'b01000101111: data <= 32'h3c8db5a4;
    11'b01000110000: data <= 32'h3eb43f1c;
    11'b01000110001: data <= 32'h3cae40a2;
    11'b01000110010: data <= 32'h396f3a06;
    11'b01000110011: data <= 32'h38fcb9f4;
    11'b01000110100: data <= 32'h31beb904;
    11'b01000110101: data <= 32'hba71a7cb;
    11'b01000110110: data <= 32'hbb92b8e6;
    11'b01000110111: data <= 32'h3830bf63;
    11'b01000111000: data <= 32'h3ff1bfe1;
    11'b01000111001: data <= 32'h3d89ba24;
    11'b01000111010: data <= 32'hb9c634b4;
    11'b01000111011: data <= 32'hbf513741;
    11'b01000111100: data <= 32'hbc4336fa;
    11'b01000111101: data <= 32'hb42e3936;
    11'b01000111110: data <= 32'hbb70350a;
    11'b01000111111: data <= 32'hbfb1ba88;
    11'b01001000000: data <= 32'hbd54bd38;
    11'b01001000001: data <= 32'h3813229b;
    11'b01001000010: data <= 32'h3e4c3f8d;
    11'b01001000011: data <= 32'h3c6d4040;
    11'b01001000100: data <= 32'h34e03a18;
    11'b01001000101: data <= 32'h2e0ea62f;
    11'b01001000110: data <= 32'ha83739bf;
    11'b01001000111: data <= 32'hb71c3d11;
    11'b01001001000: data <= 32'hb44293a4;
    11'b01001001001: data <= 32'h3c16bfc9;
    11'b01001001010: data <= 32'h4039c088;
    11'b01001001011: data <= 32'h3e03ba5c;
    11'b01001001100: data <= 32'hadc637c3;
    11'b01001001101: data <= 32'hb90c36c4;
    11'b01001001110: data <= 32'h2f7aaf7f;
    11'b01001001111: data <= 32'h32b6b384;
    11'b01001010000: data <= 32'hbd3eb690;
    11'b01001010001: data <= 32'hc14bbc6a;
    11'b01001010010: data <= 32'hbf34bd97;
    11'b01001010011: data <= 32'h3634b623;
    11'b01001010100: data <= 32'h3d903c13;
    11'b01001010101: data <= 32'h37ca3ce8;
    11'b01001010110: data <= 32'hb916381e;
    11'b01001010111: data <= 32'hb96c3907;
    11'b01001011000: data <= 32'hb4bd3f4a;
    11'b01001011001: data <= 32'hb5d04040;
    11'b01001011010: data <= 32'hb52c35a4;
    11'b01001011011: data <= 32'h3894bf04;
    11'b01001011100: data <= 32'h3e50bf14;
    11'b01001011101: data <= 32'h3e02235b;
    11'b01001011110: data <= 32'h3a0a3c96;
    11'b01001011111: data <= 32'h39a03837;
    11'b01001100000: data <= 32'h3ce0b7a2;
    11'b01001100001: data <= 32'h395bb88d;
    11'b01001100010: data <= 32'hbd03b608;
    11'b01001100011: data <= 32'hc0ebbb33;
    11'b01001100100: data <= 32'hbd39be52;
    11'b01001100101: data <= 32'h3a90bd2f;
    11'b01001100110: data <= 32'h3d27b5a7;
    11'b01001100111: data <= 32'hb10d2da9;
    11'b01001101000: data <= 32'hbd592eba;
    11'b01001101001: data <= 32'hbbe93a87;
    11'b01001101010: data <= 32'hb4cc401d;
    11'b01001101011: data <= 32'hb8a54020;
    11'b01001101100: data <= 32'hbc9332f2;
    11'b01001101101: data <= 32'hb942bde8;
    11'b01001101110: data <= 32'h38bbbb91;
    11'b01001101111: data <= 32'h3d273baf;
    11'b01001110000: data <= 32'h3d033eb8;
    11'b01001110001: data <= 32'h3d7c38b8;
    11'b01001110010: data <= 32'h3e61b675;
    11'b01001110011: data <= 32'h3a8ea427;
    11'b01001110100: data <= 32'hbb173888;
    11'b01001110101: data <= 32'hbe85b19a;
    11'b01001110110: data <= 32'hb50abe87;
    11'b01001110111: data <= 32'h3da5c039;
    11'b01001111000: data <= 32'h3d20bd8b;
    11'b01001111001: data <= 32'hb5cfb8f7;
    11'b01001111010: data <= 32'hbcc3b324;
    11'b01001111011: data <= 32'hb6d237bc;
    11'b01001111100: data <= 32'h308a3d98;
    11'b01001111101: data <= 32'hbae03cf9;
    11'b01001111110: data <= 32'hc063b413;
    11'b01001111111: data <= 32'hbfbabd39;
    11'b01010000000: data <= 32'hb499b6b0;
    11'b01010000001: data <= 32'h3b9e3d0b;
    11'b01010000010: data <= 32'h3c6d3e17;
    11'b01010000011: data <= 32'h3c1e3627;
    11'b01010000100: data <= 32'h3c65a74e;
    11'b01010000101: data <= 32'h38c63c67;
    11'b01010000110: data <= 32'hb8083faa;
    11'b01010000111: data <= 32'hba9839af;
    11'b01010001000: data <= 32'h35a9bdcf;
    11'b01010001001: data <= 32'h3e59c097;
    11'b01010001010: data <= 32'h3ce0bdd8;
    11'b01010001011: data <= 32'haad7b811;
    11'b01010001100: data <= 32'hb309b479;
    11'b01010001101: data <= 32'h3a6ead8e;
    11'b01010001110: data <= 32'h3b3436b7;
    11'b01010001111: data <= 32'hbb6e35eb;
    11'b01010010000: data <= 32'hc190b8d6;
    11'b01010010001: data <= 32'hc0ecbd05;
    11'b01010010010: data <= 32'hb848b82a;
    11'b01010010011: data <= 32'h399238f0;
    11'b01010010100: data <= 32'h376a38af;
    11'b01010010101: data <= 32'h2701b0e2;
    11'b01010010110: data <= 32'h32a134a5;
    11'b01010010111: data <= 32'h343c4019;
    11'b01010011000: data <= 32'hb50e41b2;
    11'b01010011001: data <= 32'hb8f53cf2;
    11'b01010011010: data <= 32'h300bbc8f;
    11'b01010011011: data <= 32'h3c21bf0b;
    11'b01010011100: data <= 32'h3b80b8ed;
    11'b01010011101: data <= 32'h372733a1;
    11'b01010011110: data <= 32'h3b8faf21;
    11'b01010011111: data <= 32'h3ff6b82e;
    11'b01010100000: data <= 32'h3e4eb088;
    11'b01010100001: data <= 32'hb99d31f3;
    11'b01010100010: data <= 32'hc113b671;
    11'b01010100011: data <= 32'hbfd1bcb6;
    11'b01010100100: data <= 32'hab85bc5a;
    11'b01010100101: data <= 32'h3921b898;
    11'b01010100110: data <= 32'hb392b929;
    11'b01010100111: data <= 32'hbaf1ba89;
    11'b01010101000: data <= 32'hb5013434;
    11'b01010101001: data <= 32'h337b406b;
    11'b01010101010: data <= 32'hb4e2419a;
    11'b01010101011: data <= 32'hbc6a3c69;
    11'b01010101100: data <= 32'hbb4cbb0f;
    11'b01010101101: data <= 32'ha9f3bb22;
    11'b01010101110: data <= 32'h370b37eb;
    11'b01010101111: data <= 32'h39843bbd;
    11'b01010110000: data <= 32'h3e190911;
    11'b01010110001: data <= 32'h40d1b923;
    11'b01010110010: data <= 32'h3f1f2ddd;
    11'b01010110011: data <= 32'hb51d3b6f;
    11'b01010110100: data <= 32'hbeab3675;
    11'b01010110101: data <= 32'hba9ebb76;
    11'b01010110110: data <= 32'h39afbe76;
    11'b01010110111: data <= 32'h3993be04;
    11'b01010111000: data <= 32'hb8d0bdb4;
    11'b01010111001: data <= 32'hbc15bd05;
    11'b01010111010: data <= 32'h2966b013;
    11'b01010111011: data <= 32'h39e93e0a;
    11'b01010111100: data <= 32'hb49b3f7f;
    11'b01010111101: data <= 32'hbf6237a1;
    11'b01010111110: data <= 32'hc024ba3e;
    11'b01010111111: data <= 32'hbc15b371;
    11'b01011000000: data <= 32'habd33c4c;
    11'b01011000001: data <= 32'h37063c19;
    11'b01011000010: data <= 32'h3c8db3d5;
    11'b01011000011: data <= 32'h3f5eb868;
    11'b01011000100: data <= 32'h3dc03b1f;
    11'b01011000101: data <= 32'h9950404c;
    11'b01011000110: data <= 32'hba063d99;
    11'b01011000111: data <= 32'h2e70b852;
    11'b01011001000: data <= 32'h3c6fbe97;
    11'b01011001001: data <= 32'h38f9be1d;
    11'b01011001010: data <= 32'hb872bd1f;
    11'b01011001011: data <= 32'hb5efbcf3;
    11'b01011001100: data <= 32'h3c86b92e;
    11'b01011001101: data <= 32'h3e763714;
    11'b01011001110: data <= 32'haedc3a1c;
    11'b01011001111: data <= 32'hc07bae48;
    11'b01011010000: data <= 32'hc115b9f3;
    11'b01011010001: data <= 32'hbd18ae20;
    11'b01011010010: data <= 32'hb4c53a00;
    11'b01011010011: data <= 32'hb1ce33be;
    11'b01011010100: data <= 32'h2baebb30;
    11'b01011010101: data <= 32'h39ebb80c;
    11'b01011010110: data <= 32'h3b133e75;
    11'b01011010111: data <= 32'h30af4209;
    11'b01011011000: data <= 32'hb55c3fe1;
    11'b01011011001: data <= 32'h321bb1fc;
    11'b01011011010: data <= 32'h39cdbc67;
    11'b01011011011: data <= 32'h3387b8ed;
    11'b01011011100: data <= 32'hb57ab5b0;
    11'b01011011101: data <= 32'h385dbaea;
    11'b01011011110: data <= 32'h4080bc1d;
    11'b01011011111: data <= 32'h40bdb4e5;
    11'b01011100000: data <= 32'h32e93444;
    11'b01011100001: data <= 32'hbfc9adbd;
    11'b01011100010: data <= 32'hbfe4b8aa;
    11'b01011100011: data <= 32'hb93fb5f9;
    11'b01011100100: data <= 32'hb1a6b186;
    11'b01011100101: data <= 32'hba93bb52;
    11'b01011100110: data <= 32'hbbfdbeae;
    11'b01011100111: data <= 32'had61b975;
    11'b01011101000: data <= 32'h391e3ebf;
    11'b01011101001: data <= 32'h32ca41d4;
    11'b01011101010: data <= 32'hb84a3ef1;
    11'b01011101011: data <= 32'hb87fac54;
    11'b01011101100: data <= 32'hb44ab48a;
    11'b01011101101: data <= 32'hb640391d;
    11'b01011101110: data <= 32'hb4b43950;
    11'b01011101111: data <= 32'h3c02b832;
    11'b01011110000: data <= 32'h413fbcb0;
    11'b01011110001: data <= 32'h4109b575;
    11'b01011110010: data <= 32'h381039af;
    11'b01011110011: data <= 32'hbc7138e5;
    11'b01011110100: data <= 32'hb9bbb273;
    11'b01011110101: data <= 32'h362eb95b;
    11'b01011110110: data <= 32'h2f42bb97;
    11'b01011110111: data <= 32'hbcbebea1;
    11'b01011111000: data <= 32'hbd9bc035;
    11'b01011111001: data <= 32'ha8f6bc24;
    11'b01011111010: data <= 32'h3c103c00;
    11'b01011111011: data <= 32'h35c33f7f;
    11'b01011111100: data <= 32'hbc173ae1;
    11'b01011111101: data <= 32'hbe26b244;
    11'b01011111110: data <= 32'hbcd635b3;
    11'b01011111111: data <= 32'hbb7a3dd0;
    11'b01100000000: data <= 32'hb8863c28;
    11'b01100000001: data <= 32'h38d6b8ea;
    11'b01100000010: data <= 32'h3fd5bcc8;
    11'b01100000011: data <= 32'h3fd7320e;
    11'b01100000100: data <= 32'h38e03ee4;
    11'b01100000101: data <= 32'hb33d3e4d;
    11'b01100000110: data <= 32'h36eb3463;
    11'b01100000111: data <= 32'h3c6fb8ff;
    11'b01100001000: data <= 32'h3309bb78;
    11'b01100001001: data <= 32'hbceebdbe;
    11'b01100001010: data <= 32'hbc1abfa8;
    11'b01100001011: data <= 32'h3a8fbd78;
    11'b01100001100: data <= 32'h3f67a853;
    11'b01100001101: data <= 32'h39393874;
    11'b01100001110: data <= 32'hbd29a979;
    11'b01100001111: data <= 32'hbfc4b5da;
    11'b01100010000: data <= 32'hbda03880;
    11'b01100010001: data <= 32'hbc343d9d;
    11'b01100010010: data <= 32'hbc263812;
    11'b01100010011: data <= 32'hb71abcd9;
    11'b01100010100: data <= 32'h3954bd1e;
    11'b01100010101: data <= 32'h3c5539f8;
    11'b01100010110: data <= 32'h384240ff;
    11'b01100010111: data <= 32'h339d4036;
    11'b01100011000: data <= 32'h3a5e387c;
    11'b01100011001: data <= 32'h3c01b1a8;
    11'b01100011010: data <= 32'hadbea92a;
    11'b01100011011: data <= 32'hbc9eb576;
    11'b01100011100: data <= 32'hb4e7bcef;
    11'b01100011101: data <= 32'h3f4bbe0d;
    11'b01100011110: data <= 32'h412aba76;
    11'b01100011111: data <= 32'h3bb1b2c3;
    11'b01100100000: data <= 32'hbc2db55e;
    11'b01100100001: data <= 32'hbd82b4f8;
    11'b01100100010: data <= 32'hb92436ac;
    11'b01100100011: data <= 32'hb936399e;
    11'b01100100100: data <= 32'hbdcab815;
    11'b01100100101: data <= 32'hbe0dbfe5;
    11'b01100100110: data <= 32'hb6c9bdf3;
    11'b01100100111: data <= 32'h381d3a89;
    11'b01100101000: data <= 32'h375840c4;
    11'b01100101001: data <= 32'h31093f02;
    11'b01100101010: data <= 32'h34913711;
    11'b01100101011: data <= 32'h317e36db;
    11'b01100101100: data <= 32'hb9ab3cde;
    11'b01100101101: data <= 32'hbcb63b7d;
    11'b01100101110: data <= 32'h2e95b86e;
    11'b01100101111: data <= 32'h4057bdf1;
    11'b01100110000: data <= 32'h4148bb91;
    11'b01100110001: data <= 32'h3c3fa69e;
    11'b01100110010: data <= 32'hb6403180;
    11'b01100110011: data <= 32'hafa02b26;
    11'b01100110100: data <= 32'h392b331e;
    11'b01100110101: data <= 32'ha41123e4;
    11'b01100110110: data <= 32'hbe75bcdc;
    11'b01100110111: data <= 32'hc000c0b1;
    11'b01100111000: data <= 32'hb933bece;
    11'b01100111001: data <= 32'h394c3475;
    11'b01100111010: data <= 32'h38943d5c;
    11'b01100111011: data <= 32'hb2b7392c;
    11'b01100111100: data <= 32'hb880a6fd;
    11'b01100111101: data <= 32'hb9ba3ad9;
    11'b01100111110: data <= 32'hbce34034;
    11'b01100111111: data <= 32'hbd753e5f;
    11'b01101000000: data <= 32'hb1f2b618;
    11'b01101000001: data <= 32'h3e02bdc8;
    11'b01101000010: data <= 32'h3f80b854;
    11'b01101000011: data <= 32'h3ab53a9c;
    11'b01101000100: data <= 32'h346c3c3e;
    11'b01101000101: data <= 32'h3c5b3831;
    11'b01101000110: data <= 32'h3ea2338e;
    11'b01101000111: data <= 32'h362ba8b9;
    11'b01101001000: data <= 32'hbe45bbea;
    11'b01101001001: data <= 32'hbefebfed;
    11'b01101001010: data <= 32'h2535bef3;
    11'b01101001011: data <= 32'h3d97b859;
    11'b01101001100: data <= 32'h3af2a78c;
    11'b01101001101: data <= 32'hb767b86c;
    11'b01101001110: data <= 32'hbbf0b829;
    11'b01101001111: data <= 32'hbb473b81;
    11'b01101010000: data <= 32'hbccd4057;
    11'b01101010001: data <= 32'hbe543d1b;
    11'b01101010010: data <= 32'hbc25baca;
    11'b01101010011: data <= 32'h314abe21;
    11'b01101010100: data <= 32'h399ea859;
    11'b01101010101: data <= 32'h36ab3e5b;
    11'b01101010110: data <= 32'h38b63e57;
    11'b01101010111: data <= 32'h3e4539b3;
    11'b01101011000: data <= 32'h3f2c37a8;
    11'b01101011001: data <= 32'h33ba3974;
    11'b01101011010: data <= 32'hbded3089;
    11'b01101011011: data <= 32'hbc6abc10;
    11'b01101011100: data <= 32'h3bcebe1c;
    11'b01101011101: data <= 32'h403bbc93;
    11'b01101011110: data <= 32'h3c75bb44;
    11'b01101011111: data <= 32'hb5e7bc76;
    11'b01101100000: data <= 32'hb897b95f;
    11'b01101100001: data <= 32'haf7b3a23;
    11'b01101100010: data <= 32'hb84f3e40;
    11'b01101100011: data <= 32'hbe923569;
    11'b01101100100: data <= 32'hbfabbe59;
    11'b01101100101: data <= 32'hbc1ebed5;
    11'b01101100110: data <= 32'hb12d307d;
    11'b01101100111: data <= 32'h2e033e5c;
    11'b01101101000: data <= 32'h37553cd8;
    11'b01101101001: data <= 32'h3ca835ca;
    11'b01101101010: data <= 32'h3c513a09;
    11'b01101101011: data <= 32'hb5653efe;
    11'b01101101100: data <= 32'hbdfb3e13;
    11'b01101101101: data <= 32'hb915a5e2;
    11'b01101101110: data <= 32'h3da4bcd8;
    11'b01101101111: data <= 32'h4054bcd0;
    11'b01101110000: data <= 32'h3c15bab9;
    11'b01101110001: data <= 32'ha33fba19;
    11'b01101110010: data <= 32'h37fab5f2;
    11'b01101110011: data <= 32'h3d0f3899;
    11'b01101110100: data <= 32'h36b33ad9;
    11'b01101110101: data <= 32'hbdf5b6d1;
    11'b01101110110: data <= 32'hc099bfd8;
    11'b01101110111: data <= 32'hbd85bf13;
    11'b01101111000: data <= 32'hb2acb064;
    11'b01101111001: data <= 32'h2ea039c2;
    11'b01101111010: data <= 32'h2e032537;
    11'b01101111011: data <= 32'h354bb6d9;
    11'b01101111100: data <= 32'h31273abf;
    11'b01101111101: data <= 32'hbae34102;
    11'b01101111110: data <= 32'hbe48409c;
    11'b01101111111: data <= 32'hb9a33624;
    11'b01110000000: data <= 32'h3b39bc18;
    11'b01110000001: data <= 32'h3d4eba54;
    11'b01110000010: data <= 32'h37cfa80d;
    11'b01110000011: data <= 32'h34ee2fe5;
    11'b01110000100: data <= 32'h3e432ee1;
    11'b01110000101: data <= 32'h40d33820;
    11'b01110000110: data <= 32'h3c5c3905;
    11'b01110000111: data <= 32'hbcffb592;
    11'b01110001000: data <= 32'hc00bbe2a;
    11'b01110001001: data <= 32'hba37be12;
    11'b01110001010: data <= 32'h37c6b8f5;
    11'b01110001011: data <= 32'h3667b802;
    11'b01110001100: data <= 32'hb26ebd47;
    11'b01110001101: data <= 32'hb36abce4;
    11'b01110001110: data <= 32'hb1483986;
    11'b01110001111: data <= 32'hba77410f;
    11'b01110010000: data <= 32'hbe244027;
    11'b01110010001: data <= 32'hbcec97f3;
    11'b01110010010: data <= 32'hb480bc5b;
    11'b01110010011: data <= 32'h21dbb42b;
    11'b01110010100: data <= 32'hb4283a99;
    11'b01110010101: data <= 32'h35953a19;
    11'b01110010110: data <= 32'h3fee3495;
    11'b01110010111: data <= 32'h41503863;
    11'b01110011000: data <= 32'h3c4a3c30;
    11'b01110011001: data <= 32'hbc723906;
    11'b01110011010: data <= 32'hbd73b711;
    11'b01110011011: data <= 32'h339bbbc1;
    11'b01110011100: data <= 32'h3d30bb59;
    11'b01110011101: data <= 32'h393cbd36;
    11'b01110011110: data <= 32'hb462c006;
    11'b01110011111: data <= 32'had20be32;
    11'b01110100000: data <= 32'h379136e4;
    11'b01110100001: data <= 32'ha71f3fa1;
    11'b01110100010: data <= 32'hbd083c70;
    11'b01110100011: data <= 32'hbf2bba74;
    11'b01110100100: data <= 32'hbd8cbd21;
    11'b01110100101: data <= 32'hbc04295a;
    11'b01110100110: data <= 32'hba753c3c;
    11'b01110100111: data <= 32'h2d963853;
    11'b01110101000: data <= 32'h3e40b11f;
    11'b01110101001: data <= 32'h3fc83806;
    11'b01110101010: data <= 32'h37553f26;
    11'b01110101011: data <= 32'hbc923f9d;
    11'b01110101100: data <= 32'hba6239be;
    11'b01110101101: data <= 32'h3afbb61d;
    11'b01110101110: data <= 32'h3dfbba6d;
    11'b01110101111: data <= 32'h37d5bcd9;
    11'b01110110000: data <= 32'hb2d5beca;
    11'b01110110001: data <= 32'h395fbd03;
    11'b01110110010: data <= 32'h3efb33ed;
    11'b01110110011: data <= 32'h3c6a3c85;
    11'b01110110100: data <= 32'hba643198;
    11'b01110110101: data <= 32'hbfd4bd50;
    11'b01110110110: data <= 32'hbed3bd32;
    11'b01110110111: data <= 32'hbc7f26a6;
    11'b01110111000: data <= 32'hbacf37f2;
    11'b01110111001: data <= 32'hb49db846;
    11'b01110111010: data <= 32'h396cbc7d;
    11'b01110111011: data <= 32'h3b1b3438;
    11'b01110111100: data <= 32'hb2954097;
    11'b01110111101: data <= 32'hbcce414d;
    11'b01110111110: data <= 32'hb91f3cee;
    11'b01110111111: data <= 32'h3944ad83;
    11'b01111000000: data <= 32'h3a3db591;
    11'b01111000001: data <= 32'hb295b5d8;
    11'b01111000010: data <= 32'hb352b9a8;
    11'b01111000011: data <= 32'h3ddeb930;
    11'b01111000100: data <= 32'h41b2322f;
    11'b01111000101: data <= 32'h3fa839b0;
    11'b01111000110: data <= 32'hb653a5e7;
    11'b01111000111: data <= 32'hbe65bc2c;
    11'b01111001000: data <= 32'hbc48bb3c;
    11'b01111001001: data <= 32'hb5ceafbe;
    11'b01111001010: data <= 32'hb748b706;
    11'b01111001011: data <= 32'hb888bf4c;
    11'b01111001100: data <= 32'ha950c02b;
    11'b01111001101: data <= 32'h34e3aea1;
    11'b01111001110: data <= 32'hb4ce4066;
    11'b01111001111: data <= 32'hbc3340c9;
    11'b01111010000: data <= 32'hbac03a8e;
    11'b01111010001: data <= 32'hb371b2d9;
    11'b01111010010: data <= 32'hb7a93159;
    11'b01111010011: data <= 32'hbc9038f3;
    11'b01111010100: data <= 32'hb724314d;
    11'b01111010101: data <= 32'h3eebb4fa;
    11'b01111010110: data <= 32'h42223087;
    11'b01111010111: data <= 32'h3fa53aa3;
    11'b01111011000: data <= 32'hb466393f;
    11'b01111011001: data <= 32'hbb89a0e1;
    11'b01111011010: data <= 32'h2a4cb106;
    11'b01111011011: data <= 32'h3941b00c;
    11'b01111011100: data <= 32'ha8febc39;
    11'b01111011101: data <= 32'hb98ac100;
    11'b01111011110: data <= 32'hb138c0f0;
    11'b01111011111: data <= 32'h392cb65d;
    11'b01111100000: data <= 32'h365b3e3d;
    11'b01111100001: data <= 32'hb89c3d5c;
    11'b01111100010: data <= 32'hbc59b14c;
    11'b01111100011: data <= 32'hbc82b882;
    11'b01111100100: data <= 32'hbdef37f5;
    11'b01111100101: data <= 32'hbf2d3c63;
    11'b01111100110: data <= 32'hba613391;
    11'b01111100111: data <= 32'h3d10b93d;
    11'b01111101000: data <= 32'h4092ad6f;
    11'b01111101001: data <= 32'h3c9a3cf8;
    11'b01111101010: data <= 32'hb72c3ecc;
    11'b01111101011: data <= 32'hb5da3c91;
    11'b01111101100: data <= 32'h3b37389e;
    11'b01111101101: data <= 32'h3c903050;
    11'b01111101110: data <= 32'had27bb27;
    11'b01111101111: data <= 32'hba50c044;
    11'b01111110000: data <= 32'h3437c023;
    11'b01111110001: data <= 32'h3eaeb76c;
    11'b01111110010: data <= 32'h3e113a3a;
    11'b01111110011: data <= 32'h2bf932ba;
    11'b01111110100: data <= 32'hbc39bbb8;
    11'b01111110101: data <= 32'hbd62b9c8;
    11'b01111110110: data <= 32'hbe4838e2;
    11'b01111110111: data <= 32'hbf213acc;
    11'b01111111000: data <= 32'hbc5fb89f;
    11'b01111111001: data <= 32'h3607be63;
    11'b01111111010: data <= 32'h3c39b82f;
    11'b01111111011: data <= 32'h33063e0a;
    11'b01111111100: data <= 32'hb95140a3;
    11'b01111111101: data <= 32'haedf3e91;
    11'b01111111110: data <= 32'h3bea3afa;
    11'b01111111111: data <= 32'h39933876;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    