
module memory_rom_55(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3b4dbd26;
    11'b00000000001: data <= 32'h37beba74;
    11'b00000000010: data <= 32'hb82e39ac;
    11'b00000000011: data <= 32'hbe853b54;
    11'b00000000100: data <= 32'hbe1aba5a;
    11'b00000000101: data <= 32'hb4eac0a4;
    11'b00000000110: data <= 32'h34b3bf74;
    11'b00000000111: data <= 32'hb7aeb3ce;
    11'b00000001000: data <= 32'hbc8039f2;
    11'b00000001001: data <= 32'hb45d3b45;
    11'b00000001010: data <= 32'h3b613cd6;
    11'b00000001011: data <= 32'h36693e71;
    11'b00000001100: data <= 32'hbdee3cb5;
    11'b00000001101: data <= 32'hc05c2c2e;
    11'b00000001110: data <= 32'hb873b5c3;
    11'b00000001111: data <= 32'h3e383434;
    11'b00000010000: data <= 32'h401c388d;
    11'b00000010001: data <= 32'h3d2ab3ec;
    11'b00000010010: data <= 32'h3aecbaf9;
    11'b00000010011: data <= 32'h3bdb2d81;
    11'b00000010100: data <= 32'h38bb3e16;
    11'b00000010101: data <= 32'hb6143c73;
    11'b00000010110: data <= 32'hba2ebcc2;
    11'b00000010111: data <= 32'hb40ec1a7;
    11'b00000011000: data <= 32'h2b71c042;
    11'b00000011001: data <= 32'hb68bb705;
    11'b00000011010: data <= 32'hb8b4316c;
    11'b00000011011: data <= 32'h3488b222;
    11'b00000011100: data <= 32'h3b5695a2;
    11'b00000011101: data <= 32'hb4433b67;
    11'b00000011110: data <= 32'hc0b43d1c;
    11'b00000011111: data <= 32'hc18738be;
    11'b00000100000: data <= 32'hbaf2a677;
    11'b00000100001: data <= 32'h3c573037;
    11'b00000100010: data <= 32'h3cab34c9;
    11'b00000100011: data <= 32'h349ead84;
    11'b00000100100: data <= 32'h3613acc2;
    11'b00000100101: data <= 32'h3d573c8d;
    11'b00000100110: data <= 32'h3dd9408a;
    11'b00000100111: data <= 32'h35983da4;
    11'b00000101000: data <= 32'hb86fbbd2;
    11'b00000101001: data <= 32'hb506c0a5;
    11'b00000101010: data <= 32'h344ebde7;
    11'b00000101011: data <= 32'h35a3b2c9;
    11'b00000101100: data <= 32'h36f5b6d7;
    11'b00000101101: data <= 32'h3c06bd71;
    11'b00000101110: data <= 32'h3c50bc31;
    11'b00000101111: data <= 32'hb64537b5;
    11'b00000110000: data <= 32'hc0a43d23;
    11'b00000110001: data <= 32'hc11137e2;
    11'b00000110010: data <= 32'hbb30b8b4;
    11'b00000110011: data <= 32'h3585b983;
    11'b00000110100: data <= 32'hb0d5b3ab;
    11'b00000110101: data <= 32'hbb6ca552;
    11'b00000110110: data <= 32'hb0a63655;
    11'b00000110111: data <= 32'h3dce3e31;
    11'b00000111000: data <= 32'h3e9340db;
    11'b00000111001: data <= 32'h301c3e89;
    11'b00000111010: data <= 32'hbc4ab39a;
    11'b00000111011: data <= 32'hb8d8bc44;
    11'b00000111100: data <= 32'h389cb4a6;
    11'b00000111101: data <= 32'h3c7033fd;
    11'b00000111110: data <= 32'h3ca8ba1a;
    11'b00000111111: data <= 32'h3dacbfbc;
    11'b00001000000: data <= 32'h3d78bd0a;
    11'b00001000001: data <= 32'h32643954;
    11'b00001000010: data <= 32'hbd483d7b;
    11'b00001000011: data <= 32'hbe502837;
    11'b00001000100: data <= 32'hb903be0b;
    11'b00001000101: data <= 32'hb3efbe51;
    11'b00001000110: data <= 32'hbc75b9cb;
    11'b00001000111: data <= 32'hbe49b2c0;
    11'b00001001000: data <= 32'hb42b2da3;
    11'b00001001001: data <= 32'h3dc23b71;
    11'b00001001010: data <= 32'h3cd03f4f;
    11'b00001001011: data <= 32'hba343e80;
    11'b00001001100: data <= 32'hbfd438b2;
    11'b00001001101: data <= 32'hbc0731df;
    11'b00001001110: data <= 32'h3903395a;
    11'b00001001111: data <= 32'h3cc03881;
    11'b00001010000: data <= 32'h3bd5ba45;
    11'b00001010001: data <= 32'h3cbbbecf;
    11'b00001010010: data <= 32'h3e67b8a7;
    11'b00001010011: data <= 32'h3cae3d8e;
    11'b00001010100: data <= 32'h2b023e66;
    11'b00001010101: data <= 32'hb7ecb4f4;
    11'b00001010110: data <= 32'hb46bc000;
    11'b00001010111: data <= 32'hb6d6bf3b;
    11'b00001011000: data <= 32'hbceaba33;
    11'b00001011001: data <= 32'hbd1ab883;
    11'b00001011010: data <= 32'h31cabb0d;
    11'b00001011011: data <= 32'h3de6b64c;
    11'b00001011100: data <= 32'h39033a89;
    11'b00001011101: data <= 32'hbe633da3;
    11'b00001011110: data <= 32'hc1053c21;
    11'b00001011111: data <= 32'hbce1399f;
    11'b00001100000: data <= 32'h353e3a7a;
    11'b00001100001: data <= 32'h3688370b;
    11'b00001100010: data <= 32'haff9b949;
    11'b00001100011: data <= 32'h3630bc18;
    11'b00001100100: data <= 32'h3e863649;
    11'b00001100101: data <= 32'h3fc24038;
    11'b00001100110: data <= 32'h3bba3f5d;
    11'b00001100111: data <= 32'h25e3b2ee;
    11'b00001101000: data <= 32'hb0d6be56;
    11'b00001101001: data <= 32'hb3bfbc43;
    11'b00001101010: data <= 32'hb8e2b436;
    11'b00001101011: data <= 32'hb5cdbac4;
    11'b00001101100: data <= 32'h3b00bfc0;
    11'b00001101101: data <= 32'h3e78be78;
    11'b00001101110: data <= 32'h36e42a3d;
    11'b00001101111: data <= 32'hbe853cc3;
    11'b00001110000: data <= 32'hc06a3b81;
    11'b00001110001: data <= 32'hbbfe34d2;
    11'b00001110010: data <= 32'haf953046;
    11'b00001110011: data <= 32'hba5cab8b;
    11'b00001110100: data <= 32'hbe0eb8d9;
    11'b00001110101: data <= 32'hb7adb83c;
    11'b00001110110: data <= 32'h3df13ac1;
    11'b00001110111: data <= 32'h4034406f;
    11'b00001111000: data <= 32'h3b5b3f6c;
    11'b00001111001: data <= 32'hb4fe3427;
    11'b00001111010: data <= 32'hb615b704;
    11'b00001111011: data <= 32'h28903493;
    11'b00001111100: data <= 32'h30213862;
    11'b00001111101: data <= 32'h362dbb27;
    11'b00001111110: data <= 32'h3d05c0f2;
    11'b00001111111: data <= 32'h3efbc008;
    11'b00010000000: data <= 32'h3a5c21f5;
    11'b00010000001: data <= 32'hb9de3cb9;
    11'b00010000010: data <= 32'hbc63381b;
    11'b00010000011: data <= 32'hb613b889;
    11'b00010000100: data <= 32'hb687b9fe;
    11'b00010000101: data <= 32'hbed2b838;
    11'b00010000110: data <= 32'hc0b5b978;
    11'b00010000111: data <= 32'hbad7b938;
    11'b00010001000: data <= 32'h3d5e352e;
    11'b00010001001: data <= 32'h3ec63dea;
    11'b00010001010: data <= 32'h2e673e0e;
    11'b00010001011: data <= 32'hbca33a33;
    11'b00010001100: data <= 32'hba2f39fb;
    11'b00010001101: data <= 32'h30f43dcf;
    11'b00010001110: data <= 32'h358f3ca2;
    11'b00010001111: data <= 32'h34a1b9f4;
    11'b00010010000: data <= 32'h3b46c086;
    11'b00010010001: data <= 32'h3eb1bdca;
    11'b00010010010: data <= 32'h3dd9394e;
    11'b00010010011: data <= 32'h388f3d98;
    11'b00010010100: data <= 32'h326e305c;
    11'b00010010101: data <= 32'h34cebc9f;
    11'b00010010110: data <= 32'hb611bc38;
    11'b00010010111: data <= 32'hbf52b7f1;
    11'b00010011000: data <= 32'hc064ba29;
    11'b00010011001: data <= 32'hb82fbd58;
    11'b00010011010: data <= 32'h3d67bb62;
    11'b00010011011: data <= 32'h3c6d3412;
    11'b00010011100: data <= 32'hba413b8e;
    11'b00010011101: data <= 32'hbf1c3bd4;
    11'b00010011110: data <= 32'hbb723d12;
    11'b00010011111: data <= 32'h2cf23f09;
    11'b00010100000: data <= 32'hb1843cc2;
    11'b00010100001: data <= 32'hb9dfb893;
    11'b00010100010: data <= 32'hadcbbe5c;
    11'b00010100011: data <= 32'h3d5cb72a;
    11'b00010100100: data <= 32'h3fdb3dbc;
    11'b00010100101: data <= 32'h3de33e6e;
    11'b00010100110: data <= 32'h3b4c2ac4;
    11'b00010100111: data <= 32'h3907bbbe;
    11'b00010101000: data <= 32'haf48b653;
    11'b00010101001: data <= 32'hbce9326b;
    11'b00010101010: data <= 32'hbd2ab98e;
    11'b00010101011: data <= 32'h326ac038;
    11'b00010101100: data <= 32'h3debc042;
    11'b00010101101: data <= 32'h3a34b9d7;
    11'b00010101110: data <= 32'hbc0d3791;
    11'b00010101111: data <= 32'hbe3c3a22;
    11'b00010110000: data <= 32'hb8653b1a;
    11'b00010110001: data <= 32'ha7a53c83;
    11'b00010110010: data <= 32'hbc5d3984;
    11'b00010110011: data <= 32'hc032b81a;
    11'b00010110100: data <= 32'hbcc2bbfc;
    11'b00010110101: data <= 32'h3b333184;
    11'b00010110110: data <= 32'h3fe33e83;
    11'b00010110111: data <= 32'h3dc93df7;
    11'b00010111000: data <= 32'h394b32f4;
    11'b00010111001: data <= 32'h3702ae65;
    11'b00010111010: data <= 32'h317b3b69;
    11'b00010111011: data <= 32'hb6c63d03;
    11'b00010111100: data <= 32'hb679b6a6;
    11'b00010111101: data <= 32'h3961c0e9;
    11'b00010111110: data <= 32'h3e0bc118;
    11'b00010111111: data <= 32'h3ae6bb20;
    11'b00011000000: data <= 32'hb625360a;
    11'b00011000001: data <= 32'hb7bf351b;
    11'b00011000010: data <= 32'h34fea535;
    11'b00011000011: data <= 32'h274f3082;
    11'b00011000100: data <= 32'hbf253035;
    11'b00011000101: data <= 32'hc1ebb836;
    11'b00011000110: data <= 32'hbee7bb0d;
    11'b00011000111: data <= 32'h38f3adff;
    11'b00011001000: data <= 32'h3e0f3b81;
    11'b00011001001: data <= 32'h38d93b58;
    11'b00011001010: data <= 32'hb4113603;
    11'b00011001011: data <= 32'ha8123ad5;
    11'b00011001100: data <= 32'h353b403b;
    11'b00011001101: data <= 32'h9da9401f;
    11'b00011001110: data <= 32'hb434acec;
    11'b00011001111: data <= 32'h363cc056;
    11'b00011010000: data <= 32'h3ceabfe3;
    11'b00011010001: data <= 32'h3cb4b2b0;
    11'b00011010010: data <= 32'h39673931;
    11'b00011010011: data <= 32'h3ab2ad05;
    11'b00011010100: data <= 32'h3ce2ba2c;
    11'b00011010101: data <= 32'h34b5b625;
    11'b00011010110: data <= 32'hbf3a2d4d;
    11'b00011010111: data <= 32'hc19db6f8;
    11'b00011011000: data <= 32'hbd9fbce8;
    11'b00011011001: data <= 32'h3932bc5b;
    11'b00011011010: data <= 32'h3b49b4e3;
    11'b00011011011: data <= 32'hb6862e28;
    11'b00011011100: data <= 32'hbc4734cb;
    11'b00011011101: data <= 32'hb4863cf7;
    11'b00011011110: data <= 32'h364540e2;
    11'b00011011111: data <= 32'hb2bf404d;
    11'b00011100000: data <= 32'hbc212f4c;
    11'b00011100001: data <= 32'hb8f3bde7;
    11'b00011100010: data <= 32'h3910baed;
    11'b00011100011: data <= 32'h3d7439e3;
    11'b00011100100: data <= 32'h3dae3bab;
    11'b00011100101: data <= 32'h3e56b454;
    11'b00011100110: data <= 32'h3ea2baf5;
    11'b00011100111: data <= 32'h390325e1;
    11'b00011101000: data <= 32'hbcb03a2e;
    11'b00011101001: data <= 32'hbf48ae75;
    11'b00011101010: data <= 32'hb849beab;
    11'b00011101011: data <= 32'h3b06c03c;
    11'b00011101100: data <= 32'h37febd5a;
    11'b00011101101: data <= 32'hbb2ab846;
    11'b00011101110: data <= 32'hbc67a822;
    11'b00011101111: data <= 32'h2c9a3a81;
    11'b00011110000: data <= 32'h38393f07;
    11'b00011110001: data <= 32'hba513e28;
    11'b00011110010: data <= 32'hc0682d46;
    11'b00011110011: data <= 32'hbf18ba99;
    11'b00011110100: data <= 32'ha0daa3b8;
    11'b00011110101: data <= 32'h3ccb3cb5;
    11'b00011110110: data <= 32'h3d4e3b20;
    11'b00011110111: data <= 32'h3d38b538;
    11'b00011111000: data <= 32'h3d9cb56b;
    11'b00011111001: data <= 32'h3abd3c8f;
    11'b00011111010: data <= 32'hb52c3f88;
    11'b00011111011: data <= 32'hb9d6369d;
    11'b00011111100: data <= 32'h31b0bf2c;
    11'b00011111101: data <= 32'h3bd9c0e4;
    11'b00011111110: data <= 32'h364ebdfd;
    11'b00011111111: data <= 32'hb8c2b8ef;
    11'b00100000000: data <= 32'hb3bab71e;
    11'b00100000001: data <= 32'h3be3b03d;
    11'b00100000010: data <= 32'h3abd38be;
    11'b00100000011: data <= 32'hbceb3a02;
    11'b00100000100: data <= 32'hc1e9a606;
    11'b00100000101: data <= 32'hc0abb860;
    11'b00100000110: data <= 32'hb5592883;
    11'b00100000111: data <= 32'h39dc39b5;
    11'b00100001000: data <= 32'h3726346f;
    11'b00100001001: data <= 32'h33c1b6ee;
    11'b00100001010: data <= 32'h39c83553;
    11'b00100001011: data <= 32'h3b27406a;
    11'b00100001100: data <= 32'h333c417a;
    11'b00100001101: data <= 32'hb4943acd;
    11'b00100001110: data <= 32'h3054bdcc;
    11'b00100001111: data <= 32'h3971bf4c;
    11'b00100010000: data <= 32'h371bb997;
    11'b00100010001: data <= 32'h3136b15c;
    11'b00100010010: data <= 32'h3b92b9ea;
    11'b00100010011: data <= 32'h3fdcbbec;
    11'b00100010100: data <= 32'h3d07b2ec;
    11'b00100010101: data <= 32'hbc953732;
    11'b00100010110: data <= 32'hc17f2b71;
    11'b00100010111: data <= 32'hbfb7b921;
    11'b00100011000: data <= 32'hb14fb92b;
    11'b00100011001: data <= 32'h32fdb61e;
    11'b00100011010: data <= 32'hb93fb906;
    11'b00100011011: data <= 32'hbab4b99f;
    11'b00100011100: data <= 32'h32cb3897;
    11'b00100011101: data <= 32'h3b5c40f2;
    11'b00100011110: data <= 32'h33fb418f;
    11'b00100011111: data <= 32'hb9e33b9e;
    11'b00100100000: data <= 32'hb9a7ba93;
    11'b00100100001: data <= 32'h97e5b91e;
    11'b00100100010: data <= 32'h367637d7;
    11'b00100100011: data <= 32'h39c7366c;
    11'b00100100100: data <= 32'h3e83baf1;
    11'b00100100101: data <= 32'h40c9bd2b;
    11'b00100100110: data <= 32'h3e39b02b;
    11'b00100100111: data <= 32'hb85d3b9e;
    11'b00100101000: data <= 32'hbec43782;
    11'b00100101001: data <= 32'hbab7baaa;
    11'b00100101010: data <= 32'h3502bdd1;
    11'b00100101011: data <= 32'haf2dbd5f;
    11'b00100101100: data <= 32'hbd4dbd27;
    11'b00100101101: data <= 32'hbcc0bc3e;
    11'b00100101110: data <= 32'h35b93092;
    11'b00100101111: data <= 32'h3c743ee4;
    11'b00100110000: data <= 32'haca13fea;
    11'b00100110001: data <= 32'hbea43982;
    11'b00100110010: data <= 32'hbf1eb429;
    11'b00100110011: data <= 32'hb9a835fa;
    11'b00100110100: data <= 32'h30f43cfd;
    11'b00100110101: data <= 32'h38b13884;
    11'b00100110110: data <= 32'h3d29bba5;
    11'b00100110111: data <= 32'h3ff1bc10;
    11'b00100111000: data <= 32'h3e4839c2;
    11'b00100111001: data <= 32'h32e43fdf;
    11'b00100111010: data <= 32'hb7453c46;
    11'b00100111011: data <= 32'h31feba96;
    11'b00100111100: data <= 32'h3955bece;
    11'b00100111101: data <= 32'hb322bdcd;
    11'b00100111110: data <= 32'hbd16bd0f;
    11'b00100111111: data <= 32'hb8e4bd44;
    11'b00101000000: data <= 32'h3ca4b9cd;
    11'b00101000001: data <= 32'h3e1836d9;
    11'b00101000010: data <= 32'hb5633b18;
    11'b00101000011: data <= 32'hc0973510;
    11'b00101000100: data <= 32'hc0969a2a;
    11'b00101000101: data <= 32'hbbc93949;
    11'b00101000110: data <= 32'hb2a83c55;
    11'b00101000111: data <= 32'hb3962d65;
    11'b00101001000: data <= 32'h2f22bca3;
    11'b00101001001: data <= 32'h3c16b863;
    11'b00101001010: data <= 32'h3d673e8f;
    11'b00101001011: data <= 32'h39c3418f;
    11'b00101001100: data <= 32'h32dd3df7;
    11'b00101001101: data <= 32'h375db835;
    11'b00101001110: data <= 32'h3839bc6f;
    11'b00101001111: data <= 32'hb42db865;
    11'b00101010000: data <= 32'hb9e8b87a;
    11'b00101010001: data <= 32'h366bbd64;
    11'b00101010010: data <= 32'h4031be17;
    11'b00101010011: data <= 32'h3fddb8bf;
    11'b00101010100: data <= 32'hb3d33418;
    11'b00101010101: data <= 32'hc02d3289;
    11'b00101010110: data <= 32'hbf34a709;
    11'b00101010111: data <= 32'hb8b032f7;
    11'b00101011000: data <= 32'hb7b8320c;
    11'b00101011001: data <= 32'hbd18ba33;
    11'b00101011010: data <= 32'hbcacbdf7;
    11'b00101011011: data <= 32'h3188b5dc;
    11'b00101011100: data <= 32'h3c9b3f85;
    11'b00101011101: data <= 32'h3a4f4180;
    11'b00101011110: data <= 32'h21663dad;
    11'b00101011111: data <= 32'hb0ddaea5;
    11'b00101100000: data <= 32'hae192313;
    11'b00101100001: data <= 32'hb6363a9c;
    11'b00101100010: data <= 32'hb4893590;
    11'b00101100011: data <= 32'h3c20bce8;
    11'b00101100100: data <= 32'h40f2bf61;
    11'b00101100101: data <= 32'h4047ba0a;
    11'b00101100110: data <= 32'h322537fd;
    11'b00101100111: data <= 32'hbc553843;
    11'b00101101000: data <= 32'hb84bafb3;
    11'b00101101001: data <= 32'h3329b729;
    11'b00101101010: data <= 32'hb867b98f;
    11'b00101101011: data <= 32'hbfc5bd9c;
    11'b00101101100: data <= 32'hbf0fbf1a;
    11'b00101101101: data <= 32'h280cb972;
    11'b00101101110: data <= 32'h3ced3cac;
    11'b00101101111: data <= 32'h38843f2c;
    11'b00101110000: data <= 32'hb9eb3abc;
    11'b00101110001: data <= 32'hbc7b322a;
    11'b00101110010: data <= 32'hba3e3c0c;
    11'b00101110011: data <= 32'hb8eb3f52;
    11'b00101110100: data <= 32'hb5a53a96;
    11'b00101110101: data <= 32'h39c3bcac;
    11'b00101110110: data <= 32'h3fbcbe9f;
    11'b00101110111: data <= 32'h3f7bae75;
    11'b00101111000: data <= 32'h39913d86;
    11'b00101111001: data <= 32'h302e3c75;
    11'b00101111010: data <= 32'h39e3adc7;
    11'b00101111011: data <= 32'h3b4db9b0;
    11'b00101111100: data <= 32'hb7b1ba81;
    11'b00101111101: data <= 32'hbfd8bd1a;
    11'b00101111110: data <= 32'hbd9cbf28;
    11'b00101111111: data <= 32'h395cbd40;
    11'b00110000000: data <= 32'h3e78ae4f;
    11'b00110000001: data <= 32'h35a23756;
    11'b00110000010: data <= 32'hbd632f85;
    11'b00110000011: data <= 32'hbe8333a9;
    11'b00110000100: data <= 32'hbbc73d6e;
    11'b00110000101: data <= 32'hba4a3f97;
    11'b00110000110: data <= 32'hbbc43853;
    11'b00110000111: data <= 32'hb6dcbd53;
    11'b00110001000: data <= 32'h39e9bd0a;
    11'b00110001001: data <= 32'h3d2a3a04;
    11'b00110001010: data <= 32'h3bbb4057;
    11'b00110001011: data <= 32'h3ac13df6;
    11'b00110001100: data <= 32'h3d082c66;
    11'b00110001101: data <= 32'h3c09b490;
    11'b00110001110: data <= 32'hb7442b75;
    11'b00110001111: data <= 32'hbe0bb5c0;
    11'b00110010000: data <= 32'hb7dabde1;
    11'b00110010001: data <= 32'h3e43bf72;
    11'b00110010010: data <= 32'h4011bc9b;
    11'b00110010011: data <= 32'h35b3b6fe;
    11'b00110010100: data <= 32'hbd10b452;
    11'b00110010101: data <= 32'hbca62f9b;
    11'b00110010110: data <= 32'hb6693c02;
    11'b00110010111: data <= 32'hb9da3c8b;
    11'b00110011000: data <= 32'hbf08b415;
    11'b00110011001: data <= 32'hbeebbe9b;
    11'b00110011010: data <= 32'hb628bc23;
    11'b00110011011: data <= 32'h3a3b3c50;
    11'b00110011100: data <= 32'h3b3b4054;
    11'b00110011101: data <= 32'h39d03d0e;
    11'b00110011110: data <= 32'h3a7b3243;
    11'b00110011111: data <= 32'h37ab38ca;
    11'b00110100000: data <= 32'hb89b3dcc;
    11'b00110100001: data <= 32'hbc343a9d;
    11'b00110100010: data <= 32'h3212bc08;
    11'b00110100011: data <= 32'h3fdbc009;
    11'b00110100100: data <= 32'h402cbd94;
    11'b00110100101: data <= 32'h384fb63d;
    11'b00110100110: data <= 32'hb7aeacb6;
    11'b00110100111: data <= 32'h2f3122fb;
    11'b00110101000: data <= 32'h397935cf;
    11'b00110101001: data <= 32'hb7123398;
    11'b00110101010: data <= 32'hc078bb37;
    11'b00110101011: data <= 32'hc0cebf6a;
    11'b00110101100: data <= 32'hba05bc90;
    11'b00110101101: data <= 32'h39753883;
    11'b00110101110: data <= 32'h39303cce;
    11'b00110101111: data <= 32'h266736c7;
    11'b00110110000: data <= 32'hb05b302e;
    11'b00110110001: data <= 32'hb2ea3d8d;
    11'b00110110010: data <= 32'hba06410c;
    11'b00110110011: data <= 32'hbbb03e39;
    11'b00110110100: data <= 32'h2a8ab9cf;
    11'b00110110101: data <= 32'h3db6bf15;
    11'b00110110110: data <= 32'h3e4eba6e;
    11'b00110110111: data <= 32'h398336eb;
    11'b00110111000: data <= 32'h38223801;
    11'b00110111001: data <= 32'h3dd124ee;
    11'b00110111010: data <= 32'h3e9ba2c2;
    11'b00110111011: data <= 32'haee6a6ae;
    11'b00110111100: data <= 32'hc055ba54;
    11'b00110111101: data <= 32'hc039bea1;
    11'b00110111110: data <= 32'hb2c1bdc1;
    11'b00110111111: data <= 32'h3c22b7bf;
    11'b00111000000: data <= 32'h36c9b25c;
    11'b00111000001: data <= 32'hb93ab8c9;
    11'b00111000010: data <= 32'hba15afff;
    11'b00111000011: data <= 32'hb6f83e7a;
    11'b00111000100: data <= 32'hba094158;
    11'b00111000101: data <= 32'hbd1b3da3;
    11'b00111000110: data <= 32'hbb11ba90;
    11'b00111000111: data <= 32'h3190bd74;
    11'b00111001000: data <= 32'h39872d98;
    11'b00111001001: data <= 32'h39053d3b;
    11'b00111001010: data <= 32'h3c5e3b4b;
    11'b00111001011: data <= 32'h40222a4e;
    11'b00111001100: data <= 32'h3fb430c9;
    11'b00111001101: data <= 32'h2776391f;
    11'b00111001110: data <= 32'hbeca3181;
    11'b00111001111: data <= 32'hbcc1bc24;
    11'b00111010000: data <= 32'h39ebbe8c;
    11'b00111010001: data <= 32'h3df2bd84;
    11'b00111010010: data <= 32'h355ebcc7;
    11'b00111010011: data <= 32'hba5bbcd3;
    11'b00111010100: data <= 32'hb7c4b670;
    11'b00111010101: data <= 32'h31553cec;
    11'b00111010110: data <= 32'hb6a43fb2;
    11'b00111010111: data <= 32'hbed638bb;
    11'b00111011000: data <= 32'hc006bcaf;
    11'b00111011001: data <= 32'hbc39bc4d;
    11'b00111011010: data <= 32'had3638c6;
    11'b00111011011: data <= 32'h35be3dea;
    11'b00111011100: data <= 32'h3b623961;
    11'b00111011101: data <= 32'h3ea1ad2a;
    11'b00111011110: data <= 32'h3da73983;
    11'b00111011111: data <= 32'haecd3f66;
    11'b00111100000: data <= 32'hbcc83ddd;
    11'b00111100001: data <= 32'hb5c5b481;
    11'b00111100010: data <= 32'h3d35be2b;
    11'b00111100011: data <= 32'h3e30be32;
    11'b00111100100: data <= 32'h34b8bcd6;
    11'b00111100101: data <= 32'hb556bc4c;
    11'b00111100110: data <= 32'h38d7b82b;
    11'b00111100111: data <= 32'h3d6b3882;
    11'b00111101000: data <= 32'h31ee3b4b;
    11'b00111101001: data <= 32'hbf97b27c;
    11'b00111101010: data <= 32'hc12ebd98;
    11'b00111101011: data <= 32'hbe07bbf7;
    11'b00111101100: data <= 32'hb4b53623;
    11'b00111101101: data <= 32'h2a9b399c;
    11'b00111101110: data <= 32'h324bb431;
    11'b00111101111: data <= 32'h3909b769;
    11'b00111110000: data <= 32'h38bc3caa;
    11'b00111110001: data <= 32'hb53341a2;
    11'b00111110010: data <= 32'hbba74098;
    11'b00111110011: data <= 32'hb32f315d;
    11'b00111110100: data <= 32'h3b9fbcc9;
    11'b00111110101: data <= 32'h3baabb6e;
    11'b00111110110: data <= 32'h3040b567;
    11'b00111110111: data <= 32'h3567b67a;
    11'b00111111000: data <= 32'h3f4fb77f;
    11'b00111111001: data <= 32'h40e32cae;
    11'b00111111010: data <= 32'h39e1366d;
    11'b00111111011: data <= 32'hbebeb481;
    11'b00111111100: data <= 32'hc086bc98;
    11'b00111111101: data <= 32'hbb97bbfa;
    11'b00111111110: data <= 32'h2f3fb55a;
    11'b00111111111: data <= 32'hb047b891;
    11'b01000000000: data <= 32'hb88bbdad;
    11'b01000000001: data <= 32'hb2bfbbcf;
    11'b01000000010: data <= 32'h31d43cd7;
    11'b01000000011: data <= 32'hb4d241d5;
    11'b01000000100: data <= 32'hbc024055;
    11'b01000000101: data <= 32'hbaa72c0e;
    11'b01000000110: data <= 32'hb138ba79;
    11'b01000000111: data <= 32'hac6d27bf;
    11'b01000001000: data <= 32'hb30739ca;
    11'b01000001001: data <= 32'h3981321d;
    11'b01000001010: data <= 32'h40c5b6fa;
    11'b01000001011: data <= 32'h41898ded;
    11'b01000001100: data <= 32'h3b4e3a00;
    11'b01000001101: data <= 32'hbcd3383f;
    11'b01000001110: data <= 32'hbd1fb63c;
    11'b01000001111: data <= 32'h3116bb10;
    11'b01000010000: data <= 32'h39e8bbc8;
    11'b01000010001: data <= 32'hb25bbe05;
    11'b01000010010: data <= 32'hbb4ac03a;
    11'b01000010011: data <= 32'hb3abbd67;
    11'b01000010100: data <= 32'h38f63a36;
    11'b01000010101: data <= 32'h3113403b;
    11'b01000010110: data <= 32'hbc773ce5;
    11'b01000010111: data <= 32'hbeb8b70a;
    11'b01000011000: data <= 32'hbd4cb873;
    11'b01000011001: data <= 32'hbbaf39b1;
    11'b01000011010: data <= 32'hb9223cba;
    11'b01000011011: data <= 32'h36f53022;
    11'b01000011100: data <= 32'h3fb7b94b;
    11'b01000011101: data <= 32'h40553348;
    11'b01000011110: data <= 32'h393b3ea8;
    11'b01000011111: data <= 32'hb9f13efc;
    11'b01000100000: data <= 32'hb4e4380f;
    11'b01000100001: data <= 32'h3befb8a8;
    11'b01000100010: data <= 32'h3be7bc13;
    11'b01000100011: data <= 32'hb4e9bdea;
    11'b01000100100: data <= 32'hb9f6bfbe;
    11'b01000100101: data <= 32'h3863bd8b;
    11'b01000100110: data <= 32'h3ee1307d;
    11'b01000100111: data <= 32'h3b553bd2;
    11'b01000101000: data <= 32'hbc3a31a4;
    11'b01000101001: data <= 32'hc031baec;
    11'b01000101010: data <= 32'hbef4b6fe;
    11'b01000101011: data <= 32'hbcb23a2e;
    11'b01000101100: data <= 32'hbb5639ad;
    11'b01000101101: data <= 32'hb46eb99e;
    11'b01000101110: data <= 32'h3a5abcd1;
    11'b01000101111: data <= 32'h3c7536d5;
    11'b01000110000: data <= 32'h338140e0;
    11'b01000110001: data <= 32'hb7da4117;
    11'b01000110010: data <= 32'h2d4a3c03;
    11'b01000110011: data <= 32'h3b99b2c2;
    11'b01000110100: data <= 32'h3829b62f;
    11'b01000110101: data <= 32'hb8fab825;
    11'b01000110110: data <= 32'hb5e5bc43;
    11'b01000110111: data <= 32'h3e36bc8f;
    11'b01000111000: data <= 32'h418db578;
    11'b01000111001: data <= 32'h3e3733a1;
    11'b01000111010: data <= 32'hba15b2c8;
    11'b01000111011: data <= 32'hbee6ba13;
    11'b01000111100: data <= 32'hbc6cb4d4;
    11'b01000111101: data <= 32'hb8d735b5;
    11'b01000111110: data <= 32'hbb71b535;
    11'b01000111111: data <= 32'hbc16bf4f;
    11'b01001000000: data <= 32'hb40bbf5d;
    11'b01001000001: data <= 32'h36573559;
    11'b01001000010: data <= 32'h2dbe40ec;
    11'b01001000011: data <= 32'hb6ca40b5;
    11'b01001000100: data <= 32'hb31b3a42;
    11'b01001000101: data <= 32'h2db728fc;
    11'b01001000110: data <= 32'hb7833869;
    11'b01001000111: data <= 32'hbc8139d5;
    11'b01001001000: data <= 32'hb271b166;
    11'b01001001001: data <= 32'h4004bb56;
    11'b01001001010: data <= 32'h421cb7f8;
    11'b01001001011: data <= 32'h3ea934a9;
    11'b01001001100: data <= 32'hb5fe353c;
    11'b01001001101: data <= 32'hba0aaaa7;
    11'b01001001110: data <= 32'h3160a539;
    11'b01001001111: data <= 32'h34e7abb0;
    11'b01001010000: data <= 32'hba57bc88;
    11'b01001010001: data <= 32'hbdadc0fd;
    11'b01001010010: data <= 32'hb886c066;
    11'b01001010011: data <= 32'h385bab0e;
    11'b01001010100: data <= 32'h37983ea3;
    11'b01001010101: data <= 32'hb5e43d0d;
    11'b01001010110: data <= 32'hba8c23b4;
    11'b01001010111: data <= 32'hbb5f2d9d;
    11'b01001011000: data <= 32'hbd673d10;
    11'b01001011001: data <= 32'hbe573dd4;
    11'b01001011010: data <= 32'hb7662cb8;
    11'b01001011011: data <= 32'h3e22bc29;
    11'b01001011100: data <= 32'h40a8b6e2;
    11'b01001011101: data <= 32'h3cb13b7a;
    11'b01001011110: data <= 32'haeca3d79;
    11'b01001011111: data <= 32'h33ae3ac0;
    11'b01001100000: data <= 32'h3d0935da;
    11'b01001100001: data <= 32'h3af9a9ad;
    11'b01001100010: data <= 32'hba27bc48;
    11'b01001100011: data <= 32'hbd95c070;
    11'b01001100100: data <= 32'hab8fc016;
    11'b01001100101: data <= 32'h3dc8b823;
    11'b01001100110: data <= 32'h3ceb3811;
    11'b01001100111: data <= 32'hb1f1a7fd;
    11'b01001101000: data <= 32'hbc7fb9df;
    11'b01001101001: data <= 32'hbd202a38;
    11'b01001101010: data <= 32'hbdfb3dcb;
    11'b01001101011: data <= 32'hbee23d17;
    11'b01001101100: data <= 32'hbc21b84a;
    11'b01001101101: data <= 32'h3636be48;
    11'b01001101110: data <= 32'h3c2eb60b;
    11'b01001101111: data <= 32'h36db3e37;
    11'b01001110000: data <= 32'ha8584030;
    11'b01001110001: data <= 32'h39d73d33;
    11'b01001110010: data <= 32'h3e0a393b;
    11'b01001110011: data <= 32'h393437c9;
    11'b01001110100: data <= 32'hbc37ae42;
    11'b01001110101: data <= 32'hbcb6bc8e;
    11'b01001110110: data <= 32'h3a12bdef;
    11'b01001110111: data <= 32'h40d2ba70;
    11'b01001111000: data <= 32'h3f6ab507;
    11'b01001111001: data <= 32'h2d63b9ba;
    11'b01001111010: data <= 32'hba74bb37;
    11'b01001111011: data <= 32'hb90d3020;
    11'b01001111100: data <= 32'hb9f53cc8;
    11'b01001111101: data <= 32'hbdc63736;
    11'b01001111110: data <= 32'hbe51be34;
    11'b01001111111: data <= 32'hb9d0c06c;
    11'b01010000000: data <= 32'h2789b7ec;
    11'b01010000001: data <= 32'ha4af3e59;
    11'b01010000010: data <= 32'haac23f84;
    11'b01010000011: data <= 32'h38ab3b70;
    11'b01010000100: data <= 32'h3b163934;
    11'b01010000101: data <= 32'hb2a73cf4;
    11'b01010000110: data <= 32'hbe4b3cd2;
    11'b01010000111: data <= 32'hbc502ab0;
    11'b01010001000: data <= 32'h3cb7bb7d;
    11'b01010001001: data <= 32'h4152bac0;
    11'b01010001010: data <= 32'h3f66b692;
    11'b01010001011: data <= 32'h3435b6f9;
    11'b01010001100: data <= 32'h926cb5a8;
    11'b01010001101: data <= 32'h398836d4;
    11'b01010001110: data <= 32'h37383b0c;
    11'b01010001111: data <= 32'hbbbfb48a;
    11'b01010010000: data <= 32'hbf54c05e;
    11'b01010010001: data <= 32'hbcb4c0fc;
    11'b01010010010: data <= 32'hae87b9d5;
    11'b01010010011: data <= 32'h318e3b58;
    11'b01010010100: data <= 32'h207239f1;
    11'b01010010101: data <= 32'h2f68aec8;
    11'b01010010110: data <= 32'ha42335cc;
    11'b01010010111: data <= 32'hbc313f28;
    11'b01010011000: data <= 32'hbff8401d;
    11'b01010011001: data <= 32'hbcf438bb;
    11'b01010011010: data <= 32'h3a72baa0;
    11'b01010011011: data <= 32'h3f92ba13;
    11'b01010011100: data <= 32'h3c732db0;
    11'b01010011101: data <= 32'h32a03765;
    11'b01010011110: data <= 32'h3a9337d7;
    11'b01010011111: data <= 32'h3f973a6f;
    11'b01010100000: data <= 32'h3d4e3aca;
    11'b01010100001: data <= 32'hb96db4a2;
    11'b01010100010: data <= 32'hbf0dbf80;
    11'b01010100011: data <= 32'hba8ec03f;
    11'b01010100100: data <= 32'h38fcbb20;
    11'b01010100101: data <= 32'h3adaabfb;
    11'b01010100110: data <= 32'h3287b947;
    11'b01010100111: data <= 32'hb209bcb4;
    11'b01010101000: data <= 32'hb69026aa;
    11'b01010101001: data <= 32'hbcae3f98;
    11'b01010101010: data <= 32'hbfd1400c;
    11'b01010101011: data <= 32'hbe2b3208;
    11'b01010101100: data <= 32'hb1a6bd08;
    11'b01010101101: data <= 32'h3810b9d3;
    11'b01010101110: data <= 32'h29843954;
    11'b01010101111: data <= 32'ha96b3cbf;
    11'b01010110000: data <= 32'h3cdb3b72;
    11'b01010110001: data <= 32'h409a3bb9;
    11'b01010110010: data <= 32'h3d603ca3;
    11'b01010110011: data <= 32'hbaa43847;
    11'b01010110100: data <= 32'hbe41b9a2;
    11'b01010110101: data <= 32'haccebcf9;
    11'b01010110110: data <= 32'h3e37babd;
    11'b01010110111: data <= 32'h3ddeba23;
    11'b01010111000: data <= 32'h3640be00;
    11'b01010111001: data <= 32'ha92dbe74;
    11'b01010111010: data <= 32'h2f1fac2c;
    11'b01010111011: data <= 32'hb57a3e9b;
    11'b01010111100: data <= 32'hbd823d33;
    11'b01010111101: data <= 32'hbf02ba15;
    11'b01010111110: data <= 32'hbca2bf88;
    11'b01010111111: data <= 32'hb951ba64;
    11'b01011000000: data <= 32'hb9a33a8b;
    11'b01011000001: data <= 32'hb4623c4f;
    11'b01011000010: data <= 32'h3c3a3800;
    11'b01011000011: data <= 32'h3f2d398b;
    11'b01011000100: data <= 32'h38ad3e59;
    11'b01011000101: data <= 32'hbd4a3eca;
    11'b01011000110: data <= 32'hbdc93922;
    11'b01011000111: data <= 32'h36b7b5e7;
    11'b01011001000: data <= 32'h3f8cb905;
    11'b01011001001: data <= 32'h3daebaa7;
    11'b01011001010: data <= 32'h356ebd6b;
    11'b01011001011: data <= 32'h3777bccf;
    11'b01011001100: data <= 32'h3d2c31fa;
    11'b01011001101: data <= 32'h3c033d5a;
    11'b01011001110: data <= 32'hb879383e;
    11'b01011001111: data <= 32'hbeddbdd2;
    11'b01011010000: data <= 32'hbe37c047;
    11'b01011010001: data <= 32'hbb95bac5;
    11'b01011010010: data <= 32'hb98c36a0;
    11'b01011010011: data <= 32'hb49c2ce0;
    11'b01011010100: data <= 32'h38ceb967;
    11'b01011010101: data <= 32'h3b242b92;
    11'b01011010110: data <= 32'hb4b53f4d;
    11'b01011010111: data <= 32'hbeee40f4;
    11'b01011011000: data <= 32'hbdd93d63;
    11'b01011011001: data <= 32'h3461a89a;
    11'b01011011010: data <= 32'h3cfcb6d9;
    11'b01011011011: data <= 32'h3875b580;
    11'b01011011100: data <= 32'haac8b7dc;
    11'b01011011101: data <= 32'h3bbeb593;
    11'b01011011110: data <= 32'h40d33887;
    11'b01011011111: data <= 32'h401c3cd2;
    11'b01011100000: data <= 32'h98af355f;
    11'b01011100001: data <= 32'hbdf4bd11;
    11'b01011100010: data <= 32'hbccebea8;
    11'b01011100011: data <= 32'hb49bb988;
    11'b01011100100: data <= 32'ha86db3e1;
    11'b01011100101: data <= 32'hadd0bcee;
    11'b01011100110: data <= 32'h3370bfba;
    11'b01011100111: data <= 32'h3594b8a5;
    11'b01011101000: data <= 32'hb83e3ef0;
    11'b01011101001: data <= 32'hbe7740de;
    11'b01011101010: data <= 32'hbdec3c26;
    11'b01011101011: data <= 32'hb662b669;
    11'b01011101100: data <= 32'ha929b62b;
    11'b01011101101: data <= 32'hb99f3450;
    11'b01011101110: data <= 32'hb9123585;
    11'b01011101111: data <= 32'h3c7f3253;
    11'b01011110000: data <= 32'h4197396c;
    11'b01011110001: data <= 32'h40633d14;
    11'b01011110010: data <= 32'ha96f3af3;
    11'b01011110011: data <= 32'hbd03b258;
    11'b01011110100: data <= 32'hb6ffb8c6;
    11'b01011110101: data <= 32'h39beb4af;
    11'b01011110110: data <= 32'h3955b97e;
    11'b01011110111: data <= 32'h2ca5c016;
    11'b01011111000: data <= 32'h31b3c109;
    11'b01011111001: data <= 32'h38d3baa8;
    11'b01011111010: data <= 32'h32063dae;
    11'b01011111011: data <= 32'hbaea3ecb;
    11'b01011111100: data <= 32'hbd572a01;
    11'b01011111101: data <= 32'hbc62bc62;
    11'b01011111110: data <= 32'hbcb5b739;
    11'b01011111111: data <= 32'hbe8438a8;
    11'b01100000000: data <= 32'hbc4e3797;
    11'b01100000001: data <= 32'h3ae9af8d;
    11'b01100000010: data <= 32'h40903413;
    11'b01100000011: data <= 32'h3db53d68;
    11'b01100000100: data <= 32'hb8a03ef1;
    11'b01100000101: data <= 32'hbc8e3c6b;
    11'b01100000110: data <= 32'h31d637ac;
    11'b01100000111: data <= 32'h3d0b31cc;
    11'b01100001000: data <= 32'h39ebb8e2;
    11'b01100001001: data <= 32'hae69bf94;
    11'b01100001010: data <= 32'h35cfc046;
    11'b01100001011: data <= 32'h3df4b893;
    11'b01100001100: data <= 32'h3ded3c6f;
    11'b01100001101: data <= 32'h316b3aab;
    11'b01100001110: data <= 32'hbbfdbaa3;
    11'b01100001111: data <= 32'hbd41bde5;
    11'b01100010000: data <= 32'hbdd5b686;
    11'b01100010001: data <= 32'hbec23782;
    11'b01100010010: data <= 32'hbc82b396;
    11'b01100010011: data <= 32'h365abcee;
    11'b01100010100: data <= 32'h3d3cb8c9;
    11'b01100010101: data <= 32'h364d3d0b;
    11'b01100010110: data <= 32'hbc71409c;
    11'b01100010111: data <= 32'hbc603f3c;
    11'b01100011000: data <= 32'h34b43b6b;
    11'b01100011001: data <= 32'h3b323786;
    11'b01100011010: data <= 32'haaafadcd;
    11'b01100011011: data <= 32'hb9a2bbd6;
    11'b01100011100: data <= 32'h382abca5;
    11'b01100011101: data <= 32'h40bfacea;
    11'b01100011110: data <= 32'h41113b87;
    11'b01100011111: data <= 32'h3b0c36a1;
    11'b01100100000: data <= 32'hb901bb44;
    11'b01100100001: data <= 32'hbb32bc56;
    11'b01100100010: data <= 32'hba1cab66;
    11'b01100100011: data <= 32'hbb9130f1;
    11'b01100100100: data <= 32'hbaa7bd30;
    11'b01100100101: data <= 32'h22e1c0f9;
    11'b01100100110: data <= 32'h3896bdb4;
    11'b01100100111: data <= 32'hae3d3bc5;
    11'b01100101000: data <= 32'hbc624056;
    11'b01100101001: data <= 32'hbb8a3de9;
    11'b01100101010: data <= 32'ha939382c;
    11'b01100101011: data <= 32'hb029371f;
    11'b01100101100: data <= 32'hbd3d383c;
    11'b01100101101: data <= 32'hbe0024a0;
    11'b01100101110: data <= 32'h36eab601;
    11'b01100101111: data <= 32'h414430f2;
    11'b01100110000: data <= 32'h41533aef;
    11'b01100110001: data <= 32'h3ac73900;
    11'b01100110010: data <= 32'hb6a9aeb6;
    11'b01100110011: data <= 32'hb000a69d;
    11'b01100110100: data <= 32'h36033894;
    11'b01100110101: data <= 32'ha67c9ca6;
    11'b01100110110: data <= 32'hb84abfd5;
    11'b01100110111: data <= 32'hb0abc229;
    11'b01100111000: data <= 32'h3837beee;
    11'b01100111001: data <= 32'h359d3913;
    11'b01100111010: data <= 32'hb5e53da2;
    11'b01100111011: data <= 32'hb87b3609;
    11'b01100111100: data <= 32'hb6dfb5da;
    11'b01100111101: data <= 32'hbc6233d4;
    11'b01100111110: data <= 32'hc0823b56;
    11'b01100111111: data <= 32'hc01836c0;
    11'b01101000000: data <= 32'h2e42b6ad;
    11'b01101000001: data <= 32'h4027b321;
    11'b01101000010: data <= 32'h3f3c39c5;
    11'b01101000011: data <= 32'h30db3caa;
    11'b01101000100: data <= 32'hb6d73c08;
    11'b01101000101: data <= 32'h38613c53;
    11'b01101000110: data <= 32'h3cac3ccc;
    11'b01101000111: data <= 32'h35253258;
    11'b01101001000: data <= 32'hb91abeff;
    11'b01101001001: data <= 32'hb15bc145;
    11'b01101001010: data <= 32'h3c54bd69;
    11'b01101001011: data <= 32'h3dbf36de;
    11'b01101001100: data <= 32'h399c3806;
    11'b01101001101: data <= 32'ha7dfb9ce;
    11'b01101001110: data <= 32'hb785bc0f;
    11'b01101001111: data <= 32'hbd313230;
    11'b01101010000: data <= 32'hc08f3bdf;
    11'b01101010001: data <= 32'hc00d28aa;
    11'b01101010010: data <= 32'hb4adbd3c;
    11'b01101010011: data <= 32'h3c47bc6d;
    11'b01101010100: data <= 32'h3891368e;
    11'b01101010101: data <= 32'hb9283e0f;
    11'b01101010110: data <= 32'hb7f73e75;
    11'b01101010111: data <= 32'h3a7d3e16;
    11'b01101011000: data <= 32'h3c7e3de4;
    11'b01101011001: data <= 32'hb3763972;
    11'b01101011010: data <= 32'hbd0aba66;
    11'b01101011011: data <= 32'hb3cfbde9;
    11'b01101011100: data <= 32'h3edbb8db;
    11'b01101011101: data <= 32'h40bf363d;
    11'b01101011110: data <= 32'h3dbaa97e;
    11'b01101011111: data <= 32'h362ebc72;
    11'b01101100000: data <= 32'ha9d7bb04;
    11'b01101100001: data <= 32'hb8853856;
    11'b01101100010: data <= 32'hbd8a3b3b;
    11'b01101100011: data <= 32'hbe04b9f8;
    11'b01101100100: data <= 32'hb857c0dd;
    11'b01101100101: data <= 32'h3357bfe5;
    11'b01101100110: data <= 32'hb2f9258a;
    11'b01101100111: data <= 32'hbb303d46;
    11'b01101101000: data <= 32'hb5f43cf2;
    11'b01101101001: data <= 32'h39a13bfd;
    11'b01101101010: data <= 32'h36323d08;
    11'b01101101011: data <= 32'hbd5f3cb3;
    11'b01101101100: data <= 32'hc0373489;
    11'b01101101101: data <= 32'hb7a3b685;
    11'b01101101110: data <= 32'h3f75ae03;
    11'b01101101111: data <= 32'h40e435ee;
    11'b01101110000: data <= 32'h3d42a9cd;
    11'b01101110001: data <= 32'h3741b8e6;
    11'b01101110010: data <= 32'h38fc242d;
    11'b01101110011: data <= 32'h392e3ced;
    11'b01101110100: data <= 32'hb24a3b69;
    11'b01101110101: data <= 32'hbb5bbd09;
    11'b01101110110: data <= 32'hb8f2c1ec;
    11'b01101110111: data <= 32'ha16dc078;
    11'b01101111000: data <= 32'had4fb349;
    11'b01101111001: data <= 32'hb5ba3910;
    11'b01101111010: data <= 32'h2c2d2c7e;
    11'b01101111011: data <= 32'h382fb04e;
    11'b01101111100: data <= 32'hb6563a2b;
    11'b01101111101: data <= 32'hc0703dd3;
    11'b01101111110: data <= 32'hc14b3ae1;
    11'b01101111111: data <= 32'hba3eb028;
    11'b01110000000: data <= 32'h3d62b41c;
    11'b01110000001: data <= 32'h3e1e31f2;
    11'b01110000010: data <= 32'h366a345c;
    11'b01110000011: data <= 32'h317c349a;
    11'b01110000100: data <= 32'h3cb73c30;
    11'b01110000101: data <= 32'h3e5f3f89;
    11'b01110000110: data <= 32'h378d3c9e;
    11'b01110000111: data <= 32'hba3bbc32;
    11'b01110001000: data <= 32'hb93bc0ea;
    11'b01110001001: data <= 32'h3511bead;
    11'b01110001010: data <= 32'h3a1bb20d;
    11'b01110001011: data <= 32'h38fab0ff;
    11'b01110001100: data <= 32'h392fbcaf;
    11'b01110001101: data <= 32'h387dbc6b;
    11'b01110001110: data <= 32'hb87b3742;
    11'b01110001111: data <= 32'hc0623e09;
    11'b01110010000: data <= 32'hc0f63995;
    11'b01110010001: data <= 32'hbbb7ba12;
    11'b01110010010: data <= 32'h3722bc20;
    11'b01110010011: data <= 32'h313db23c;
    11'b01110010100: data <= 32'hb9b137ef;
    11'b01110010101: data <= 32'hb1dc3a8c;
    11'b01110010110: data <= 32'h3d9a3dc5;
    11'b01110010111: data <= 32'h3f0e401d;
    11'b01110011000: data <= 32'h32653de9;
    11'b01110011001: data <= 32'hbd11b216;
    11'b01110011010: data <= 32'hba6abcbb;
    11'b01110011011: data <= 32'h3a4cb8f0;
    11'b01110011100: data <= 32'h3e5b2c37;
    11'b01110011101: data <= 32'h3d3fb91a;
    11'b01110011110: data <= 32'h3c0dbf0e;
    11'b01110011111: data <= 32'h3b0dbd12;
    11'b01110100000: data <= 32'h2ebe391c;
    11'b01110100001: data <= 32'hbcc53df7;
    11'b01110100010: data <= 32'hbeb12e5d;
    11'b01110100011: data <= 32'hbb5dbef5;
    11'b01110100100: data <= 32'hb507bf6f;
    11'b01110100101: data <= 32'hba98b898;
    11'b01110100110: data <= 32'hbd24358c;
    11'b01110100111: data <= 32'hb40e37b5;
    11'b01110101000: data <= 32'h3d5c3aa7;
    11'b01110101001: data <= 32'h3ce83e5c;
    11'b01110101010: data <= 32'hb9eb3ec5;
    11'b01110101011: data <= 32'hc0233a6d;
    11'b01110101100: data <= 32'hbc3e2d18;
    11'b01110101101: data <= 32'h3b753371;
    11'b01110101110: data <= 32'h3eb2346a;
    11'b01110101111: data <= 32'h3c80b954;
    11'b01110110000: data <= 32'h3af5bde6;
    11'b01110110001: data <= 32'h3d32b896;
    11'b01110110010: data <= 32'h3ce83d14;
    11'b01110110011: data <= 32'h31a93e41;
    11'b01110110100: data <= 32'hb9efb5c8;
    11'b01110110101: data <= 32'hb9e4c081;
    11'b01110110110: data <= 32'hb874c021;
    11'b01110110111: data <= 32'hbb44b949;
    11'b01110111000: data <= 32'hbbccb017;
    11'b01110111001: data <= 32'h2ebdb8cf;
    11'b01110111010: data <= 32'h3ce5b787;
    11'b01110111011: data <= 32'h38453a10;
    11'b01110111100: data <= 32'hbe4c3ec4;
    11'b01110111101: data <= 32'hc1233d70;
    11'b01110111110: data <= 32'hbd0038a7;
    11'b01110111111: data <= 32'h38a23558;
    11'b01111000000: data <= 32'h3a9e3261;
    11'b01111000001: data <= 32'h2b65b6b1;
    11'b01111000010: data <= 32'h3417b995;
    11'b01111000011: data <= 32'h3e413642;
    11'b01111000100: data <= 32'h40453f97;
    11'b01111000101: data <= 32'h3c4b3ee8;
    11'b01111000110: data <= 32'hb4dab453;
    11'b01111000111: data <= 32'hb904bf38;
    11'b01111001000: data <= 32'hb4b3bd75;
    11'b01111001001: data <= 32'hb2d5b509;
    11'b01111001010: data <= 32'hadc1b90c;
    11'b01111001011: data <= 32'h395ebf2d;
    11'b01111001100: data <= 32'h3cf6bead;
    11'b01111001101: data <= 32'h34c02f4f;
    11'b01111001110: data <= 32'hbe5c3e3d;
    11'b01111001111: data <= 32'hc0953cfe;
    11'b01111010000: data <= 32'hbca5301e;
    11'b01111010001: data <= 32'haa98b4fc;
    11'b01111010010: data <= 32'hb7c6b11c;
    11'b01111010011: data <= 32'hbd21b2ab;
    11'b01111010100: data <= 32'hb723b076;
    11'b01111010101: data <= 32'h3e453a89;
    11'b01111010110: data <= 32'h40ad3ff5;
    11'b01111010111: data <= 32'h3bfa3f47;
    11'b01111011000: data <= 32'hb8fc3580;
    11'b01111011001: data <= 32'hb9e5b8ac;
    11'b01111011010: data <= 32'h3071adc8;
    11'b01111011011: data <= 32'h38c834cc;
    11'b01111011100: data <= 32'h38ebbaf2;
    11'b01111011101: data <= 32'h3bdcc0d0;
    11'b01111011110: data <= 32'h3d85c018;
    11'b01111011111: data <= 32'h39fe2dd4;
    11'b01111100000: data <= 32'hb9283dea;
    11'b01111100001: data <= 32'hbd19399b;
    11'b01111100010: data <= 32'hba0dba68;
    11'b01111100011: data <= 32'hb865bc88;
    11'b01111100100: data <= 32'hbdefb814;
    11'b01111100101: data <= 32'hc02db350;
    11'b01111100110: data <= 32'hba20b4cb;
    11'b01111100111: data <= 32'h3da43428;
    11'b01111101000: data <= 32'h3f6d3d56;
    11'b01111101001: data <= 32'h30863ebd;
    11'b01111101010: data <= 32'hbd953c45;
    11'b01111101011: data <= 32'hbbda3972;
    11'b01111101100: data <= 32'h35dc3c0a;
    11'b01111101101: data <= 32'h3a8f3a65;
    11'b01111101110: data <= 32'h37b4ba21;
    11'b01111101111: data <= 32'h3974c058;
    11'b01111110000: data <= 32'h3de7bdde;
    11'b01111110001: data <= 32'h3e6a394d;
    11'b01111110010: data <= 32'h39c23e2a;
    11'b01111110011: data <= 32'had333240;
    11'b01111110100: data <= 32'hb3e2bda7;
    11'b01111110101: data <= 32'hb905bd90;
    11'b01111110110: data <= 32'hbe7cb792;
    11'b01111110111: data <= 32'hbfb5b6b5;
    11'b01111111000: data <= 32'hb805bc83;
    11'b01111111001: data <= 32'h3d1dbc1e;
    11'b01111111010: data <= 32'h3c98339e;
    11'b01111111011: data <= 32'hba113d54;
    11'b01111111100: data <= 32'hbfc63db6;
    11'b01111111101: data <= 32'hbc533cef;
    11'b01111111110: data <= 32'h34103d2e;
    11'b01111111111: data <= 32'h32a23ae7;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    