
module memory_rom_48(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3d4d3ae2;
    11'b00000000001: data <= 32'h3a783727;
    11'b00000000010: data <= 32'hb9f0b814;
    11'b00000000011: data <= 32'hbbb9be6a;
    11'b00000000100: data <= 32'h3a16be2e;
    11'b00000000101: data <= 32'h40a1b610;
    11'b00000000110: data <= 32'h3f6f3328;
    11'b00000000111: data <= 32'h32afb800;
    11'b00000001000: data <= 32'hba4fbc62;
    11'b00000001001: data <= 32'hbb59b326;
    11'b00000001010: data <= 32'hbcb83bc7;
    11'b00000001011: data <= 32'hbe623715;
    11'b00000001100: data <= 32'hbce2bdd4;
    11'b00000001101: data <= 32'hb04bc057;
    11'b00000001110: data <= 32'h3568b858;
    11'b00000001111: data <= 32'hb2d23e52;
    11'b00000010000: data <= 32'hb7d64024;
    11'b00000010001: data <= 32'h34e73d16;
    11'b00000010010: data <= 32'h3b363aa9;
    11'b00000010011: data <= 32'hac543be2;
    11'b00000010100: data <= 32'hbe08391b;
    11'b00000010101: data <= 32'hbc6eb596;
    11'b00000010110: data <= 32'h3cc1ba84;
    11'b00000010111: data <= 32'h41a4b59a;
    11'b00000011000: data <= 32'h4039a568;
    11'b00000011001: data <= 32'h3688b6e4;
    11'b00000011010: data <= 32'hb210b89e;
    11'b00000011011: data <= 32'h3295349d;
    11'b00000011100: data <= 32'h26eb3b51;
    11'b00000011101: data <= 32'hbb90b412;
    11'b00000011110: data <= 32'hbd72c0a4;
    11'b00000011111: data <= 32'hb978c176;
    11'b00000100000: data <= 32'h9b11babc;
    11'b00000100001: data <= 32'hae193c68;
    11'b00000100010: data <= 32'hb4133cac;
    11'b00000100011: data <= 32'h2e7b3474;
    11'b00000100100: data <= 32'h2d36362b;
    11'b00000100101: data <= 32'hbc6c3d8b;
    11'b00000100110: data <= 32'hc0703e26;
    11'b00000100111: data <= 32'hbd80362d;
    11'b00000101000: data <= 32'h3bdbb8c1;
    11'b00000101001: data <= 32'h409fb646;
    11'b00000101010: data <= 32'h3ddf3305;
    11'b00000101011: data <= 32'h32f8357f;
    11'b00000101100: data <= 32'h374236c2;
    11'b00000101101: data <= 32'h3d9d3bb1;
    11'b00000101110: data <= 32'h3c4b3c20;
    11'b00000101111: data <= 32'hb81bb657;
    11'b00000110000: data <= 32'hbd79c093;
    11'b00000110001: data <= 32'hb891c102;
    11'b00000110010: data <= 32'h3880bb31;
    11'b00000110011: data <= 32'h3994352d;
    11'b00000110100: data <= 32'h3357b17a;
    11'b00000110101: data <= 32'ha3c4bb6f;
    11'b00000110110: data <= 32'hb68caf3c;
    11'b00000110111: data <= 32'hbe073e15;
    11'b00000111000: data <= 32'hc0bd3ee3;
    11'b00000111001: data <= 32'hbe713162;
    11'b00000111010: data <= 32'h32ecbc57;
    11'b00000111011: data <= 32'h3c2bb90d;
    11'b00000111100: data <= 32'h34cd389c;
    11'b00000111101: data <= 32'hb2973c7a;
    11'b00000111110: data <= 32'h3a933c8b;
    11'b00000111111: data <= 32'h3ff53d65;
    11'b00001000000: data <= 32'h3d2a3d42;
    11'b00001000001: data <= 32'hb96c329d;
    11'b00001000010: data <= 32'hbda7bd20;
    11'b00001000011: data <= 32'hac7cbe48;
    11'b00001000100: data <= 32'h3dfcb95f;
    11'b00001000101: data <= 32'h3e3fb4f4;
    11'b00001000110: data <= 32'h3962bc9b;
    11'b00001000111: data <= 32'h30d0be4b;
    11'b00001001000: data <= 32'hae90b388;
    11'b00001001001: data <= 32'hbb1b3def;
    11'b00001001010: data <= 32'hbf273d04;
    11'b00001001011: data <= 32'hbe94b9e7;
    11'b00001001100: data <= 32'hb92fbfbd;
    11'b00001001101: data <= 32'hb31abbd9;
    11'b00001001110: data <= 32'hb9343951;
    11'b00001001111: data <= 32'hb8143cd3;
    11'b00001010000: data <= 32'h3ab03b95;
    11'b00001010001: data <= 32'h3efa3c80;
    11'b00001010010: data <= 32'h38f13e53;
    11'b00001010011: data <= 32'hbd723cd7;
    11'b00001010100: data <= 32'hbe572e83;
    11'b00001010101: data <= 32'h3510b80f;
    11'b00001010110: data <= 32'h3ffeb58f;
    11'b00001010111: data <= 32'h3f1eb800;
    11'b00001011000: data <= 32'h39c4bd0e;
    11'b00001011001: data <= 32'h3829bd26;
    11'b00001011010: data <= 32'h3b1d3164;
    11'b00001011011: data <= 32'h36fb3ddb;
    11'b00001011100: data <= 32'hba743914;
    11'b00001011101: data <= 32'hbddfbe43;
    11'b00001011110: data <= 32'hbc79c0ef;
    11'b00001011111: data <= 32'hb9f7bcb1;
    11'b00001100000: data <= 32'hba6035e0;
    11'b00001100001: data <= 32'hb6a636ae;
    11'b00001100010: data <= 32'h3956b0d5;
    11'b00001100011: data <= 32'h3c2035c9;
    11'b00001100100: data <= 32'hb5ab3ea0;
    11'b00001100101: data <= 32'hc0194005;
    11'b00001100110: data <= 32'hbf273c13;
    11'b00001100111: data <= 32'h33b4203c;
    11'b00001101000: data <= 32'h3e53b2b1;
    11'b00001101001: data <= 32'h3c2db48b;
    11'b00001101010: data <= 32'h33a2b8fa;
    11'b00001101011: data <= 32'h3ac4b626;
    11'b00001101100: data <= 32'h3fe73a8b;
    11'b00001101101: data <= 32'h3ea63e38;
    11'b00001101110: data <= 32'haac33691;
    11'b00001101111: data <= 32'hbd04be69;
    11'b00001110000: data <= 32'hbc0ac055;
    11'b00001110001: data <= 32'hb552bbc5;
    11'b00001110010: data <= 32'hb065af3a;
    11'b00001110011: data <= 32'h285cba79;
    11'b00001110100: data <= 32'h3871be23;
    11'b00001110101: data <= 32'h3808b7a5;
    11'b00001110110: data <= 32'hba763e23;
    11'b00001110111: data <= 32'hc04a405b;
    11'b00001111000: data <= 32'hbf393bc1;
    11'b00001111001: data <= 32'hb413b4f7;
    11'b00001111010: data <= 32'h36c1b644;
    11'b00001111011: data <= 32'hb4b52a59;
    11'b00001111100: data <= 32'hb84a30c5;
    11'b00001111101: data <= 32'h3b7035be;
    11'b00001111110: data <= 32'h410d3cb2;
    11'b00001111111: data <= 32'h401f3eac;
    11'b00010000000: data <= 32'h9d313a3a;
    11'b00010000001: data <= 32'hbcd6b99e;
    11'b00010000010: data <= 32'hb851bc4a;
    11'b00010000011: data <= 32'h387bb64b;
    11'b00010000100: data <= 32'h39d9b71c;
    11'b00010000101: data <= 32'h376abef4;
    11'b00010000110: data <= 32'h38cbc0bf;
    11'b00010000111: data <= 32'h38edbad2;
    11'b00010001000: data <= 32'hb49d3d7c;
    11'b00010001001: data <= 32'hbdb13ef2;
    11'b00010001010: data <= 32'hbe033051;
    11'b00010001011: data <= 32'hba7cbc8a;
    11'b00010001100: data <= 32'hba40b9df;
    11'b00010001101: data <= 32'hbdce32e4;
    11'b00010001110: data <= 32'hbc863633;
    11'b00010001111: data <= 32'h3a3a3437;
    11'b00010010000: data <= 32'h40993aae;
    11'b00010010001: data <= 32'h3df33e7e;
    11'b00010010010: data <= 32'hb9083dea;
    11'b00010010011: data <= 32'hbd7c38e5;
    11'b00010010100: data <= 32'haf0a3294;
    11'b00010010101: data <= 32'h3cb03419;
    11'b00010010110: data <= 32'h3c21b6e8;
    11'b00010010111: data <= 32'h36cfbf72;
    11'b00010011000: data <= 32'h3992c06e;
    11'b00010011001: data <= 32'h3d47b85f;
    11'b00010011010: data <= 32'h3bb13d50;
    11'b00010011011: data <= 32'hb33e3c65;
    11'b00010011100: data <= 32'hbbceba23;
    11'b00010011101: data <= 32'hbc2cbef5;
    11'b00010011110: data <= 32'hbd3abaf3;
    11'b00010011111: data <= 32'hbf0730b0;
    11'b00010100000: data <= 32'hbcb8b063;
    11'b00010100001: data <= 32'h3883ba0d;
    11'b00010100010: data <= 32'h3e57b04d;
    11'b00010100011: data <= 32'h379b3d59;
    11'b00010100100: data <= 32'hbd804007;
    11'b00010100101: data <= 32'hbe2b3e16;
    11'b00010100110: data <= 32'h91f43b46;
    11'b00010100111: data <= 32'h3bef38b4;
    11'b00010101000: data <= 32'h3613b07b;
    11'b00010101001: data <= 32'hb3d6bceb;
    11'b00010101010: data <= 32'h394fbd3a;
    11'b00010101011: data <= 32'h4041308e;
    11'b00010101100: data <= 32'h40583d9e;
    11'b00010101101: data <= 32'h39ec39d8;
    11'b00010101110: data <= 32'hb825bc0b;
    11'b00010101111: data <= 32'hba97be18;
    11'b00010110000: data <= 32'hbb47b807;
    11'b00010110001: data <= 32'hbc842000;
    11'b00010110010: data <= 32'hb9c0bc53;
    11'b00010110011: data <= 32'h372ac03c;
    11'b00010110100: data <= 32'h3b9abcd1;
    11'b00010110101: data <= 32'hb1083b6b;
    11'b00010110110: data <= 32'hbe414010;
    11'b00010110111: data <= 32'hbdb43df6;
    11'b00010111000: data <= 32'hb1c9394e;
    11'b00010111001: data <= 32'h2f0536ee;
    11'b00010111010: data <= 32'hbb743267;
    11'b00010111011: data <= 32'hbd0bb61f;
    11'b00010111100: data <= 32'h36d2b69d;
    11'b00010111101: data <= 32'h40fc38c3;
    11'b00010111110: data <= 32'h412d3dac;
    11'b00010111111: data <= 32'h3b353a86;
    11'b00011000000: data <= 32'hb65db611;
    11'b00011000001: data <= 32'hb54eb772;
    11'b00011000010: data <= 32'h28363514;
    11'b00011000011: data <= 32'hb094251b;
    11'b00011000100: data <= 32'hb232bf36;
    11'b00011000101: data <= 32'h36cfc1f4;
    11'b00011000110: data <= 32'h3a87beee;
    11'b00011000111: data <= 32'h2ea83918;
    11'b00011001000: data <= 32'hbb1c3e2f;
    11'b00011001001: data <= 32'hbb1d3901;
    11'b00011001010: data <= 32'hb61fb3cb;
    11'b00011001011: data <= 32'hbaf01e2a;
    11'b00011001100: data <= 32'hc03a367b;
    11'b00011001101: data <= 32'hc0172c18;
    11'b00011001110: data <= 32'h2e2cb43b;
    11'b00011001111: data <= 32'h4063351f;
    11'b00011010000: data <= 32'h40003ca5;
    11'b00011010001: data <= 32'h33783ca6;
    11'b00011010010: data <= 32'hb8fb3990;
    11'b00011010011: data <= 32'h2fbd3ab6;
    11'b00011010100: data <= 32'h3a8a3cc3;
    11'b00011010101: data <= 32'h362d342a;
    11'b00011010110: data <= 32'hb0cdbf4c;
    11'b00011010111: data <= 32'h3579c1a3;
    11'b00011011000: data <= 32'h3cb8bdb3;
    11'b00011011001: data <= 32'h3c6c38ff;
    11'b00011011010: data <= 32'h354a3b1f;
    11'b00011011011: data <= 32'haf3eb6b3;
    11'b00011011100: data <= 32'hb581bc39;
    11'b00011011101: data <= 32'hbd10b32e;
    11'b00011011110: data <= 32'hc0de37b6;
    11'b00011011111: data <= 32'hc048b099;
    11'b00011100000: data <= 32'hb00ebc20;
    11'b00011100001: data <= 32'h3dd5b949;
    11'b00011100010: data <= 32'h3af938ea;
    11'b00011100011: data <= 32'hb9963d93;
    11'b00011100100: data <= 32'hbb2d3dd1;
    11'b00011100101: data <= 32'h357d3e4d;
    11'b00011100110: data <= 32'h3b6b3e7c;
    11'b00011100111: data <= 32'ha32938df;
    11'b00011101000: data <= 32'hba86bca4;
    11'b00011101001: data <= 32'h2a94bf46;
    11'b00011101010: data <= 32'h3ea5b89e;
    11'b00011101011: data <= 32'h404a3a74;
    11'b00011101100: data <= 32'h3d6036fb;
    11'b00011101101: data <= 32'h37e8bb6a;
    11'b00011101110: data <= 32'ha35bbc5f;
    11'b00011101111: data <= 32'hba922f64;
    11'b00011110000: data <= 32'hbef838b1;
    11'b00011110001: data <= 32'hbe3aba06;
    11'b00011110010: data <= 32'hb0b0c069;
    11'b00011110011: data <= 32'h3a14bf26;
    11'b00011110100: data <= 32'h8340211f;
    11'b00011110101: data <= 32'hbc8e3cfd;
    11'b00011110110: data <= 32'hbaa33d6d;
    11'b00011110111: data <= 32'h36263d2c;
    11'b00011111000: data <= 32'h36113d8d;
    11'b00011111001: data <= 32'hbc803afb;
    11'b00011111010: data <= 32'hbf8fb43f;
    11'b00011111011: data <= 32'hb6a1b9b0;
    11'b00011111100: data <= 32'h3f452ff3;
    11'b00011111101: data <= 32'h40f43b23;
    11'b00011111110: data <= 32'h3dfd353a;
    11'b00011111111: data <= 32'h38b7b8fb;
    11'b00100000000: data <= 32'h36f7b3d9;
    11'b00100000001: data <= 32'h31303bec;
    11'b00100000010: data <= 32'hb88d3acb;
    11'b00100000011: data <= 32'hba56bce9;
    11'b00100000100: data <= 32'hacd2c1ed;
    11'b00100000101: data <= 32'h375fc0aa;
    11'b00100000110: data <= 32'hab4bb4fe;
    11'b00100000111: data <= 32'hb9803a16;
    11'b00100001000: data <= 32'hb4033736;
    11'b00100001001: data <= 32'h37193350;
    11'b00100001010: data <= 32'hb53039ee;
    11'b00100001011: data <= 32'hc0623bc6;
    11'b00100001100: data <= 32'hc1703513;
    11'b00100001101: data <= 32'hbaa6b41a;
    11'b00100001110: data <= 32'h3de22db7;
    11'b00100001111: data <= 32'h3f5c38ec;
    11'b00100010000: data <= 32'h399e369b;
    11'b00100010001: data <= 32'h319c3114;
    11'b00100010010: data <= 32'h3a413b74;
    11'b00100010011: data <= 32'h3c3b3fba;
    11'b00100010100: data <= 32'h34023ce9;
    11'b00100010101: data <= 32'hb7e8bc9f;
    11'b00100010110: data <= 32'hb0d2c180;
    11'b00100010111: data <= 32'h389abfbb;
    11'b00100011000: data <= 32'h3918b198;
    11'b00100011001: data <= 32'h363b3259;
    11'b00100011010: data <= 32'h38dcb981;
    11'b00100011011: data <= 32'h3954bada;
    11'b00100011100: data <= 32'hb8b133ea;
    11'b00100011101: data <= 32'hc0e83c0b;
    11'b00100011110: data <= 32'hc184356a;
    11'b00100011111: data <= 32'hbba1b9a9;
    11'b00100100000: data <= 32'h3a71b9d8;
    11'b00100100001: data <= 32'h3905a490;
    11'b00100100010: data <= 32'hb7bb36ca;
    11'b00100100011: data <= 32'hb5d239f0;
    11'b00100100100: data <= 32'h3b863e6d;
    11'b00100100101: data <= 32'h3d7e40b1;
    11'b00100100110: data <= 32'h31703e1f;
    11'b00100100111: data <= 32'hbbcfb842;
    11'b00100101000: data <= 32'hb825beb2;
    11'b00100101001: data <= 32'h3a84bad4;
    11'b00100101010: data <= 32'h3dde343c;
    11'b00100101011: data <= 32'h3d58b196;
    11'b00100101100: data <= 32'h3cf4bd86;
    11'b00100101101: data <= 32'h3c09bcdb;
    11'b00100101110: data <= 32'hb0b73617;
    11'b00100101111: data <= 32'hbec73cb1;
    11'b00100110000: data <= 32'hbfe4a511;
    11'b00100110001: data <= 32'hb9ddbe95;
    11'b00100110010: data <= 32'h3247bf1f;
    11'b00100110011: data <= 32'hb695b970;
    11'b00100110100: data <= 32'hbcf9329d;
    11'b00100110101: data <= 32'hb83538e4;
    11'b00100110110: data <= 32'h3c0f3d0e;
    11'b00100110111: data <= 32'h3c4e3fcd;
    11'b00100111000: data <= 32'hb9783e56;
    11'b00100111001: data <= 32'hbfd8345f;
    11'b00100111010: data <= 32'hbc42b6a2;
    11'b00100111011: data <= 32'h3ac93151;
    11'b00100111100: data <= 32'h3ee838cf;
    11'b00100111101: data <= 32'h3dbeb4a7;
    11'b00100111110: data <= 32'h3cdfbd49;
    11'b00100111111: data <= 32'h3d2bb922;
    11'b00101000000: data <= 32'h3a0d3c99;
    11'b00101000001: data <= 32'hb6223e1d;
    11'b00101000010: data <= 32'hbb2eb54a;
    11'b00101000011: data <= 32'hb64bc097;
    11'b00101000100: data <= 32'had57c08f;
    11'b00101000101: data <= 32'hb9a4bb78;
    11'b00101000110: data <= 32'hbc59b14f;
    11'b00101000111: data <= 32'hacdfb382;
    11'b00101001000: data <= 32'h3cad2cee;
    11'b00101001001: data <= 32'h38883c0a;
    11'b00101001010: data <= 32'hbe743da2;
    11'b00101001011: data <= 32'hc17f3a81;
    11'b00101001100: data <= 32'hbdd63447;
    11'b00101001101: data <= 32'h3879371c;
    11'b00101001110: data <= 32'h3c7f37b8;
    11'b00101001111: data <= 32'h3845b4a9;
    11'b00101010000: data <= 32'h384fba0b;
    11'b00101010001: data <= 32'h3d7b35f0;
    11'b00101010010: data <= 32'h3e60401a;
    11'b00101010011: data <= 32'h39373fb6;
    11'b00101010100: data <= 32'hb452b434;
    11'b00101010101: data <= 32'hb470c02d;
    11'b00101010110: data <= 32'ha8ecbf26;
    11'b00101010111: data <= 32'hb3c0b88b;
    11'b00101011000: data <= 32'hb26eb7b7;
    11'b00101011001: data <= 32'h39ecbd3c;
    11'b00101011010: data <= 32'h3dc9bcd9;
    11'b00101011011: data <= 32'h359a31a5;
    11'b00101011100: data <= 32'hbf6e3ce5;
    11'b00101011101: data <= 32'hc16e3b0a;
    11'b00101011110: data <= 32'hbd962b2f;
    11'b00101011111: data <= 32'h2ed8b0f4;
    11'b00101100000: data <= 32'ha6d6ae21;
    11'b00101100001: data <= 32'hbac1b5c6;
    11'b00101100010: data <= 32'hb57db436;
    11'b00101100011: data <= 32'h3d1f3c04;
    11'b00101100100: data <= 32'h3fb940d3;
    11'b00101100101: data <= 32'h3a864030;
    11'b00101100110: data <= 32'hb8013205;
    11'b00101100111: data <= 32'hb888bc43;
    11'b00101101000: data <= 32'h2eddb83c;
    11'b00101101001: data <= 32'h375132a8;
    11'b00101101010: data <= 32'h396eb8bc;
    11'b00101101011: data <= 32'h3d5bc001;
    11'b00101101100: data <= 32'h3ed4bf42;
    11'b00101101101: data <= 32'h394d2747;
    11'b00101101110: data <= 32'hbc8e3d1b;
    11'b00101101111: data <= 32'hbf1238ec;
    11'b00101110000: data <= 32'hbad9b9c2;
    11'b00101110001: data <= 32'hb385bc71;
    11'b00101110010: data <= 32'hbc36b9e8;
    11'b00101110011: data <= 32'hbf69b85f;
    11'b00101110100: data <= 32'hba83b50f;
    11'b00101110101: data <= 32'h3cd93989;
    11'b00101110110: data <= 32'h3ede3f85;
    11'b00101110111: data <= 32'h30b83f6d;
    11'b00101111000: data <= 32'hbd7339de;
    11'b00101111001: data <= 32'hbc633187;
    11'b00101111010: data <= 32'h302439eb;
    11'b00101111011: data <= 32'h39f83b07;
    11'b00101111100: data <= 32'h3a5fb840;
    11'b00101111101: data <= 32'h3cd7c007;
    11'b00101111110: data <= 32'h3ef4bdcc;
    11'b00101111111: data <= 32'h3d4d3925;
    11'b00110000000: data <= 32'h30a93e70;
    11'b00110000001: data <= 32'hb722358f;
    11'b00110000010: data <= 32'hb13abd6a;
    11'b00110000011: data <= 32'hb4eabe74;
    11'b00110000100: data <= 32'hbd9fbb51;
    11'b00110000101: data <= 32'hbfafb9be;
    11'b00110000110: data <= 32'hb86dbb9b;
    11'b00110000111: data <= 32'h3d4fb776;
    11'b00110001000: data <= 32'h3d1639a2;
    11'b00110001001: data <= 32'hb9d33d46;
    11'b00110001010: data <= 32'hc0463c2a;
    11'b00110001011: data <= 32'hbdc53b34;
    11'b00110001100: data <= 32'ha1893d0d;
    11'b00110001101: data <= 32'h351a3be6;
    11'b00110001110: data <= 32'hacefb785;
    11'b00110001111: data <= 32'h3507be19;
    11'b00110010000: data <= 32'h3dd9b82f;
    11'b00110010001: data <= 32'h3fa93e0e;
    11'b00110010010: data <= 32'h3cdc3fed;
    11'b00110010011: data <= 32'h371d3511;
    11'b00110010100: data <= 32'h3319bd23;
    11'b00110010101: data <= 32'hb16cbc97;
    11'b00110010110: data <= 32'hbc19b5be;
    11'b00110010111: data <= 32'hbc9eb99a;
    11'b00110011000: data <= 32'h32babf19;
    11'b00110011001: data <= 32'h3e60bf1f;
    11'b00110011010: data <= 32'h3c01b67a;
    11'b00110011011: data <= 32'hbc483a9b;
    11'b00110011100: data <= 32'hc0423bd8;
    11'b00110011101: data <= 32'hbce23a2d;
    11'b00110011110: data <= 32'hb12b3a89;
    11'b00110011111: data <= 32'hb8bc37e2;
    11'b00110100000: data <= 32'hbde4b845;
    11'b00110100001: data <= 32'hbac8bc11;
    11'b00110100010: data <= 32'h3c233189;
    11'b00110100011: data <= 32'h402e3f9c;
    11'b00110100100: data <= 32'h3dd4400c;
    11'b00110100101: data <= 32'h366b380c;
    11'b00110100110: data <= 32'h2b18b7be;
    11'b00110100111: data <= 32'ha20b2fef;
    11'b00110101000: data <= 32'hb575398f;
    11'b00110101001: data <= 32'hb3e4b743;
    11'b00110101010: data <= 32'h3aacc08f;
    11'b00110101011: data <= 32'h3f11c0ea;
    11'b00110101100: data <= 32'h3c62ba2d;
    11'b00110101101: data <= 32'hb86f39b0;
    11'b00110101110: data <= 32'hbcb2397c;
    11'b00110101111: data <= 32'hb69a2882;
    11'b00110110000: data <= 32'hb089b02e;
    11'b00110110001: data <= 32'hbda7b15e;
    11'b00110110010: data <= 32'hc11bb954;
    11'b00110110011: data <= 32'hbe45bb33;
    11'b00110110100: data <= 32'h3a022921;
    11'b00110110101: data <= 32'h3f483d7d;
    11'b00110110110: data <= 32'h3ac13e29;
    11'b00110110111: data <= 32'hb6a43991;
    11'b00110111000: data <= 32'hb79f3853;
    11'b00110111001: data <= 32'h28e13ddb;
    11'b00110111010: data <= 32'h2c983e90;
    11'b00110111011: data <= 32'h266eb054;
    11'b00110111100: data <= 32'h39c6c06a;
    11'b00110111101: data <= 32'h3e56c050;
    11'b00110111110: data <= 32'h3db0b3b9;
    11'b00110111111: data <= 32'h381a3c13;
    11'b00111000000: data <= 32'h32ee3673;
    11'b00111000001: data <= 32'h389bb975;
    11'b00111000010: data <= 32'h2d4dba14;
    11'b00111000011: data <= 32'hbe9eb5fc;
    11'b00111000100: data <= 32'hc165b94d;
    11'b00111000101: data <= 32'hbdb9bce8;
    11'b00111000110: data <= 32'h3a74bb3a;
    11'b00111000111: data <= 32'h3d72304d;
    11'b00111001000: data <= 32'had363990;
    11'b00111001001: data <= 32'hbd273967;
    11'b00111001010: data <= 32'hbae03c89;
    11'b00111001011: data <= 32'h28214026;
    11'b00111001100: data <= 32'had753fab;
    11'b00111001101: data <= 32'hb9222705;
    11'b00111001110: data <= 32'hb323becb;
    11'b00111001111: data <= 32'h3c03bcd5;
    11'b00111010000: data <= 32'h3ea83996;
    11'b00111010001: data <= 32'h3db63db8;
    11'b00111010010: data <= 32'h3cd33463;
    11'b00111010011: data <= 32'h3cb2babe;
    11'b00111010100: data <= 32'h35e7b7d7;
    11'b00111010101: data <= 32'hbcf632da;
    11'b00111010110: data <= 32'hbfbdb5b9;
    11'b00111010111: data <= 32'hb90ebecb;
    11'b00111011000: data <= 32'h3c6ec018;
    11'b00111011001: data <= 32'h3c17bc53;
    11'b00111011010: data <= 32'hb8f1aa97;
    11'b00111011011: data <= 32'hbdda36ad;
    11'b00111011100: data <= 32'hb8ff3ba5;
    11'b00111011101: data <= 32'h308b3ea2;
    11'b00111011110: data <= 32'hb9373db5;
    11'b00111011111: data <= 32'hbf70ab41;
    11'b00111100000: data <= 32'hbdf9bc93;
    11'b00111100001: data <= 32'h349fb5a6;
    11'b00111100010: data <= 32'h3e623d07;
    11'b00111100011: data <= 32'h3e673dec;
    11'b00111100100: data <= 32'h3cdd338c;
    11'b00111100101: data <= 32'h3c3cb5eb;
    11'b00111100110: data <= 32'h384338cc;
    11'b00111100111: data <= 32'hb8313d7f;
    11'b00111101000: data <= 32'hbb333245;
    11'b00111101001: data <= 32'h30c5bfb1;
    11'b00111101010: data <= 32'h3d3cc146;
    11'b00111101011: data <= 32'h3b69be1a;
    11'b00111101100: data <= 32'hb681b456;
    11'b00111101101: data <= 32'hb98a2cfc;
    11'b00111101110: data <= 32'h347a3216;
    11'b00111101111: data <= 32'h37a238ef;
    11'b00111110000: data <= 32'hbcab3908;
    11'b00111110001: data <= 32'hc1abb372;
    11'b00111110010: data <= 32'hc0a0baf9;
    11'b00111110011: data <= 32'hb0dbb28f;
    11'b00111110100: data <= 32'h3cf23b54;
    11'b00111110101: data <= 32'h3ba43b54;
    11'b00111110110: data <= 32'h356d2f4c;
    11'b00111110111: data <= 32'h36b9355a;
    11'b00111111000: data <= 32'h38433f4d;
    11'b00111111001: data <= 32'h20ba40e0;
    11'b00111111010: data <= 32'hb5fa39c4;
    11'b00111111011: data <= 32'h335ebedc;
    11'b00111111100: data <= 32'h3c48c097;
    11'b00111111101: data <= 32'h3ba3bbbd;
    11'b00111111110: data <= 32'h355a2eb8;
    11'b00111111111: data <= 32'h3898b12d;
    11'b01000000000: data <= 32'h3d9cb8f7;
    11'b01000000001: data <= 32'h3b9cb3a7;
    11'b01000000010: data <= 32'hbceb3346;
    11'b01000000011: data <= 32'hc1ddb27d;
    11'b01000000100: data <= 32'hc05dbb6a;
    11'b01000000101: data <= 32'hacb1ba94;
    11'b01000000110: data <= 32'h3a68b1fe;
    11'b01000000111: data <= 32'ha9cfac7f;
    11'b01000001000: data <= 32'hb9dbb217;
    11'b01000001001: data <= 32'hb0f839b1;
    11'b01000001010: data <= 32'h383440c4;
    11'b01000001011: data <= 32'h2de74183;
    11'b01000001100: data <= 32'hb9c53b4d;
    11'b01000001101: data <= 32'hb888bccd;
    11'b01000001110: data <= 32'h35a2bd22;
    11'b01000001111: data <= 32'h3b203086;
    11'b01000010000: data <= 32'h3c013996;
    11'b01000010001: data <= 32'h3e05b447;
    11'b01000010010: data <= 32'h4029bbe8;
    11'b01000010011: data <= 32'h3d4ab46b;
    11'b01000010100: data <= 32'hba373938;
    11'b01000010101: data <= 32'hc0393329;
    11'b01000010110: data <= 32'hbcfbbc55;
    11'b01000010111: data <= 32'h363fbec7;
    11'b01000011000: data <= 32'h37f6bd5a;
    11'b01000011001: data <= 32'hba14bb72;
    11'b01000011010: data <= 32'hbcccb8bb;
    11'b01000011011: data <= 32'hae44374a;
    11'b01000011100: data <= 32'h39dc3fa9;
    11'b01000011101: data <= 32'hb1494054;
    11'b01000011110: data <= 32'hbe9a398e;
    11'b01000011111: data <= 32'hbf0eb97a;
    11'b01000100000: data <= 32'hb805b460;
    11'b01000100001: data <= 32'h39023bd5;
    11'b01000100010: data <= 32'h3c3a3b84;
    11'b01000100011: data <= 32'h3de4b600;
    11'b01000100100: data <= 32'h3fa2ba7a;
    11'b01000100101: data <= 32'h3d913821;
    11'b01000100110: data <= 32'hadfc3ee9;
    11'b01000100111: data <= 32'hbb8d3b75;
    11'b01000101000: data <= 32'hb271bc47;
    11'b01000101001: data <= 32'h3a57c042;
    11'b01000101010: data <= 32'h35c3befb;
    11'b01000101011: data <= 32'hba98bc90;
    11'b01000101100: data <= 32'hb9dabb19;
    11'b01000101101: data <= 32'h39a8b4ac;
    11'b01000101110: data <= 32'h3ce73a14;
    11'b01000101111: data <= 32'hb6963c81;
    11'b01000110000: data <= 32'hc0e234fe;
    11'b01000110001: data <= 32'hc119b65f;
    11'b01000110010: data <= 32'hbbd8302c;
    11'b01000110011: data <= 32'h340c3b90;
    11'b01000110100: data <= 32'h367937e4;
    11'b01000110101: data <= 32'h37fcb932;
    11'b01000110110: data <= 32'h3c3ab649;
    11'b01000110111: data <= 32'h3cc43e21;
    11'b01000111000: data <= 32'h36ee4186;
    11'b01000111001: data <= 32'hb1d73e26;
    11'b01000111010: data <= 32'h3221ba50;
    11'b01000111011: data <= 32'h3992bf01;
    11'b01000111100: data <= 32'h3407bc6d;
    11'b01000111101: data <= 32'hb616b8bb;
    11'b01000111110: data <= 32'h34e8bb94;
    11'b01000111111: data <= 32'h3f34bc56;
    11'b01001000000: data <= 32'h3f45b4f3;
    11'b01001000001: data <= 32'hb5963695;
    11'b01001000010: data <= 32'hc0f1318e;
    11'b01001000011: data <= 32'hc0b5b571;
    11'b01001000100: data <= 32'hba30b208;
    11'b01001000101: data <= 32'ha8a72dc1;
    11'b01001000110: data <= 32'hb89bb756;
    11'b01001000111: data <= 32'hba1ebc65;
    11'b01001001000: data <= 32'h3194b1fb;
    11'b01001001001: data <= 32'h3bf23ffc;
    11'b01001001010: data <= 32'h38ce4211;
    11'b01001001011: data <= 32'hb38f3e9a;
    11'b01001001100: data <= 32'hb566b60d;
    11'b01001001101: data <= 32'h26e7ba00;
    11'b01001001110: data <= 32'h265431a6;
    11'b01001001111: data <= 32'h2ce534be;
    11'b01001010000: data <= 32'h3c7abac8;
    11'b01001010001: data <= 32'h40e6be09;
    11'b01001010010: data <= 32'h4053b90c;
    11'b01001010011: data <= 32'h2a3e3866;
    11'b01001010100: data <= 32'hbe993839;
    11'b01001010101: data <= 32'hbd0cb54a;
    11'b01001010110: data <= 32'ha8a1ba8e;
    11'b01001010111: data <= 32'hb038bb5b;
    11'b01001011000: data <= 32'hbd4ebd3c;
    11'b01001011001: data <= 32'hbe06be1c;
    11'b01001011010: data <= 32'hac96b709;
    11'b01001011011: data <= 32'h3c663e0d;
    11'b01001011100: data <= 32'h3801409e;
    11'b01001011101: data <= 32'hbb3a3cc1;
    11'b01001011110: data <= 32'hbd7aabec;
    11'b01001011111: data <= 32'hba9d3484;
    11'b01001100000: data <= 32'hb50c3d1c;
    11'b01001100001: data <= 32'h2d513ad6;
    11'b01001100010: data <= 32'h3c39ba9a;
    11'b01001100011: data <= 32'h4059bde2;
    11'b01001100100: data <= 32'h400faf3c;
    11'b01001100101: data <= 32'h386b3dbd;
    11'b01001100110: data <= 32'hb7723cf1;
    11'b01001100111: data <= 32'h2879b27b;
    11'b01001101000: data <= 32'h398abc9f;
    11'b01001101001: data <= 32'haf2bbd1d;
    11'b01001101010: data <= 32'hbe0dbdc8;
    11'b01001101011: data <= 32'hbd48beb0;
    11'b01001101100: data <= 32'h3827bc27;
    11'b01001101101: data <= 32'h3e553583;
    11'b01001101110: data <= 32'h364c3c1f;
    11'b01001101111: data <= 32'hbe37379f;
    11'b01001110000: data <= 32'hc02e29ba;
    11'b01001110001: data <= 32'hbd0c3a51;
    11'b01001110010: data <= 32'hb8c13e22;
    11'b01001110011: data <= 32'hb75e3932;
    11'b01001110100: data <= 32'h2c6bbc49;
    11'b01001110101: data <= 32'h3c6bbcd3;
    11'b01001110110: data <= 32'h3e0839d6;
    11'b01001110111: data <= 32'h3b1240c5;
    11'b01001111000: data <= 32'h361b3f4b;
    11'b01001111001: data <= 32'h39cb2920;
    11'b01001111010: data <= 32'h3aefbaba;
    11'b01001111011: data <= 32'hb15eb8fc;
    11'b01001111100: data <= 32'hbce7b9a6;
    11'b01001111101: data <= 32'hb7c0bdbc;
    11'b01001111110: data <= 32'h3e0cbe86;
    11'b01001111111: data <= 32'h405aba5d;
    11'b01010000000: data <= 32'h3783240c;
    11'b01010000001: data <= 32'hbe6828d6;
    11'b01010000010: data <= 32'hbf7d250c;
    11'b01010000011: data <= 32'hbb2f3901;
    11'b01010000100: data <= 32'hb8f93b3d;
    11'b01010000101: data <= 32'hbd02b1c2;
    11'b01010000110: data <= 32'hbd05be24;
    11'b01010000111: data <= 32'hace1bc3b;
    11'b01010001000: data <= 32'h3be03cae;
    11'b01010001001: data <= 32'h3b7d4143;
    11'b01010001010: data <= 32'h379a3f43;
    11'b01010001011: data <= 32'h37243380;
    11'b01010001100: data <= 32'h3593a007;
    11'b01010001101: data <= 32'hb69339b3;
    11'b01010001110: data <= 32'hbae4378c;
    11'b01010001111: data <= 32'h344bbbf6;
    11'b01010010000: data <= 32'h4043bfa6;
    11'b01010010001: data <= 32'h40e0bd03;
    11'b01010010010: data <= 32'h399cafa6;
    11'b01010010011: data <= 32'hbb5c3299;
    11'b01010010100: data <= 32'hb9da2879;
    11'b01010010101: data <= 32'h2f532f42;
    11'b01010010110: data <= 32'hb608a088;
    11'b01010010111: data <= 32'hbf5cbbf8;
    11'b01010011000: data <= 32'hc03ebfac;
    11'b01010011001: data <= 32'hb8ecbcca;
    11'b01010011010: data <= 32'h3aee3a5e;
    11'b01010011011: data <= 32'h3a903f75;
    11'b01010011100: data <= 32'hab3a3c67;
    11'b01010011101: data <= 32'hb7473317;
    11'b01010011110: data <= 32'hb75e3ad4;
    11'b01010011111: data <= 32'hb9e73fb9;
    11'b01010100000: data <= 32'hba5b3d5b;
    11'b01010100001: data <= 32'h3483b9b0;
    11'b01010100010: data <= 32'h3f4abf53;
    11'b01010100011: data <= 32'h402bbb08;
    11'b01010100100: data <= 32'h3b2f38cf;
    11'b01010100101: data <= 32'h2df53acb;
    11'b01010100110: data <= 32'h396b3181;
    11'b01010100111: data <= 32'h3ca9b379;
    11'b01010101000: data <= 32'hac07b69c;
    11'b01010101001: data <= 32'hbfd2bc70;
    11'b01010101010: data <= 32'hc02abf88;
    11'b01010101011: data <= 32'hb315be17;
    11'b01010101100: data <= 32'h3d07b2ac;
    11'b01010101101: data <= 32'h39da37b3;
    11'b01010101110: data <= 32'hb96a2bdc;
    11'b01010101111: data <= 32'hbcbf2052;
    11'b01010110000: data <= 32'hbb0e3d0f;
    11'b01010110001: data <= 32'hbb1040ac;
    11'b01010110010: data <= 32'hbc703d74;
    11'b01010110011: data <= 32'hb86dbaa5;
    11'b01010110100: data <= 32'h3945be54;
    11'b01010110101: data <= 32'h3cf5ae49;
    11'b01010110110: data <= 32'h3b263e20;
    11'b01010110111: data <= 32'h3a993db6;
    11'b01010111000: data <= 32'h3e153531;
    11'b01010111001: data <= 32'h3e69ae54;
    11'b01010111010: data <= 32'h29eb2f05;
    11'b01010111011: data <= 32'hbeb1b4a9;
    11'b01010111100: data <= 32'hbd54bd5b;
    11'b01010111101: data <= 32'h39bfbf1b;
    11'b01010111110: data <= 32'h3f5bbce0;
    11'b01010111111: data <= 32'h3a09b988;
    11'b01011000000: data <= 32'hbad8b964;
    11'b01011000001: data <= 32'hbc53b326;
    11'b01011000010: data <= 32'hb74c3c5c;
    11'b01011000011: data <= 32'hb9143f43;
    11'b01011000100: data <= 32'hbe4b38f7;
    11'b01011000101: data <= 32'hbef4bd18;
    11'b01011000110: data <= 32'hb970bda3;
    11'b01011000111: data <= 32'h364436de;
    11'b01011001000: data <= 32'h39943f79;
    11'b01011001001: data <= 32'h3b1a3d81;
    11'b01011001010: data <= 32'h3d7b3484;
    11'b01011001011: data <= 32'h3cd636e6;
    11'b01011001100: data <= 32'hb1083d39;
    11'b01011001101: data <= 32'hbd383c28;
    11'b01011001110: data <= 32'hb840b878;
    11'b01011001111: data <= 32'h3da3bf18;
    11'b01011010000: data <= 32'h4026be7f;
    11'b01011010001: data <= 32'h3a56bbc8;
    11'b01011010010: data <= 32'hb71db967;
    11'b01011010011: data <= 32'hacdeb470;
    11'b01011010100: data <= 32'h399838ad;
    11'b01011010101: data <= 32'ha9a03b1e;
    11'b01011010110: data <= 32'hbf69b3d7;
    11'b01011010111: data <= 32'hc112be99;
    11'b01011011000: data <= 32'hbd86bd98;
    11'b01011011001: data <= 32'h2b4d34a7;
    11'b01011011010: data <= 32'h37923cec;
    11'b01011011011: data <= 32'h35d23843;
    11'b01011011100: data <= 32'h37dbac6e;
    11'b01011011101: data <= 32'h360c3bc8;
    11'b01011011110: data <= 32'hb7d140e2;
    11'b01011011111: data <= 32'hbc844029;
    11'b01011100000: data <= 32'hb51ba384;
    11'b01011100001: data <= 32'h3ce6be2a;
    11'b01011100010: data <= 32'h3e75bd01;
    11'b01011100011: data <= 32'h3959b4e3;
    11'b01011100100: data <= 32'h33f7a9b4;
    11'b01011100101: data <= 32'h3cf8b054;
    11'b01011100110: data <= 32'h3fbe314f;
    11'b01011100111: data <= 32'h388a352f;
    11'b01011101000: data <= 32'hbf19b7ac;
    11'b01011101001: data <= 32'hc0f9be22;
    11'b01011101010: data <= 32'hbc48bdbb;
    11'b01011101011: data <= 32'h364fb672;
    11'b01011101100: data <= 32'h3607ab6a;
    11'b01011101101: data <= 32'hb4cfb998;
    11'b01011101110: data <= 32'hb5d8b8e1;
    11'b01011101111: data <= 32'hb1023c9e;
    11'b01011110000: data <= 32'hb8a941a7;
    11'b01011110001: data <= 32'hbcc44070;
    11'b01011110010: data <= 32'hbae1a86f;
    11'b01011110011: data <= 32'h3130bd0b;
    11'b01011110100: data <= 32'h38a2b718;
    11'b01011110101: data <= 32'h351339b5;
    11'b01011110110: data <= 32'h39c73912;
    11'b01011110111: data <= 32'h401e9f1f;
    11'b01011111000: data <= 32'h41082dd1;
    11'b01011111001: data <= 32'h3a9c3898;
    11'b01011111010: data <= 32'hbdb83362;
    11'b01011111011: data <= 32'hbee0ba7f;
    11'b01011111100: data <= 32'hacd7bd55;
    11'b01011111101: data <= 32'h3c3abc88;
    11'b01011111110: data <= 32'h364ebcca;
    11'b01011111111: data <= 32'hb92ebe6f;
    11'b01100000000: data <= 32'hb80cbc2b;
    11'b01100000001: data <= 32'h30e83b0f;
    11'b01100000010: data <= 32'hb1cb4096;
    11'b01100000011: data <= 32'hbd3d3dd2;
    11'b01100000100: data <= 32'hbf03b841;
    11'b01100000101: data <= 32'hbc8cbc5d;
    11'b01100000110: data <= 32'hb77b32f8;
    11'b01100000111: data <= 32'hb0293d13;
    11'b01100001000: data <= 32'h393439a3;
    11'b01100001001: data <= 32'h3f9bb18d;
    11'b01100001010: data <= 32'h404834c0;
    11'b01100001011: data <= 32'h38d43de7;
    11'b01100001100: data <= 32'hbc413e0d;
    11'b01100001101: data <= 32'hba8031d8;
    11'b01100001110: data <= 32'h3a79bc26;
    11'b01100001111: data <= 32'h3daebd78;
    11'b01100010000: data <= 32'h356abde6;
    11'b01100010001: data <= 32'hb841beaf;
    11'b01100010010: data <= 32'h32b7bc7d;
    11'b01100010011: data <= 32'h3d0135e5;
    11'b01100010100: data <= 32'h39073d25;
    11'b01100010101: data <= 32'hbd1036c4;
    11'b01100010110: data <= 32'hc0b1bc24;
    11'b01100010111: data <= 32'hbf59bc11;
    11'b01100011000: data <= 32'hbb43357c;
    11'b01100011001: data <= 32'hb6ed3b4c;
    11'b01100011010: data <= 32'h2e38ac71;
    11'b01100011011: data <= 32'h3bb0b9e6;
    11'b01100011100: data <= 32'h3cb237ff;
    11'b01100011101: data <= 32'h30c540c5;
    11'b01100011110: data <= 32'hbacf411c;
    11'b01100011111: data <= 32'hb5e53afd;
    11'b01100100000: data <= 32'h3b2ab959;
    11'b01100100001: data <= 32'h3c2cbb7e;
    11'b01100100010: data <= 32'h24d2ba1f;
    11'b01100100011: data <= 32'hb1c9bb89;
    11'b01100100100: data <= 32'h3d25bafd;
    11'b01100100101: data <= 32'h40faac52;
    11'b01100100110: data <= 32'h3db0382a;
    11'b01100100111: data <= 32'hbbfdacb3;
    11'b01100101000: data <= 32'hc06abc16;
    11'b01100101001: data <= 32'hbdfebb08;
    11'b01100101010: data <= 32'hb822a37f;
    11'b01100101011: data <= 32'hb73dafe1;
    11'b01100101100: data <= 32'hb89abd34;
    11'b01100101101: data <= 32'hac30bdf3;
    11'b01100101110: data <= 32'h36433725;
    11'b01100101111: data <= 32'hac45414d;
    11'b01100110000: data <= 32'hba2d415c;
    11'b01100110001: data <= 32'hb8b03ac8;
    11'b01100110010: data <= 32'h2e0db6ca;
    11'b01100110011: data <= 32'h23b1af89;
    11'b01100110100: data <= 32'hb87c365c;
    11'b01100110101: data <= 32'h2515a856;
    11'b01100110110: data <= 32'h3fd6b8e0;
    11'b01100110111: data <= 32'h4225b402;
    11'b01100111000: data <= 32'h3ee7377c;
    11'b01100111001: data <= 32'hb92335e2;
    11'b01100111010: data <= 32'hbdabb52a;
    11'b01100111011: data <= 32'hb623b85c;
    11'b01100111100: data <= 32'h3598b71b;
    11'b01100111101: data <= 32'hb4bcbc64;
    11'b01100111110: data <= 32'hbc01c075;
    11'b01100111111: data <= 32'hb7c6c008;
    11'b01101000000: data <= 32'h36d32f13;
    11'b01101000001: data <= 32'h34a74028;
    11'b01101000010: data <= 32'hb9513f46;
    11'b01101000011: data <= 32'hbca431b5;
    11'b01101000100: data <= 32'hbc15b62c;
    11'b01101000101: data <= 32'hbc4138cd;
    11'b01101000110: data <= 32'hbc9c3cd6;
    11'b01101000111: data <= 32'hb15e3506;
    11'b01101001000: data <= 32'h3efab9a6;
    11'b01101001001: data <= 32'h4140b405;
    11'b01101001010: data <= 32'h3d7b3c2d;
    11'b01101001011: data <= 32'hb6383dcb;
    11'b01101001100: data <= 32'hb77939ab;
    11'b01101001101: data <= 32'h39e3ac0f;
    11'b01101001110: data <= 32'h3becb81a;
    11'b01101001111: data <= 32'hb41cbd35;
    11'b01101010000: data <= 32'hbc43c07f;
    11'b01101010001: data <= 32'hadf8c006;
    11'b01101010010: data <= 32'h3d3ab51a;
    11'b01101010011: data <= 32'h3c883c22;
    11'b01101010100: data <= 32'hb6813893;
    11'b01101010101: data <= 32'hbe2db8c6;
    11'b01101010110: data <= 32'hbe84b6d4;
    11'b01101010111: data <= 32'hbdf73b09;
    11'b01101011000: data <= 32'hbdb63cad;
    11'b01101011001: data <= 32'hb966b341;
    11'b01101011010: data <= 32'h3a25bd28;
    11'b01101011011: data <= 32'h3ddeb46f;
    11'b01101011100: data <= 32'h393f3ed5;
    11'b01101011101: data <= 32'hb4e840c3;
    11'b01101011110: data <= 32'h2edb3da8;
    11'b01101011111: data <= 32'h3c873564;
    11'b01101100000: data <= 32'h3ae6ad2f;
    11'b01101100001: data <= 32'hb89db86c;
    11'b01101100010: data <= 32'hbb92bd6f;
    11'b01101100011: data <= 32'h39b7be1a;
    11'b01101100100: data <= 32'h40d6b8f3;
    11'b01101100101: data <= 32'h3fdb3117;
    11'b01101100110: data <= 32'haaa3b33a;
    11'b01101100111: data <= 32'hbd6cbacf;
    11'b01101101000: data <= 32'hbcfbb507;
    11'b01101101001: data <= 32'hbbc739fa;
    11'b01101101010: data <= 32'hbcfc36b4;
    11'b01101101011: data <= 32'hbcdfbd45;
    11'b01101101100: data <= 32'hb596c02f;
    11'b01101101101: data <= 32'h3648b76e;
    11'b01101101110: data <= 32'h30fe3f84;
    11'b01101101111: data <= 32'hb48140e7;
    11'b01101110000: data <= 32'h2e803d30;
    11'b01101110001: data <= 32'h390936d7;
    11'b01101110010: data <= 32'h9f383906;
    11'b01101110011: data <= 32'hbcdc3980;
    11'b01101110100: data <= 32'hbb56b195;
    11'b01101110101: data <= 32'h3d01bbc0;
    11'b01101110110: data <= 32'h41e2b9c1;
    11'b01101110111: data <= 32'h406dada8;
    11'b01101111000: data <= 32'h3290ae0f;
    11'b01101111001: data <= 32'hb928b558;
    11'b01101111010: data <= 32'haba62cd2;
    11'b01101111011: data <= 32'h30c23822;
    11'b01101111100: data <= 32'hba63b62b;
    11'b01101111101: data <= 32'hbe27c05c;
    11'b01101111110: data <= 32'hbb8ec135;
    11'b01101111111: data <= 32'h2f01ba0f;
    11'b01110000000: data <= 32'h34d83d67;
    11'b01110000001: data <= 32'hb0473e1a;
    11'b01110000010: data <= 32'hb41c3665;
    11'b01110000011: data <= 32'hb48d3209;
    11'b01110000100: data <= 32'hbc0f3cea;
    11'b01110000101: data <= 32'hbf4f3ea0;
    11'b01110000110: data <= 32'hbc7837f1;
    11'b01110000111: data <= 32'h3c2eba9a;
    11'b01110001000: data <= 32'h40deb9e2;
    11'b01110001001: data <= 32'h3ea6343f;
    11'b01110001010: data <= 32'h329c3a0d;
    11'b01110001011: data <= 32'h320338ea;
    11'b01110001100: data <= 32'h3cd038d9;
    11'b01110001101: data <= 32'h3c74381f;
    11'b01110001110: data <= 32'hb7e6b87c;
    11'b01110001111: data <= 32'hbe5cc04b;
    11'b01110010000: data <= 32'hba2cc0e4;
    11'b01110010001: data <= 32'h39e2bbc5;
    11'b01110010010: data <= 32'h3c2b36a2;
    11'b01110010011: data <= 32'h321430ad;
    11'b01110010100: data <= 32'hb836b993;
    11'b01110010101: data <= 32'hbaa0b065;
    11'b01110010110: data <= 32'hbd983ddf;
    11'b01110010111: data <= 32'hbffa3f51;
    11'b01110011000: data <= 32'hbdd2336a;
    11'b01110011001: data <= 32'h312cbd1f;
    11'b01110011010: data <= 32'h3c9ebaa3;
    11'b01110011011: data <= 32'h39153a3e;
    11'b01110011100: data <= 32'ha0193e5d;
    11'b01110011101: data <= 32'h39993d21;
    11'b01110011110: data <= 32'h3f393b91;
    11'b01110011111: data <= 32'h3d213aa6;
    11'b01110100000: data <= 32'hb93d2f6d;
    11'b01110100001: data <= 32'hbe1fbc99;
    11'b01110100010: data <= 32'hb067beaa;
    11'b01110100011: data <= 32'h3edfbbca;
    11'b01110100100: data <= 32'h3f58b61b;
    11'b01110100101: data <= 32'h3839bad4;
    11'b01110100110: data <= 32'hb65fbd13;
    11'b01110100111: data <= 32'hb7dab2ef;
    11'b01110101000: data <= 32'hba4f3d86;
    11'b01110101001: data <= 32'hbe343d14;
    11'b01110101010: data <= 32'hbedbb99b;
    11'b01110101011: data <= 32'hbaf0c015;
    11'b01110101100: data <= 32'haf5cbc24;
    11'b01110101101: data <= 32'hb2713baa;
    11'b01110101110: data <= 32'hb2b03eb9;
    11'b01110101111: data <= 32'h39c33c5e;
    11'b01110110000: data <= 32'h3e073a89;
    11'b01110110001: data <= 32'h38cf3d21;
    11'b01110110010: data <= 32'hbcf53d11;
    11'b01110110011: data <= 32'hbe2f330c;
    11'b01110110100: data <= 32'h35c4ba15;
    11'b01110110101: data <= 32'h4078ba87;
    11'b01110110110: data <= 32'h400fb910;
    11'b01110110111: data <= 32'h38e8bb7d;
    11'b01110111000: data <= 32'h2e07bbc9;
    11'b01110111001: data <= 32'h38e22e57;
    11'b01110111010: data <= 32'h380d3cd8;
    11'b01110111011: data <= 32'hba083856;
    11'b01110111100: data <= 32'hbf03be22;
    11'b01110111101: data <= 32'hbdc7c108;
    11'b01110111110: data <= 32'hb8f6bcd3;
    11'b01110111111: data <= 32'hb4fc38d6;
    11'b01111000000: data <= 32'hb1463a9e;
    11'b01111000001: data <= 32'h36d7289d;
    11'b01111000010: data <= 32'h39a033b5;
    11'b01111000011: data <= 32'hb59e3e5e;
    11'b01111000100: data <= 32'hbf504066;
    11'b01111000101: data <= 32'hbeaf3c79;
    11'b01111000110: data <= 32'h3488b530;
    11'b01111000111: data <= 32'h3f26b987;
    11'b01111001000: data <= 32'h3d5cb571;
    11'b01111001001: data <= 32'h34d0b335;
    11'b01111001010: data <= 32'h391daef3;
    11'b01111001011: data <= 32'h3f4f38ea;
    11'b01111001100: data <= 32'h3ecd3cb6;
    11'b01111001101: data <= 32'hb00b3485;
    11'b01111001110: data <= 32'hbe80be32;
    11'b01111001111: data <= 32'hbd48c07b;
    11'b01111010000: data <= 32'hb122bc8e;
    11'b01111010001: data <= 32'h34f3ab88;
    11'b01111010010: data <= 32'h307ab805;
    11'b01111010011: data <= 32'h3135bd2a;
    11'b01111010100: data <= 32'h2f95b6e5;
    11'b01111010101: data <= 32'hba2e3e77;
    11'b01111010110: data <= 32'hbfa440d0;
    11'b01111010111: data <= 32'hbf153c2a;
    11'b01111011000: data <= 32'hb599b8f9;
    11'b01111011001: data <= 32'h3877ba01;
    11'b01111011010: data <= 32'h2d8b30a3;
    11'b01111011011: data <= 32'hb46138e0;
    11'b01111011100: data <= 32'h3b4738aa;
    11'b01111011101: data <= 32'h40e73b32;
    11'b01111011110: data <= 32'h40283d37;
    11'b01111011111: data <= 32'hadab39ea;
    11'b01111100000: data <= 32'hbe05b8d4;
    11'b01111100001: data <= 32'hb9d7bcfd;
    11'b01111100010: data <= 32'h3a47ba3a;
    11'b01111100011: data <= 32'h3c6eb8c3;
    11'b01111100100: data <= 32'h372abe0e;
    11'b01111100101: data <= 32'h30dfc02f;
    11'b01111100110: data <= 32'h3455ba03;
    11'b01111100111: data <= 32'hb2fa3dc0;
    11'b01111101000: data <= 32'hbd193f95;
    11'b01111101001: data <= 32'hbeb531c1;
    11'b01111101010: data <= 32'hbc71bd74;
    11'b01111101011: data <= 32'hb9bbbb89;
    11'b01111101100: data <= 32'hbbfe36a5;
    11'b01111101101: data <= 32'hba113ac6;
    11'b01111101110: data <= 32'h3a6f3731;
    11'b01111101111: data <= 32'h406738de;
    11'b01111110000: data <= 32'h3e013db7;
    11'b01111110001: data <= 32'hb8ff3e7d;
    11'b01111110010: data <= 32'hbe0a3a1d;
    11'b01111110011: data <= 32'hb1a8ad18;
    11'b01111110100: data <= 32'h3da7b4ca;
    11'b01111110101: data <= 32'h3d6eb97e;
    11'b01111110110: data <= 32'h367cbe97;
    11'b01111110111: data <= 32'h35abbfbd;
    11'b01111111000: data <= 32'h3c76b82c;
    11'b01111111001: data <= 32'h3c443d02;
    11'b01111111010: data <= 32'hb2ca3c92;
    11'b01111111011: data <= 32'hbd77b9d9;
    11'b01111111100: data <= 32'hbdfbbf90;
    11'b01111111101: data <= 32'hbd16bc12;
    11'b01111111110: data <= 32'hbd2334f5;
    11'b01111111111: data <= 32'hbac1335f;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    