
module memory_rom_52(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3e09b76d;
    11'b00000000001: data <= 32'h3af5b56f;
    11'b00000000010: data <= 32'hbad833c6;
    11'b00000000011: data <= 32'hbf66b46c;
    11'b00000000100: data <= 32'hb9b4be44;
    11'b00000000101: data <= 32'h3cb9c00c;
    11'b00000000110: data <= 32'h3d77bd2a;
    11'b00000000111: data <= 32'hb3a9b7be;
    11'b00000001000: data <= 32'hbd62ae40;
    11'b00000001001: data <= 32'hba213875;
    11'b00000001010: data <= 32'ha0303e18;
    11'b00000001011: data <= 32'hb9623e0f;
    11'b00000001100: data <= 32'hbf962474;
    11'b00000001101: data <= 32'hbf0bbd21;
    11'b00000001110: data <= 32'hb2cab8f0;
    11'b00000001111: data <= 32'h3c4b3ca9;
    11'b00000010000: data <= 32'h3d1e3ed1;
    11'b00000010001: data <= 32'h3cb138b1;
    11'b00000010010: data <= 32'h3cdeb125;
    11'b00000010011: data <= 32'h39c33965;
    11'b00000010100: data <= 32'hb77a3e44;
    11'b00000010101: data <= 32'hbbd5391e;
    11'b00000010110: data <= 32'h2febbdb1;
    11'b00000010111: data <= 32'h3e1fc0c8;
    11'b00000011000: data <= 32'h3d5ebe93;
    11'b00000011001: data <= 32'habe7b8c0;
    11'b00000011010: data <= 32'hb88ab330;
    11'b00000011011: data <= 32'h358b2607;
    11'b00000011100: data <= 32'h39ca387e;
    11'b00000011101: data <= 32'hba4b3889;
    11'b00000011110: data <= 32'hc14cb6e7;
    11'b00000011111: data <= 32'hc117bce2;
    11'b00000100000: data <= 32'hb94cb85b;
    11'b00000100001: data <= 32'h3a413a2d;
    11'b00000100010: data <= 32'h39e83b94;
    11'b00000100011: data <= 32'h347b2eb3;
    11'b00000100100: data <= 32'h358d31b1;
    11'b00000100101: data <= 32'h35c23ee7;
    11'b00000100110: data <= 32'hb37b4161;
    11'b00000100111: data <= 32'hb8ac3d46;
    11'b00000101000: data <= 32'h313fbc7d;
    11'b00000101001: data <= 32'h3cb2c00f;
    11'b00000101010: data <= 32'h3c72bbf9;
    11'b00000101011: data <= 32'h36802a58;
    11'b00000101100: data <= 32'h38e0acce;
    11'b00000101101: data <= 32'h3e87b767;
    11'b00000101110: data <= 32'h3df3b164;
    11'b00000101111: data <= 32'hb8ef3087;
    11'b00000110000: data <= 32'hc141b67d;
    11'b00000110001: data <= 32'hc099bca4;
    11'b00000110010: data <= 32'hb57cbc0b;
    11'b00000110011: data <= 32'h398eb550;
    11'b00000110100: data <= 32'h2599b489;
    11'b00000110101: data <= 32'hb9c8b8aa;
    11'b00000110110: data <= 32'hb5a7336e;
    11'b00000110111: data <= 32'h3285403d;
    11'b00000111000: data <= 32'hb1ff41d9;
    11'b00000111001: data <= 32'hbb303d71;
    11'b00000111010: data <= 32'hb99abace;
    11'b00000111011: data <= 32'h31a5bcd7;
    11'b00000111100: data <= 32'h39133020;
    11'b00000111101: data <= 32'h39d13b01;
    11'b00000111110: data <= 32'h3d922e88;
    11'b00000111111: data <= 32'h409db951;
    11'b00001000000: data <= 32'h3f62b109;
    11'b00001000001: data <= 32'hb4293935;
    11'b00001000010: data <= 32'hbf8a345d;
    11'b00001000011: data <= 32'hbd0cbb8d;
    11'b00001000100: data <= 32'h36eebe51;
    11'b00001000101: data <= 32'h3a1fbd99;
    11'b00001000110: data <= 32'hb723bd04;
    11'b00001000111: data <= 32'hbc75bc80;
    11'b00001001000: data <= 32'hb411ad3f;
    11'b00001001001: data <= 32'h38923e7e;
    11'b00001001010: data <= 32'hb179405c;
    11'b00001001011: data <= 32'hbe733a6e;
    11'b00001001100: data <= 32'hbf9fb9e1;
    11'b00001001101: data <= 32'hbb3ab76f;
    11'b00001001110: data <= 32'h2dca3b58;
    11'b00001001111: data <= 32'h38c83cac;
    11'b00001010000: data <= 32'h3d08a730;
    11'b00001010001: data <= 32'h3fe9b8fb;
    11'b00001010010: data <= 32'h3e783835;
    11'b00001010011: data <= 32'h2c7a3f45;
    11'b00001010100: data <= 32'hbb7b3d2c;
    11'b00001010101: data <= 32'hb248b873;
    11'b00001010110: data <= 32'h3c07bf05;
    11'b00001010111: data <= 32'h3a16bec2;
    11'b00001011000: data <= 32'hb807bd74;
    11'b00001011001: data <= 32'hb94bbce6;
    11'b00001011010: data <= 32'h3983b8a8;
    11'b00001011011: data <= 32'h3da038c2;
    11'b00001011100: data <= 32'ha3343c1d;
    11'b00001011101: data <= 32'hc044304a;
    11'b00001011110: data <= 32'hc13bb9be;
    11'b00001011111: data <= 32'hbd8db1e4;
    11'b00001100000: data <= 32'hb36c3ac0;
    11'b00001100001: data <= 32'h2af938be;
    11'b00001100010: data <= 32'h34ebb8d4;
    11'b00001100011: data <= 32'h3b7ab88d;
    11'b00001100100: data <= 32'h3c323d46;
    11'b00001100101: data <= 32'h33b441b7;
    11'b00001100110: data <= 32'hb5c54013;
    11'b00001100111: data <= 32'h30f4b158;
    11'b00001101000: data <= 32'h3accbd64;
    11'b00001101001: data <= 32'h3749bbe8;
    11'b00001101010: data <= 32'hb52eb8a7;
    11'b00001101011: data <= 32'h3392bb25;
    11'b00001101100: data <= 32'h3f89bbfb;
    11'b00001101101: data <= 32'h4087b49c;
    11'b00001101110: data <= 32'h34c634d6;
    11'b00001101111: data <= 32'hc00cab4c;
    11'b00001110000: data <= 32'hc0a2b8dc;
    11'b00001110001: data <= 32'hbbbfb5e9;
    11'b00001110010: data <= 32'hb19a2845;
    11'b00001110011: data <= 32'hb8c5b84c;
    11'b00001110100: data <= 32'hba9cbda0;
    11'b00001110101: data <= 32'haa90b9a2;
    11'b00001110110: data <= 32'h394a3e59;
    11'b00001110111: data <= 32'h34e54215;
    11'b00001111000: data <= 32'hb687400a;
    11'b00001111001: data <= 32'hb6761f6c;
    11'b00001111010: data <= 32'ha81ab89f;
    11'b00001111011: data <= 32'hb0bd3409;
    11'b00001111100: data <= 32'hb3633815;
    11'b00001111101: data <= 32'h3ae1b7a3;
    11'b00001111110: data <= 32'h4105bcc2;
    11'b00001111111: data <= 32'h4137b830;
    11'b00010000000: data <= 32'h38e237f8;
    11'b00010000001: data <= 32'hbd3a37be;
    11'b00010000010: data <= 32'hbcb4b446;
    11'b00010000011: data <= 32'h2a71b973;
    11'b00010000100: data <= 32'h3032bac0;
    11'b00010000101: data <= 32'hbc21bdda;
    11'b00010000110: data <= 32'hbdc6bfeb;
    11'b00010000111: data <= 32'hb455bc1f;
    11'b00010001000: data <= 32'h3aee3c58;
    11'b00010001001: data <= 32'h36e84069;
    11'b00010001010: data <= 32'hbace3d01;
    11'b00010001011: data <= 32'hbd90ae4a;
    11'b00010001100: data <= 32'hbc442ff9;
    11'b00010001101: data <= 32'hba1d3cfe;
    11'b00010001110: data <= 32'hb6e03c7f;
    11'b00010001111: data <= 32'h3987b6b7;
    11'b00010010000: data <= 32'h4036bcef;
    11'b00010010001: data <= 32'h4069af63;
    11'b00010010010: data <= 32'h39f43db1;
    11'b00010010011: data <= 32'hb67a3dce;
    11'b00010010100: data <= 32'h2d2d332e;
    11'b00010010101: data <= 32'h3b90b9de;
    11'b00010010110: data <= 32'h3567bc45;
    11'b00010010111: data <= 32'hbc9abe0e;
    11'b00010011000: data <= 32'hbd0dbfcf;
    11'b00010011001: data <= 32'h3696bd7c;
    11'b00010011010: data <= 32'h3e8a2e84;
    11'b00010011011: data <= 32'h39b13b05;
    11'b00010011100: data <= 32'hbcd0343e;
    11'b00010011101: data <= 32'hc002b4fa;
    11'b00010011110: data <= 32'hbe08370e;
    11'b00010011111: data <= 32'hbc0d3dc4;
    11'b00010100000: data <= 32'hbae53aa1;
    11'b00010100001: data <= 32'hb341bb44;
    11'b00010100010: data <= 32'h3b3dbd3d;
    11'b00010100011: data <= 32'h3d55379c;
    11'b00010100100: data <= 32'h396440ae;
    11'b00010100101: data <= 32'h31db4055;
    11'b00010100110: data <= 32'h398c38bc;
    11'b00010100111: data <= 32'h3c5ab624;
    11'b00010101000: data <= 32'h30a0b61c;
    11'b00010101001: data <= 32'hbc64b8c1;
    11'b00010101010: data <= 32'hb8b8bd5e;
    11'b00010101011: data <= 32'h3dd5be2f;
    11'b00010101100: data <= 32'h40f1ba36;
    11'b00010101101: data <= 32'h3c32ae96;
    11'b00010101110: data <= 32'hbc64b3e2;
    11'b00010101111: data <= 32'hbecdb581;
    11'b00010110000: data <= 32'hbbca35f0;
    11'b00010110001: data <= 32'hb9b73afe;
    11'b00010110010: data <= 32'hbd26b021;
    11'b00010110011: data <= 32'hbd61bec5;
    11'b00010110100: data <= 32'hb536be0a;
    11'b00010110101: data <= 32'h38df3996;
    11'b00010110110: data <= 32'h388240fe;
    11'b00010110111: data <= 32'h3379401d;
    11'b00010111000: data <= 32'h36473891;
    11'b00010111001: data <= 32'h367e3217;
    11'b00010111010: data <= 32'hb6f83aba;
    11'b00010111011: data <= 32'hbc6739d6;
    11'b00010111100: data <= 32'hab50b8aa;
    11'b00010111101: data <= 32'h4015be23;
    11'b00010111110: data <= 32'h4180bc5a;
    11'b00010111111: data <= 32'h3cdeb198;
    11'b00011000000: data <= 32'hb8512c14;
    11'b00011000001: data <= 32'hb899a982;
    11'b00011000010: data <= 32'h343031a1;
    11'b00011000011: data <= 32'hac69300a;
    11'b00011000100: data <= 32'hbe01bbf5;
    11'b00011000101: data <= 32'hc009c074;
    11'b00011000110: data <= 32'hba8ebefb;
    11'b00011000111: data <= 32'h38683506;
    11'b00011001000: data <= 32'h38fc3eae;
    11'b00011001001: data <= 32'had643c5d;
    11'b00011001010: data <= 32'hb6e6307e;
    11'b00011001011: data <= 32'hb863394c;
    11'b00011001100: data <= 32'hbc253f83;
    11'b00011001101: data <= 32'hbd0c3e7c;
    11'b00011001110: data <= 32'hb0e2b362;
    11'b00011001111: data <= 32'h3e90bdeb;
    11'b00011010000: data <= 32'h405aba6c;
    11'b00011010001: data <= 32'h3c353876;
    11'b00011010010: data <= 32'h30633b67;
    11'b00011010011: data <= 32'h39b93727;
    11'b00011010100: data <= 32'h3dc1304f;
    11'b00011010101: data <= 32'h3757b00e;
    11'b00011010110: data <= 32'hbdf4bc2d;
    11'b00011010111: data <= 32'hbfcfc020;
    11'b00011011000: data <= 32'hb5a8bf4d;
    11'b00011011001: data <= 32'h3cbbb756;
    11'b00011011010: data <= 32'h3b38350a;
    11'b00011011011: data <= 32'hb631b1a5;
    11'b00011011100: data <= 32'hbc1fb6a1;
    11'b00011011101: data <= 32'hbbdc3a8c;
    11'b00011011110: data <= 32'hbcbd405a;
    11'b00011011111: data <= 32'hbdec3e42;
    11'b00011100000: data <= 32'hbb0db866;
    11'b00011100001: data <= 32'h36afbe2e;
    11'b00011100010: data <= 32'h3c1eb4a0;
    11'b00011100011: data <= 32'h39043daf;
    11'b00011100100: data <= 32'h38533e7f;
    11'b00011100101: data <= 32'h3db239ff;
    11'b00011100110: data <= 32'h3f5e3532;
    11'b00011100111: data <= 32'h378d3669;
    11'b00011101000: data <= 32'hbd9faf00;
    11'b00011101001: data <= 32'hbd7ebcca;
    11'b00011101010: data <= 32'h38d7be96;
    11'b00011101011: data <= 32'h3ff6bc8b;
    11'b00011101100: data <= 32'h3cd2ba08;
    11'b00011101101: data <= 32'hb637bbc5;
    11'b00011101110: data <= 32'hbaceb98d;
    11'b00011101111: data <= 32'hb704398f;
    11'b00011110000: data <= 32'hb9463edb;
    11'b00011110001: data <= 32'hbe4739d1;
    11'b00011110010: data <= 32'hbf2bbd27;
    11'b00011110011: data <= 32'hbb27beee;
    11'b00011110100: data <= 32'h1c5f9f8c;
    11'b00011110101: data <= 32'h335d3eac;
    11'b00011110110: data <= 32'h38113e0c;
    11'b00011110111: data <= 32'h3cf1384a;
    11'b00011111000: data <= 32'h3d4138bc;
    11'b00011111001: data <= 32'ha8e03dae;
    11'b00011111010: data <= 32'hbda33d27;
    11'b00011111011: data <= 32'hba94b00c;
    11'b00011111100: data <= 32'h3cfcbd41;
    11'b00011111101: data <= 32'h408abd57;
    11'b00011111110: data <= 32'h3ce0bb8c;
    11'b00011111111: data <= 32'hae39bad0;
    11'b00100000000: data <= 32'h2d6cb7f1;
    11'b00100000001: data <= 32'h3ae73805;
    11'b00100000010: data <= 32'h34c43bdc;
    11'b00100000011: data <= 32'hbdc2b14a;
    11'b00100000100: data <= 32'hc0a6bf52;
    11'b00100000101: data <= 32'hbe07bf6a;
    11'b00100000110: data <= 32'hb482b15c;
    11'b00100000111: data <= 32'h309e3c0e;
    11'b00100001000: data <= 32'h31ea37cd;
    11'b00100001001: data <= 32'h3753b23c;
    11'b00100001010: data <= 32'h35da39b4;
    11'b00100001011: data <= 32'hb92e4099;
    11'b00100001100: data <= 32'hbdfb4099;
    11'b00100001101: data <= 32'hb9e937cf;
    11'b00100001110: data <= 32'h3c00bc46;
    11'b00100001111: data <= 32'h3e9bbc19;
    11'b00100010000: data <= 32'h3a30b477;
    11'b00100010001: data <= 32'h3370a83d;
    11'b00100010010: data <= 32'h3cd49e3e;
    11'b00100010011: data <= 32'h405236b5;
    11'b00100010100: data <= 32'h3c7838c3;
    11'b00100010101: data <= 32'hbcc4b59c;
    11'b00100010110: data <= 32'hc06cbe8d;
    11'b00100010111: data <= 32'hbc82bebb;
    11'b00100011000: data <= 32'h3448b8dd;
    11'b00100011001: data <= 32'h3678b175;
    11'b00100011010: data <= 32'hb065bb37;
    11'b00100011011: data <= 32'hb376bc42;
    11'b00100011100: data <= 32'hb1e138c2;
    11'b00100011101: data <= 32'hba4d410d;
    11'b00100011110: data <= 32'hbe0340b1;
    11'b00100011111: data <= 32'hbca334b3;
    11'b00100100000: data <= 32'haabdbc56;
    11'b00100100001: data <= 32'h3638b803;
    11'b00100100010: data <= 32'h24d2391b;
    11'b00100100011: data <= 32'h354c3a0e;
    11'b00100100100: data <= 32'h3f4e34e8;
    11'b00100100101: data <= 32'h415d3711;
    11'b00100100110: data <= 32'h3d333ac9;
    11'b00100100111: data <= 32'hbc1636a7;
    11'b00100101000: data <= 32'hbe7db956;
    11'b00100101001: data <= 32'hb0b1bcb0;
    11'b00100101010: data <= 32'h3c8ebbac;
    11'b00100101011: data <= 32'h39d1bc89;
    11'b00100101100: data <= 32'hb43cbf54;
    11'b00100101101: data <= 32'hb4a4be3d;
    11'b00100101110: data <= 32'h324d357a;
    11'b00100101111: data <= 32'hb1a44018;
    11'b00100110000: data <= 32'hbd153e0e;
    11'b00100110001: data <= 32'hbef0b7a5;
    11'b00100110010: data <= 32'hbcfcbd2b;
    11'b00100110011: data <= 32'hba4bb01f;
    11'b00100110100: data <= 32'hb91c3c56;
    11'b00100110101: data <= 32'h30033a68;
    11'b00100110110: data <= 32'h3e7327df;
    11'b00100110111: data <= 32'h406136a1;
    11'b00100111000: data <= 32'h3a593e22;
    11'b00100111001: data <= 32'hbc263ebe;
    11'b00100111010: data <= 32'hbc07387e;
    11'b00100111011: data <= 32'h3946b853;
    11'b00100111100: data <= 32'h3e45bb87;
    11'b00100111101: data <= 32'h39a0bd25;
    11'b00100111110: data <= 32'hb380bf1e;
    11'b00100111111: data <= 32'h3536bda4;
    11'b00101000000: data <= 32'h3d753093;
    11'b00101000001: data <= 32'h3b813d15;
    11'b00101000010: data <= 32'hba8937d1;
    11'b00101000011: data <= 32'hc006bca2;
    11'b00101000100: data <= 32'hbf3dbd99;
    11'b00101000101: data <= 32'hbcb0ac24;
    11'b00101000110: data <= 32'hba9939d6;
    11'b00101000111: data <= 32'hb384ad5e;
    11'b00101001000: data <= 32'h3a69bacc;
    11'b00101001001: data <= 32'h3c91325f;
    11'b00101001010: data <= 32'h2bac4043;
    11'b00101001011: data <= 32'hbc864146;
    11'b00101001100: data <= 32'hb9e33d37;
    11'b00101001101: data <= 32'h3988b076;
    11'b00101001110: data <= 32'h3c5fb871;
    11'b00101001111: data <= 32'h2ff3b8c3;
    11'b00101010000: data <= 32'hb3aabb2a;
    11'b00101010001: data <= 32'h3c9aba8e;
    11'b00101010010: data <= 32'h412f2d2d;
    11'b00101010011: data <= 32'h3fa439db;
    11'b00101010100: data <= 32'hb5c52a0e;
    11'b00101010101: data <= 32'hbf1fbc79;
    11'b00101010110: data <= 32'hbd9ebc79;
    11'b00101010111: data <= 32'hb8c2b1d4;
    11'b00101011000: data <= 32'hb7f8b0c5;
    11'b00101011001: data <= 32'hb844bd97;
    11'b00101011010: data <= 32'ha126bf91;
    11'b00101011011: data <= 32'h35c3b183;
    11'b00101011100: data <= 32'hb3bb4066;
    11'b00101011101: data <= 32'hbc3b414f;
    11'b00101011110: data <= 32'hbad73c7c;
    11'b00101011111: data <= 32'haaeeb1b0;
    11'b00101100000: data <= 32'had8ea9b2;
    11'b00101100001: data <= 32'hba8436ad;
    11'b00101100010: data <= 32'hb6e32e57;
    11'b00101100011: data <= 32'h3e4eb577;
    11'b00101100100: data <= 32'h422c2b10;
    11'b00101100101: data <= 32'h404a39b0;
    11'b00101100110: data <= 32'hb1363813;
    11'b00101100111: data <= 32'hbcbbb3c6;
    11'b00101101000: data <= 32'hb588b6c2;
    11'b00101101001: data <= 32'h3739b2f9;
    11'b00101101010: data <= 32'ha3bfbb23;
    11'b00101101011: data <= 32'hb973c09b;
    11'b00101101100: data <= 32'hb4edc0f5;
    11'b00101101101: data <= 32'h3717b80f;
    11'b00101101110: data <= 32'h341e3ebc;
    11'b00101101111: data <= 32'hb9383f09;
    11'b00101110000: data <= 32'hbc6732a0;
    11'b00101110001: data <= 32'hbc04b840;
    11'b00101110010: data <= 32'hbcf43546;
    11'b00101110011: data <= 32'hbe6c3c4b;
    11'b00101110100: data <= 32'hba3236e4;
    11'b00101110101: data <= 32'h3d2db7c7;
    11'b00101110110: data <= 32'h4116afea;
    11'b00101110111: data <= 32'h3e213c45;
    11'b00101111000: data <= 32'hb4ca3e12;
    11'b00101111001: data <= 32'hb8973bab;
    11'b00101111010: data <= 32'h39263605;
    11'b00101111011: data <= 32'h3c9fa002;
    11'b00101111100: data <= 32'h2f08bb8d;
    11'b00101111101: data <= 32'hba30c06d;
    11'b00101111110: data <= 32'ha14ac08a;
    11'b00101111111: data <= 32'h3d58b8f5;
    11'b00110000000: data <= 32'h3d583b4f;
    11'b00110000001: data <= 32'ha0653894;
    11'b00110000010: data <= 32'hbc90b9e0;
    11'b00110000011: data <= 32'hbdbeba6a;
    11'b00110000100: data <= 32'hbe6737c9;
    11'b00110000101: data <= 32'hbf203c14;
    11'b00110000110: data <= 32'hbc5fb188;
    11'b00110000111: data <= 32'h37b4bd44;
    11'b00110001000: data <= 32'h3d6bb84d;
    11'b00110001001: data <= 32'h38723d92;
    11'b00110001010: data <= 32'hb883409e;
    11'b00110001011: data <= 32'hb3983ec3;
    11'b00110001100: data <= 32'h3baa3a90;
    11'b00110001101: data <= 32'h3bc0363a;
    11'b00110001110: data <= 32'hb66db38b;
    11'b00110001111: data <= 32'hbbcbbcd9;
    11'b00110010000: data <= 32'h3828bdd8;
    11'b00110010001: data <= 32'h40c3b816;
    11'b00110010010: data <= 32'h409d3550;
    11'b00110010011: data <= 32'h3852b041;
    11'b00110010100: data <= 32'hbab9bbea;
    11'b00110010101: data <= 32'hbbefb8e3;
    11'b00110010110: data <= 32'hbb71386b;
    11'b00110010111: data <= 32'hbd193725;
    11'b00110011000: data <= 32'hbceebd24;
    11'b00110011001: data <= 32'hb5aec0ba;
    11'b00110011010: data <= 32'h3540bc2c;
    11'b00110011011: data <= 32'ha9dd3d5b;
    11'b00110011100: data <= 32'hb8dd4087;
    11'b00110011101: data <= 32'hb22d3dc2;
    11'b00110011110: data <= 32'h382f3930;
    11'b00110011111: data <= 32'h1fe53a25;
    11'b00110100000: data <= 32'hbd623a59;
    11'b00110100001: data <= 32'hbd541f7a;
    11'b00110100010: data <= 32'h3a3ab976;
    11'b00110100011: data <= 32'h4196b64c;
    11'b00110100100: data <= 32'h40fe3189;
    11'b00110100101: data <= 32'h394024b7;
    11'b00110100110: data <= 32'hb55fb5a1;
    11'b00110100111: data <= 32'h2d5a2d54;
    11'b00110101000: data <= 32'h351739a6;
    11'b00110101001: data <= 32'hb7ffadc6;
    11'b00110101010: data <= 32'hbcdfc02d;
    11'b00110101011: data <= 32'hba1dc1dd;
    11'b00110101100: data <= 32'h2eafbd68;
    11'b00110101101: data <= 32'h32343af8;
    11'b00110101110: data <= 32'hb31f3d61;
    11'b00110101111: data <= 32'hb39f3589;
    11'b00110110000: data <= 32'hb20d25bd;
    11'b00110110001: data <= 32'hbc193bc6;
    11'b00110110010: data <= 32'hc0483e26;
    11'b00110110011: data <= 32'hbed1391a;
    11'b00110110100: data <= 32'h37efb860;
    11'b00110110101: data <= 32'h406eb834;
    11'b00110110110: data <= 32'h3eee354d;
    11'b00110110111: data <= 32'h346b3a1c;
    11'b00110111000: data <= 32'h2ecf39b2;
    11'b00110111001: data <= 32'h3c933b3e;
    11'b00110111010: data <= 32'h3d3f3bfa;
    11'b00110111011: data <= 32'hacf3ae11;
    11'b00110111100: data <= 32'hbceebfd4;
    11'b00110111101: data <= 32'hb938c133;
    11'b00110111110: data <= 32'h39bdbd09;
    11'b00110111111: data <= 32'h3c733409;
    11'b00111000000: data <= 32'h37412e3c;
    11'b00111000001: data <= 32'hb0e9bb01;
    11'b00111000010: data <= 32'hb839b876;
    11'b00111000011: data <= 32'hbd5b3c17;
    11'b00111000100: data <= 32'hc0773e9c;
    11'b00111000101: data <= 32'hbf77353a;
    11'b00111000110: data <= 32'hb210bcc6;
    11'b00111000111: data <= 32'h3bc8bbbe;
    11'b00111001000: data <= 32'h37d237f9;
    11'b00111001001: data <= 32'hb4dc3dae;
    11'b00111001010: data <= 32'h35043d8d;
    11'b00111001011: data <= 32'h3e713d36;
    11'b00111001100: data <= 32'h3db53d2d;
    11'b00111001101: data <= 32'hb6093826;
    11'b00111001110: data <= 32'hbdcbbb42;
    11'b00111001111: data <= 32'hb4c9be2e;
    11'b00111010000: data <= 32'h3e5fbab5;
    11'b00111010001: data <= 32'h4008b1dc;
    11'b00111010010: data <= 32'h3bebb9f6;
    11'b00111010011: data <= 32'h2ecabdc3;
    11'b00111010100: data <= 32'hb075b8dc;
    11'b00111010101: data <= 32'hb8fe3c54;
    11'b00111010110: data <= 32'hbe083d0f;
    11'b00111010111: data <= 32'hbed9b8b2;
    11'b00111011000: data <= 32'hbafac051;
    11'b00111011001: data <= 32'hb1b1bdf4;
    11'b00111011010: data <= 32'hb6e836e5;
    11'b00111011011: data <= 32'hb8f13d90;
    11'b00111011100: data <= 32'h35373c60;
    11'b00111011101: data <= 32'h3d733b99;
    11'b00111011110: data <= 32'h39853da5;
    11'b00111011111: data <= 32'hbce43d96;
    11'b00111100000: data <= 32'hbf5b36c8;
    11'b00111100001: data <= 32'hae87b720;
    11'b00111100010: data <= 32'h3feab6c8;
    11'b00111100011: data <= 32'h4055b481;
    11'b00111100100: data <= 32'h3bbcba3d;
    11'b00111100101: data <= 32'h3649bc36;
    11'b00111100110: data <= 32'h3a65a888;
    11'b00111100111: data <= 32'h39cd3d1c;
    11'b00111101000: data <= 32'hb6aa3a9e;
    11'b00111101001: data <= 32'hbd85bd53;
    11'b00111101010: data <= 32'hbcc5c162;
    11'b00111101011: data <= 32'hb8a9becd;
    11'b00111101100: data <= 32'hb77c302b;
    11'b00111101101: data <= 32'hb62c38ad;
    11'b00111101110: data <= 32'h351eadc1;
    11'b00111101111: data <= 32'h3a3e25b3;
    11'b00111110000: data <= 32'hb4093d2a;
    11'b00111110001: data <= 32'hbff0400f;
    11'b00111110010: data <= 32'hc0503cea;
    11'b00111110011: data <= 32'hb44ea083;
    11'b00111110100: data <= 32'h3df5b5d6;
    11'b00111110101: data <= 32'h3d49b0c4;
    11'b00111110110: data <= 32'h34f0b1fb;
    11'b00111110111: data <= 32'h3828af28;
    11'b00111111000: data <= 32'h3ef33a02;
    11'b00111111001: data <= 32'h3f8b3e35;
    11'b00111111010: data <= 32'h353c3a12;
    11'b00111111011: data <= 32'hbca9bd0c;
    11'b00111111100: data <= 32'hbc56c095;
    11'b00111111101: data <= 32'hb068bd72;
    11'b00111111110: data <= 32'h34b5b22e;
    11'b00111111111: data <= 32'h33c8b84f;
    11'b01000000000: data <= 32'h36b4bde4;
    11'b01000000001: data <= 32'h36d7bb27;
    11'b01000000010: data <= 32'hb8d13c50;
    11'b01000000011: data <= 32'hc00d403f;
    11'b01000000100: data <= 32'hc03a3c61;
    11'b01000000101: data <= 32'hb984b769;
    11'b01000000110: data <= 32'h35deb9e8;
    11'b01000000111: data <= 32'hacf5a392;
    11'b01000001000: data <= 32'hb8ec3708;
    11'b01000001001: data <= 32'h36fb3895;
    11'b01000001010: data <= 32'h40513c76;
    11'b01000001011: data <= 32'h405f3ec4;
    11'b01000001100: data <= 32'h34113c95;
    11'b01000001101: data <= 32'hbd20b52d;
    11'b01000001110: data <= 32'hba28bc5d;
    11'b01000001111: data <= 32'h395eb8ca;
    11'b01000010000: data <= 32'h3cb6b521;
    11'b01000010001: data <= 32'h3a15bd47;
    11'b01000010010: data <= 32'h3890c076;
    11'b01000010011: data <= 32'h3914bcd2;
    11'b01000010100: data <= 32'h21dc3c02;
    11'b01000010101: data <= 32'hbcb03f14;
    11'b01000010110: data <= 32'hbe86346d;
    11'b01000010111: data <= 32'hbc3abd84;
    11'b01000011000: data <= 32'hb9acbcfb;
    11'b01000011001: data <= 32'hbccaa4c5;
    11'b01000011010: data <= 32'hbce83859;
    11'b01000011011: data <= 32'h346535e1;
    11'b01000011100: data <= 32'h3fbd3943;
    11'b01000011101: data <= 32'h3e463e07;
    11'b01000011110: data <= 32'hb8133edc;
    11'b01000011111: data <= 32'hbe9f3b64;
    11'b01000100000: data <= 32'hb85932d4;
    11'b01000100001: data <= 32'h3c9530a4;
    11'b01000100010: data <= 32'h3d9bb29b;
    11'b01000100011: data <= 32'h3943bd75;
    11'b01000100100: data <= 32'h38c3bff2;
    11'b01000100101: data <= 32'h3d22ba04;
    11'b01000100110: data <= 32'h3d163cac;
    11'b01000100111: data <= 32'h2fc53d50;
    11'b01000101000: data <= 32'hbb93b821;
    11'b01000101001: data <= 32'hbc85bfdf;
    11'b01000101010: data <= 32'hbc70bd9b;
    11'b01000101011: data <= 32'hbd9cae80;
    11'b01000101100: data <= 32'hbc9f96d4;
    11'b01000101101: data <= 32'h32f7b9d2;
    11'b01000101110: data <= 32'h3d77b769;
    11'b01000101111: data <= 32'h38e73c1b;
    11'b01000110000: data <= 32'hbd3f4026;
    11'b01000110001: data <= 32'hbfc33ed7;
    11'b01000110010: data <= 32'hb84f3abb;
    11'b01000110011: data <= 32'h3b123698;
    11'b01000110100: data <= 32'h39262077;
    11'b01000110101: data <= 32'hb1afba5a;
    11'b01000110110: data <= 32'h35dabc44;
    11'b01000110111: data <= 32'h3fba2af3;
    11'b01000111000: data <= 32'h40ce3db7;
    11'b01000111001: data <= 32'h3c4e3c87;
    11'b01000111010: data <= 32'hb7a3b920;
    11'b01000111011: data <= 32'hbb34be9f;
    11'b01000111100: data <= 32'hb985bb45;
    11'b01000111101: data <= 32'hb994ad8c;
    11'b01000111110: data <= 32'hb848baa9;
    11'b01000111111: data <= 32'h3501c025;
    11'b01001000000: data <= 32'h3b66be6b;
    11'b01001000001: data <= 32'h2e8c3823;
    11'b01001000010: data <= 32'hbdc24003;
    11'b01001000011: data <= 32'hbf163e65;
    11'b01001000100: data <= 32'hb92f37ac;
    11'b01001000101: data <= 32'h29f32d77;
    11'b01001000110: data <= 32'hb9b630c9;
    11'b01001000111: data <= 32'hbd58af3b;
    11'b01001001000: data <= 32'ha9e1b415;
    11'b01001001001: data <= 32'h4051380d;
    11'b01001001010: data <= 32'h41703de7;
    11'b01001001011: data <= 32'h3c853cf9;
    11'b01001001100: data <= 32'hb8012649;
    11'b01001001101: data <= 32'hb881b803;
    11'b01001001110: data <= 32'h30bd2dbe;
    11'b01001001111: data <= 32'h3473305a;
    11'b01001010000: data <= 32'h2c28bd90;
    11'b01001010001: data <= 32'h3677c1b0;
    11'b01001010010: data <= 32'h3b2ec028;
    11'b01001010011: data <= 32'h375c34cc;
    11'b01001010100: data <= 32'hb9253e6b;
    11'b01001010101: data <= 32'hbc403a24;
    11'b01001010110: data <= 32'hb93eb7de;
    11'b01001010111: data <= 32'hba4bb7da;
    11'b01001011000: data <= 32'hbf6431bd;
    11'b01001011001: data <= 32'hc04931da;
    11'b01001011010: data <= 32'hb664b334;
    11'b01001011011: data <= 32'h3f6d2f86;
    11'b01001011100: data <= 32'h40343c59;
    11'b01001011101: data <= 32'h35903dd2;
    11'b01001011110: data <= 32'hbb603c10;
    11'b01001011111: data <= 32'hb51e3a86;
    11'b01001100000: data <= 32'h3a353c3d;
    11'b01001100001: data <= 32'h39b637dc;
    11'b01001100010: data <= 32'h2996bd4e;
    11'b01001100011: data <= 32'h3415c138;
    11'b01001100100: data <= 32'h3cd3be94;
    11'b01001100101: data <= 32'h3dd537b8;
    11'b01001100110: data <= 32'h39443c9b;
    11'b01001100111: data <= 32'hb02bb0ac;
    11'b01001101000: data <= 32'hb716bd14;
    11'b01001101001: data <= 32'hbc32b9ea;
    11'b01001101010: data <= 32'hc0253385;
    11'b01001101011: data <= 32'hc045aa34;
    11'b01001101100: data <= 32'hb7abbc3c;
    11'b01001101101: data <= 32'h3d16bc01;
    11'b01001101110: data <= 32'h3c35358e;
    11'b01001101111: data <= 32'hb8f23dfb;
    11'b01001110000: data <= 32'hbd383e8b;
    11'b01001110001: data <= 32'hb2b73de6;
    11'b01001110010: data <= 32'h3a5f3dc1;
    11'b01001110011: data <= 32'h32c83a37;
    11'b01001110100: data <= 32'hba36b9d4;
    11'b01001110101: data <= 32'hb358be7c;
    11'b01001110110: data <= 32'h3e0fb99f;
    11'b01001110111: data <= 32'h40cc3ab9;
    11'b01001111000: data <= 32'h3e9d3b09;
    11'b01001111001: data <= 32'h37ffb82d;
    11'b01001111010: data <= 32'hadb5bcd3;
    11'b01001111011: data <= 32'hb8a8b472;
    11'b01001111100: data <= 32'hbd4a37da;
    11'b01001111101: data <= 32'hbda9b845;
    11'b01001111110: data <= 32'hb4bac065;
    11'b01001111111: data <= 32'h3a39c060;
    11'b01010000000: data <= 32'h351fb5d2;
    11'b01010000001: data <= 32'hbbe93cff;
    11'b01010000010: data <= 32'hbcbf3dd0;
    11'b01010000011: data <= 32'hae733c5e;
    11'b01010000100: data <= 32'h34d13c39;
    11'b01010000101: data <= 32'hbb6f3ace;
    11'b01010000110: data <= 32'hbfeea212;
    11'b01010000111: data <= 32'hbb01b8f1;
    11'b01010001000: data <= 32'h3e10a3bf;
    11'b01010001001: data <= 32'h413e3baf;
    11'b01010001010: data <= 32'h3ed53a69;
    11'b01010001011: data <= 32'h3788b204;
    11'b01010001100: data <= 32'h32e9b46f;
    11'b01010001101: data <= 32'h34923a1f;
    11'b01010001110: data <= 32'hb1e63bc1;
    11'b01010001111: data <= 32'hb8beba9f;
    11'b01010010000: data <= 32'haf1fc1b5;
    11'b01010010001: data <= 32'h38c1c15e;
    11'b01010010010: data <= 32'h35c8b908;
    11'b01010010011: data <= 32'hb6d23aaf;
    11'b01010010100: data <= 32'hb71c38b7;
    11'b01010010101: data <= 32'h310fa33f;
    11'b01010010110: data <= 32'hb3af347b;
    11'b01010010111: data <= 32'hbfba3a35;
    11'b01010011000: data <= 32'hc1aa3687;
    11'b01010011001: data <= 32'hbd51b4a5;
    11'b01010011010: data <= 32'h3c9db121;
    11'b01010011011: data <= 32'h3fd73878;
    11'b01010011100: data <= 32'h3a8e39fe;
    11'b01010011101: data <= 32'hafa637df;
    11'b01010011110: data <= 32'h35b03b28;
    11'b01010011111: data <= 32'h3c0b3f32;
    11'b01010100000: data <= 32'h38373de7;
    11'b01010100001: data <= 32'hb5cdb93f;
    11'b01010100010: data <= 32'hb3e2c122;
    11'b01010100011: data <= 32'h3938c059;
    11'b01010100100: data <= 32'h3c26b50f;
    11'b01010100101: data <= 32'h39b73792;
    11'b01010100110: data <= 32'h3885b673;
    11'b01010100111: data <= 32'h388abc2e;
    11'b01010101000: data <= 32'hb591b32b;
    11'b01010101001: data <= 32'hc0303a51;
    11'b01010101010: data <= 32'hc1903673;
    11'b01010101011: data <= 32'hbd4dba62;
    11'b01010101100: data <= 32'h3915bc68;
    11'b01010101101: data <= 32'h3abeb42c;
    11'b01010101110: data <= 32'hb60e3873;
    11'b01010101111: data <= 32'hba0d3b52;
    11'b01010110000: data <= 32'h36623dee;
    11'b01010110001: data <= 32'h3ced4058;
    11'b01010110010: data <= 32'h35903eef;
    11'b01010110011: data <= 32'hbbe7adf8;
    11'b01010110100: data <= 32'hba6abe10;
    11'b01010110101: data <= 32'h39aabc18;
    11'b01010110110: data <= 32'h3efc3498;
    11'b01010110111: data <= 32'h3e83348f;
    11'b01010111000: data <= 32'h3ce6bba2;
    11'b01010111001: data <= 32'h3b9ebd32;
    11'b01010111010: data <= 32'h2fce2634;
    11'b01010111011: data <= 32'hbd253c65;
    11'b01010111100: data <= 32'hbf8831b9;
    11'b01010111101: data <= 32'hbb52beb8;
    11'b01010111110: data <= 32'h338fc064;
    11'b01010111111: data <= 32'ha973bc20;
    11'b01011000000: data <= 32'hbc3e3311;
    11'b01011000001: data <= 32'hbaf6397e;
    11'b01011000010: data <= 32'h384d3c2d;
    11'b01011000011: data <= 32'h3bf23e96;
    11'b01011000100: data <= 32'hb8223e71;
    11'b01011000101: data <= 32'hc02c383c;
    11'b01011000110: data <= 32'hbe1db609;
    11'b01011000111: data <= 32'h388aa80b;
    11'b01011001000: data <= 32'h3f843942;
    11'b01011001001: data <= 32'h3e84328d;
    11'b01011001010: data <= 32'h3c61baf2;
    11'b01011001011: data <= 32'h3c6bb94a;
    11'b01011001100: data <= 32'h3b413b92;
    11'b01011001101: data <= 32'ha77f3eae;
    11'b01011001110: data <= 32'hba252c41;
    11'b01011001111: data <= 32'hb774c06a;
    11'b01011010000: data <= 32'h2d02c147;
    11'b01011010001: data <= 32'hb392bcf7;
    11'b01011010010: data <= 32'hba6cadff;
    11'b01011010011: data <= 32'hb44eaf7f;
    11'b01011010100: data <= 32'h3b23b14f;
    11'b01011010101: data <= 32'h395038c6;
    11'b01011010110: data <= 32'hbd703d10;
    11'b01011010111: data <= 32'hc1c63b30;
    11'b01011011000: data <= 32'hbfe2316f;
    11'b01011011001: data <= 32'h33ee307d;
    11'b01011011010: data <= 32'h3cfe36c5;
    11'b01011011011: data <= 32'h392e2c2f;
    11'b01011011100: data <= 32'h3426b6be;
    11'b01011011101: data <= 32'h3bde3529;
    11'b01011011110: data <= 32'h3e413fb7;
    11'b01011011111: data <= 32'h3b144069;
    11'b01011100000: data <= 32'hb2bd3408;
    11'b01011100001: data <= 32'hb672bfac;
    11'b01011100010: data <= 32'h2c63c018;
    11'b01011100011: data <= 32'h3234b9bd;
    11'b01011100100: data <= 32'h2feeb2f7;
    11'b01011100101: data <= 32'h397cbc24;
    11'b01011100110: data <= 32'h3d76bd8a;
    11'b01011100111: data <= 32'h38fbb3a6;
    11'b01011101000: data <= 32'hbdf63c35;
    11'b01011101001: data <= 32'hc1893b7c;
    11'b01011101010: data <= 32'hbf31ada9;
    11'b01011101011: data <= 32'hac2ab87c;
    11'b01011101100: data <= 32'h326cb541;
    11'b01011101101: data <= 32'hb9ccb2ec;
    11'b01011101110: data <= 32'hb9abaf2e;
    11'b01011101111: data <= 32'h3a373acd;
    11'b01011110000: data <= 32'h3f324080;
    11'b01011110001: data <= 32'h3b9f40ae;
    11'b01011110010: data <= 32'hb88e3937;
    11'b01011110011: data <= 32'hbaf3bb6a;
    11'b01011110100: data <= 32'h25fab9e1;
    11'b01011110101: data <= 32'h39fe32b4;
    11'b01011110110: data <= 32'h3b96b089;
    11'b01011110111: data <= 32'h3d3cbe51;
    11'b01011111000: data <= 32'h3eb8bf86;
    11'b01011111001: data <= 32'h3bd5b47c;
    11'b01011111010: data <= 32'hb9d13cf8;
    11'b01011111011: data <= 32'hbee43a7b;
    11'b01011111100: data <= 32'hbc52ba49;
    11'b01011111101: data <= 32'hb24bbe26;
    11'b01011111110: data <= 32'hb94abc4b;
    11'b01011111111: data <= 32'hbe97b843;
    11'b01100000000: data <= 32'hbc8ab47d;
    11'b01100000001: data <= 32'h3a1e3709;
    11'b01100000010: data <= 32'h3e993e67;
    11'b01100000011: data <= 32'h34b23fc3;
    11'b01100000100: data <= 32'hbe183c0e;
    11'b01100000101: data <= 32'hbe4931ac;
    11'b01100000110: data <= 32'hb08637e8;
    11'b01100000111: data <= 32'h3b1d3b4e;
    11'b01100001000: data <= 32'h3baaa8f8;
    11'b01100001001: data <= 32'h3c52be43;
    11'b01100001010: data <= 32'h3e62bddb;
    11'b01100001011: data <= 32'h3e193779;
    11'b01100001100: data <= 32'h37d63f23;
    11'b01100001101: data <= 32'hb6093a08;
    11'b01100001110: data <= 32'hb482bd19;
    11'b01100001111: data <= 32'hb07ebfe0;
    11'b01100010000: data <= 32'hbb48bcd7;
    11'b01100010001: data <= 32'hbe7fb948;
    11'b01100010010: data <= 32'hb9e9bb05;
    11'b01100010011: data <= 32'h3c4cb9d7;
    11'b01100010100: data <= 32'h3d973551;
    11'b01100010101: data <= 32'hb7863cf7;
    11'b01100010110: data <= 32'hc0953c93;
    11'b01100010111: data <= 32'hbfdc3a19;
    11'b01100011000: data <= 32'hb53a3b52;
    11'b01100011001: data <= 32'h36ca3b5b;
    11'b01100011010: data <= 32'h220aaf0e;
    11'b01100011011: data <= 32'h29a5bcd4;
    11'b01100011100: data <= 32'h3c82b8bf;
    11'b01100011101: data <= 32'h3fb53d98;
    11'b01100011110: data <= 32'h3db44095;
    11'b01100011111: data <= 32'h370c3ad9;
    11'b01100100000: data <= 32'h2ba0bc6e;
    11'b01100100001: data <= 32'haa7cbd9e;
    11'b01100100010: data <= 32'hb893b812;
    11'b01100100011: data <= 32'hbabbb759;
    11'b01100100100: data <= 32'h308abe29;
    11'b01100100101: data <= 32'h3e23bfd6;
    11'b01100100110: data <= 32'h3d46ba2a;
    11'b01100100111: data <= 32'hb97339b6;
    11'b01100101000: data <= 32'hc0643c2e;
    11'b01100101001: data <= 32'hbe9238bc;
    11'b01100101010: data <= 32'hb58d3634;
    11'b01100101011: data <= 32'hb60f3457;
    11'b01100101100: data <= 32'hbd74b629;
    11'b01100101101: data <= 32'hbcc5bb37;
    11'b01100101110: data <= 32'h38a5a67f;
    11'b01100101111: data <= 32'h3ff73ef4;
    11'b01100110000: data <= 32'h3e4a409f;
    11'b01100110001: data <= 32'h34883c04;
    11'b01100110010: data <= 32'hb43fb572;
    11'b01100110011: data <= 32'had43aded;
    11'b01100110100: data <= 32'haabd3978;
    11'b01100110101: data <= 32'ha3fea6d7;
    11'b01100110110: data <= 32'h3a38bf8a;
    11'b01100110111: data <= 32'h3f14c10c;
    11'b01100111000: data <= 32'h3de2bc28;
    11'b01100111001: data <= 32'haf8939c6;
    11'b01100111010: data <= 32'hbc9d3b18;
    11'b01100111011: data <= 32'hb95caa29;
    11'b01100111100: data <= 32'haf7cb86b;
    11'b01100111101: data <= 32'hbc18b79c;
    11'b01100111110: data <= 32'hc0b2b93b;
    11'b01100111111: data <= 32'hbf7bbb55;
    11'b01101000000: data <= 32'h357eb43c;
    11'b01101000001: data <= 32'h3f213c65;
    11'b01101000010: data <= 32'h3bdd3eb4;
    11'b01101000011: data <= 32'hb8c93c0c;
    11'b01101000100: data <= 32'hbb9e384c;
    11'b01101000101: data <= 32'hb32a3cc8;
    11'b01101000110: data <= 32'h32243ea5;
    11'b01101000111: data <= 32'h3047357e;
    11'b01101001000: data <= 32'h388bbf21;
    11'b01101001001: data <= 32'h3dedc05e;
    11'b01101001010: data <= 32'h3ebab663;
    11'b01101001011: data <= 32'h3af73ce2;
    11'b01101001100: data <= 32'h33e53a90;
    11'b01101001101: data <= 32'h36bab8ca;
    11'b01101001110: data <= 32'h33d3bc5c;
    11'b01101001111: data <= 32'hbc9eb91b;
    11'b01101010000: data <= 32'hc0d0b8ee;
    11'b01101010001: data <= 32'hbe78bcd9;
    11'b01101010010: data <= 32'h38a0bcd9;
    11'b01101010011: data <= 32'h3e16b2f0;
    11'b01101010100: data <= 32'h32253967;
    11'b01101010101: data <= 32'hbdc33a70;
    11'b01101010110: data <= 32'hbd813bce;
    11'b01101010111: data <= 32'hb4893ed1;
    11'b01101011000: data <= 32'ha2763f66;
    11'b01101011001: data <= 32'hb8d33630;
    11'b01101011010: data <= 32'hb80abda2;
    11'b01101011011: data <= 32'h39bcbd40;
    11'b01101011100: data <= 32'h3eeb389c;
    11'b01101011101: data <= 32'h3e8d3f09;
    11'b01101011110: data <= 32'h3ca13aaa;
    11'b01101011111: data <= 32'h3be0b930;
    11'b01101100000: data <= 32'h37edb9c0;
    11'b01101100001: data <= 32'hba482d87;
    11'b01101100010: data <= 32'hbe98b055;
    11'b01101100011: data <= 32'hb9d0be11;
    11'b01101100100: data <= 32'h3c40c083;
    11'b01101100101: data <= 32'h3d89bdaa;
    11'b01101100110: data <= 32'hb23baf1d;
    11'b01101100111: data <= 32'hbe1337f0;
    11'b01101101000: data <= 32'hbc2e3a07;
    11'b01101101001: data <= 32'haa7e3ce4;
    11'b01101101010: data <= 32'hb77d3ceb;
    11'b01101101011: data <= 32'hbf252e8a;
    11'b01101101100: data <= 32'hbf5abc44;
    11'b01101101101: data <= 32'haf9cb8dc;
    11'b01101101110: data <= 32'h3e273c4a;
    11'b01101101111: data <= 32'h3ed43f26;
    11'b01101110000: data <= 32'h3c433a16;
    11'b01101110001: data <= 32'h39dcb2af;
    11'b01101110010: data <= 32'h37b33664;
    11'b01101110011: data <= 32'hb3ce3d7d;
    11'b01101110100: data <= 32'hb9c538d6;
    11'b01101110101: data <= 32'h2a1bbe46;
    11'b01101110110: data <= 32'h3d4cc171;
    11'b01101110111: data <= 32'h3d6abf12;
    11'b01101111000: data <= 32'h2c4ab337;
    11'b01101111001: data <= 32'hb95b3483;
    11'b01101111010: data <= 32'h22e12e12;
    11'b01101111011: data <= 32'h37ea32de;
    11'b01101111100: data <= 32'hba5b35e2;
    11'b01101111101: data <= 32'hc14eb2a4;
    11'b01101111110: data <= 32'hc13abb82;
    11'b01101111111: data <= 32'hb837b899;
    11'b01110000000: data <= 32'h3ce838ff;
    11'b01110000001: data <= 32'h3c5f3c52;
    11'b01110000010: data <= 32'h30b73752;
    11'b01110000011: data <= 32'ha8f7355d;
    11'b01110000100: data <= 32'h34b53e3a;
    11'b01110000101: data <= 32'h2edb40ee;
    11'b01110000110: data <= 32'hb5533cc4;
    11'b01110000111: data <= 32'h2759bd45;
    11'b01110001000: data <= 32'h3be6c0af;
    11'b01110001001: data <= 32'h3d13bc7a;
    11'b01110001010: data <= 32'h39bd3521;
    11'b01110001011: data <= 32'h38b8340d;
    11'b01110001100: data <= 32'h3cedb845;
    11'b01110001101: data <= 32'h3c75b83b;
    11'b01110001110: data <= 32'hb9db24b8;
    11'b01110001111: data <= 32'hc152b0bc;
    11'b01110010000: data <= 32'hc0c4bbbc;
    11'b01110010001: data <= 32'hb4a1bcc1;
    11'b01110010010: data <= 32'h3be0b853;
    11'b01110010011: data <= 32'h33c1aad7;
    11'b01110010100: data <= 32'hbaf3a959;
    11'b01110010101: data <= 32'hb9203854;
    11'b01110010110: data <= 32'h335d4002;
    11'b01110010111: data <= 32'h30514169;
    11'b01110011000: data <= 32'hb9fd3d20;
    11'b01110011001: data <= 32'hbb12bb76;
    11'b01110011010: data <= 32'h2dfebdb1;
    11'b01110011011: data <= 32'h3c030fa7;
    11'b01110011100: data <= 32'h3cdf3c18;
    11'b01110011101: data <= 32'h3db934a6;
    11'b01110011110: data <= 32'h3f86ba3c;
    11'b01110011111: data <= 32'h3ddeb75c;
    11'b01110100000: data <= 32'hb5113896;
    11'b01110100001: data <= 32'hbf6f3726;
    11'b01110100010: data <= 32'hbd83bb9b;
    11'b01110100011: data <= 32'h3576bfc3;
    11'b01110100100: data <= 32'h3b13bea3;
    11'b01110100101: data <= 32'hb4f0bba5;
    11'b01110100110: data <= 32'hbcebb812;
    11'b01110100111: data <= 32'hb7d2336a;
    11'b01110101000: data <= 32'h386f3dee;
    11'b01110101001: data <= 32'h9fc34003;
    11'b01110101010: data <= 32'hbe813b09;
    11'b01110101011: data <= 32'hc040b910;
    11'b01110101100: data <= 32'hbb0bb8a5;
    11'b01110101101: data <= 32'h38ce3a14;
    11'b01110101110: data <= 32'h3ca13cf4;
    11'b01110101111: data <= 32'h3d3230ec;
    11'b01110110000: data <= 32'h3e5db916;
    11'b01110110001: data <= 32'h3d803591;
    11'b01110110010: data <= 32'h320c3f08;
    11'b01110110011: data <= 32'hba8a3d5b;
    11'b01110110100: data <= 32'hb5c6b9ff;
    11'b01110110101: data <= 32'h3a61c078;
    11'b01110110110: data <= 32'h3a8abfe2;
    11'b01110110111: data <= 32'hb520bc4c;
    11'b01110111000: data <= 32'hb987b991;
    11'b01110111001: data <= 32'h3752b68c;
    11'b01110111010: data <= 32'h3d063614;
    11'b01110111011: data <= 32'haa933b69;
    11'b01110111100: data <= 32'hc09435f6;
    11'b01110111101: data <= 32'hc1b9b7f0;
    11'b01110111110: data <= 32'hbd58b4cc;
    11'b01110111111: data <= 32'h342538f9;
    11'b01111000000: data <= 32'h38413948;
    11'b01111000001: data <= 32'h34d2b4cc;
    11'b01111000010: data <= 32'h390db646;
    11'b01111000011: data <= 32'h3bfe3d1a;
    11'b01111000100: data <= 32'h3835419e;
    11'b01111000101: data <= 32'hb2a24006;
    11'b01111000110: data <= 32'hac9bb691;
    11'b01111000111: data <= 32'h38dfbf41;
    11'b01111001000: data <= 32'h38cbbd04;
    11'b01111001001: data <= 32'h258bb60b;
    11'b01111001010: data <= 32'h351bb874;
    11'b01111001011: data <= 32'h3e88bc0b;
    11'b01111001100: data <= 32'h3ffeb879;
    11'b01111001101: data <= 32'h30e43464;
    11'b01111001110: data <= 32'hc070342d;
    11'b01111001111: data <= 32'hc125b6a5;
    11'b01111010000: data <= 32'hbbeab8da;
    11'b01111010001: data <= 32'h30d4b46e;
    11'b01111010010: data <= 32'hb4a8b6d0;
    11'b01111010011: data <= 32'hbb1abb99;
    11'b01111010100: data <= 32'hb433b604;
    11'b01111010101: data <= 32'h39f53e75;
    11'b01111010110: data <= 32'h390f4203;
    11'b01111010111: data <= 32'hb53b4014;
    11'b01111011000: data <= 32'hb99faf83;
    11'b01111011001: data <= 32'hb328bb4a;
    11'b01111011010: data <= 32'h314e24d2;
    11'b01111011011: data <= 32'h34a938d0;
    11'b01111011100: data <= 32'h3c17b515;
    11'b01111011101: data <= 32'h4081bd39;
    11'b01111011110: data <= 32'h40adba2b;
    11'b01111011111: data <= 32'h38363847;
    11'b01111100000: data <= 32'hbdad3a31;
    11'b01111100001: data <= 32'hbdbbb35a;
    11'b01111100010: data <= 32'haea3bc64;
    11'b01111100011: data <= 32'h3414bcee;
    11'b01111100100: data <= 32'hbaf3bd3f;
    11'b01111100101: data <= 32'hbe0dbdd4;
    11'b01111100110: data <= 32'hb6a3b996;
    11'b01111100111: data <= 32'h3bb03c4e;
    11'b01111101000: data <= 32'h39314062;
    11'b01111101001: data <= 32'hbb663da7;
    11'b01111101010: data <= 32'hbf08a28d;
    11'b01111101011: data <= 32'hbcc1ab50;
    11'b01111101100: data <= 32'hb52f3c1c;
    11'b01111101101: data <= 32'h31353c85;
    11'b01111101110: data <= 32'h3ad4b51f;
    11'b01111101111: data <= 32'h3f7cbd36;
    11'b01111110000: data <= 32'h401fb404;
    11'b01111110001: data <= 32'h3adb3e0a;
    11'b01111110010: data <= 32'hb5ff3e9f;
    11'b01111110011: data <= 32'hb1bf2e2a;
    11'b01111110100: data <= 32'h395ebd17;
    11'b01111110101: data <= 32'h3592bdef;
    11'b01111110110: data <= 32'hbbffbd76;
    11'b01111110111: data <= 32'hbd10be0a;
    11'b01111111000: data <= 32'h34d0bcc9;
    11'b01111111001: data <= 32'h3e93a6ed;
    11'b01111111010: data <= 32'h3a0a3b23;
    11'b01111111011: data <= 32'hbdb238b3;
    11'b01111111100: data <= 32'hc0d2ab86;
    11'b01111111101: data <= 32'hbe6a3520;
    11'b01111111110: data <= 32'hb8b33cba;
    11'b01111111111: data <= 32'hb5cf3a6e;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    