
module memory_rom_6(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbe01b829;
    11'b00000000001: data <= 32'hba48b3a3;
    11'b00000000010: data <= 32'h3b74365f;
    11'b00000000011: data <= 32'h3cf23da4;
    11'b00000000100: data <= 32'hb86c3e99;
    11'b00000000101: data <= 32'hc0753a78;
    11'b00000000110: data <= 32'hbf1031c3;
    11'b00000000111: data <= 32'h24e6389d;
    11'b00000001000: data <= 32'h3c213b0d;
    11'b00000001001: data <= 32'h3b6dacf3;
    11'b00000001010: data <= 32'h3bb3bcfb;
    11'b00000001011: data <= 32'h3df8b96e;
    11'b00000001100: data <= 32'h3de63d1d;
    11'b00000001101: data <= 32'h3843401f;
    11'b00000001110: data <= 32'hb374372a;
    11'b00000001111: data <= 32'haf55bec3;
    11'b00000010000: data <= 32'h2082c02f;
    11'b00000010001: data <= 32'hb90ebc6c;
    11'b00000010010: data <= 32'hbc33b8f4;
    11'b00000010011: data <= 32'ha9bbbc03;
    11'b00000010100: data <= 32'h3d92bb47;
    11'b00000010101: data <= 32'h3c3d31d7;
    11'b00000010110: data <= 32'hbc903c54;
    11'b00000010111: data <= 32'hc16b3b66;
    11'b00000011000: data <= 32'hbfc93776;
    11'b00000011001: data <= 32'hb2bd3830;
    11'b00000011010: data <= 32'h34b337f0;
    11'b00000011011: data <= 32'hb4cbb4d6;
    11'b00000011100: data <= 32'hb18ebb10;
    11'b00000011101: data <= 32'h3c45312a;
    11'b00000011110: data <= 32'h3f5f4025;
    11'b00000011111: data <= 32'h3cc340ed;
    11'b00000100000: data <= 32'h30593958;
    11'b00000100001: data <= 32'hb090bcac;
    11'b00000100010: data <= 32'h9d0bbc90;
    11'b00000100011: data <= 32'hb1a8b29d;
    11'b00000100100: data <= 32'hb03fb6c1;
    11'b00000100101: data <= 32'h3ae6bead;
    11'b00000100110: data <= 32'h3f6cbfc8;
    11'b00000100111: data <= 32'h3c96b87b;
    11'b00000101000: data <= 32'hbbbf3ace;
    11'b00000101001: data <= 32'hc05e3ac8;
    11'b00000101010: data <= 32'hbd8d2baf;
    11'b00000101011: data <= 32'hb3fcb4ad;
    11'b00000101100: data <= 32'hb8d3b526;
    11'b00000101101: data <= 32'hbe7bb946;
    11'b00000101110: data <= 32'hbcbab9f5;
    11'b00000101111: data <= 32'h39be3628;
    11'b00000110000: data <= 32'h3f644008;
    11'b00000110001: data <= 32'h3c06408b;
    11'b00000110010: data <= 32'hb6c43b22;
    11'b00000110011: data <= 32'hb9d9b1f7;
    11'b00000110100: data <= 32'hb0a53478;
    11'b00000110101: data <= 32'h335b3b3b;
    11'b00000110110: data <= 32'h3739ae29;
    11'b00000110111: data <= 32'h3ccfbfa2;
    11'b00000111000: data <= 32'h3fd3c046;
    11'b00000111001: data <= 32'h3dd1b603;
    11'b00000111010: data <= 32'hacab3c9d;
    11'b00000111011: data <= 32'hbb143a22;
    11'b00000111100: data <= 32'hb5e4b899;
    11'b00000111101: data <= 32'hac48bc8f;
    11'b00000111110: data <= 32'hbc9abb4a;
    11'b00000111111: data <= 32'hc086bb25;
    11'b00001000000: data <= 32'hbdb4bbe9;
    11'b00001000001: data <= 32'h39ffb459;
    11'b00001000010: data <= 32'h3e903c11;
    11'b00001000011: data <= 32'h34803e08;
    11'b00001000100: data <= 32'hbd883b7d;
    11'b00001000101: data <= 32'hbd9e3946;
    11'b00001000110: data <= 32'hb5633d4b;
    11'b00001000111: data <= 32'h328f3e20;
    11'b00001001000: data <= 32'h30e72c91;
    11'b00001001001: data <= 32'h38c6bedf;
    11'b00001001010: data <= 32'h3e17be19;
    11'b00001001011: data <= 32'h3ef93806;
    11'b00001001100: data <= 32'h3bf93f0a;
    11'b00001001101: data <= 32'h36af3a5a;
    11'b00001001110: data <= 32'h37f6baff;
    11'b00001001111: data <= 32'h31aabd13;
    11'b00001010000: data <= 32'hbc7ab9ad;
    11'b00001010001: data <= 32'hbfcaba01;
    11'b00001010010: data <= 32'hba8ebdc9;
    11'b00001010011: data <= 32'h3cabbdc1;
    11'b00001010100: data <= 32'h3ddbb5cb;
    11'b00001010101: data <= 32'hb57c38d2;
    11'b00001010110: data <= 32'hbfb03a31;
    11'b00001010111: data <= 32'hbe353b36;
    11'b00001011000: data <= 32'hb5e43db0;
    11'b00001011001: data <= 32'hb42a3d47;
    11'b00001011010: data <= 32'hbb7fad76;
    11'b00001011011: data <= 32'hb974bd7a;
    11'b00001011100: data <= 32'h3a03b97b;
    11'b00001011101: data <= 32'h3f383d53;
    11'b00001011110: data <= 32'h3e5b4049;
    11'b00001011111: data <= 32'h3b9e3ae3;
    11'b00001100000: data <= 32'h397bb8b0;
    11'b00001100001: data <= 32'h3441b721;
    11'b00001100010: data <= 32'hb9733517;
    11'b00001100011: data <= 32'hbc42b2d3;
    11'b00001100100: data <= 32'h2e36bf2a;
    11'b00001100101: data <= 32'h3e7fc0c8;
    11'b00001100110: data <= 32'h3dc4bd20;
    11'b00001100111: data <= 32'hb5d42f2e;
    11'b00001101000: data <= 32'hbe0f386b;
    11'b00001101001: data <= 32'hbb0e380f;
    11'b00001101010: data <= 32'had69395f;
    11'b00001101011: data <= 32'hbaad382f;
    11'b00001101100: data <= 32'hc054b711;
    11'b00001101101: data <= 32'hbf7fbca3;
    11'b00001101110: data <= 32'h2ec9b4ec;
    11'b00001101111: data <= 32'h3e7d3d8a;
    11'b00001110000: data <= 32'h3d9e3f74;
    11'b00001110001: data <= 32'h37cd3a51;
    11'b00001110010: data <= 32'h31032d3f;
    11'b00001110011: data <= 32'h30443b02;
    11'b00001110100: data <= 32'hb38c3e79;
    11'b00001110101: data <= 32'hb5da3704;
    11'b00001110110: data <= 32'h384dbf36;
    11'b00001110111: data <= 32'h3ea7c123;
    11'b00001111000: data <= 32'h3df5bcdf;
    11'b00001111001: data <= 32'h338734f9;
    11'b00001111010: data <= 32'hb511371b;
    11'b00001111011: data <= 32'h353cb09c;
    11'b00001111100: data <= 32'h371cb40a;
    11'b00001111101: data <= 32'hbc7eb0f1;
    11'b00001111110: data <= 32'hc18fb921;
    11'b00001111111: data <= 32'hc087bcc1;
    11'b00010000000: data <= 32'ha2ddb989;
    11'b00010000001: data <= 32'h3d6e37d6;
    11'b00010000010: data <= 32'h39653b5b;
    11'b00010000011: data <= 32'hb81a37a7;
    11'b00010000100: data <= 32'hb8b0392c;
    11'b00010000101: data <= 32'ha9e83f8a;
    11'b00010000110: data <= 32'hadc440d6;
    11'b00010000111: data <= 32'hb6b93a73;
    11'b00010001000: data <= 32'h295fbe14;
    11'b00010001001: data <= 32'h3c46bfd1;
    11'b00010001010: data <= 32'h3db6b552;
    11'b00010001011: data <= 32'h3c0a3bb0;
    11'b00010001100: data <= 32'h3b8d378b;
    11'b00010001101: data <= 32'h3d8eb897;
    11'b00010001110: data <= 32'h3b7db8bf;
    11'b00010001111: data <= 32'hbbb0ac47;
    11'b00010010000: data <= 32'hc0eeb5d7;
    11'b00010010001: data <= 32'hbebebd41;
    11'b00010010010: data <= 32'h36a4be3c;
    11'b00010010011: data <= 32'h3cbabab7;
    11'b00010010100: data <= 32'haa03b269;
    11'b00010010101: data <= 32'hbcef2674;
    11'b00010010110: data <= 32'hbacb39c4;
    11'b00010010111: data <= 32'h26363ff0;
    11'b00010011000: data <= 32'hb40b408b;
    11'b00010011001: data <= 32'hbcdd396e;
    11'b00010011010: data <= 32'hbcb6bca6;
    11'b00010011011: data <= 32'h2cd6bc2c;
    11'b00010011100: data <= 32'h3ca8392d;
    11'b00010011101: data <= 32'h3d993dd6;
    11'b00010011110: data <= 32'h3deb3779;
    11'b00010011111: data <= 32'h3ebbb86b;
    11'b00010100000: data <= 32'h3c69aac4;
    11'b00010100001: data <= 32'hb7f73b25;
    11'b00010100010: data <= 32'hbe1f363c;
    11'b00010100011: data <= 32'hb92fbd40;
    11'b00010100100: data <= 32'h3bdbc090;
    11'b00010100101: data <= 32'h3c76bf09;
    11'b00010100110: data <= 32'hb4cabab4;
    11'b00010100111: data <= 32'hbc5fb543;
    11'b00010101000: data <= 32'hb4223467;
    11'b00010101001: data <= 32'h38163ccc;
    11'b00010101010: data <= 32'hb79f3d8d;
    11'b00010101011: data <= 32'hc063333a;
    11'b00010101100: data <= 32'hc0bdbb73;
    11'b00010101101: data <= 32'hba06b780;
    11'b00010101110: data <= 32'h3a583ba0;
    11'b00010101111: data <= 32'h3c863d16;
    11'b00010110000: data <= 32'h3bf732e2;
    11'b00010110001: data <= 32'h3c6fb34c;
    11'b00010110010: data <= 32'h3b2f3c09;
    11'b00010110011: data <= 32'ha9934061;
    11'b00010110100: data <= 32'hb9553d02;
    11'b00010110101: data <= 32'h27a6bc59;
    11'b00010110110: data <= 32'h3c84c0af;
    11'b00010110111: data <= 32'h3c0cbec0;
    11'b00010111000: data <= 32'ha763b91d;
    11'b00010111001: data <= 32'hb11eb671;
    11'b00010111010: data <= 32'h3b8ab621;
    11'b00010111011: data <= 32'h3d14307f;
    11'b00010111100: data <= 32'hb7ce37e0;
    11'b00010111101: data <= 32'hc153ae23;
    11'b00010111110: data <= 32'hc186babb;
    11'b00010111111: data <= 32'hbb5db85c;
    11'b00011000000: data <= 32'h3821353a;
    11'b00011000001: data <= 32'h36283589;
    11'b00011000010: data <= 32'haf45b55b;
    11'b00011000011: data <= 32'h318b27b5;
    11'b00011000100: data <= 32'h38b73f64;
    11'b00011000101: data <= 32'h32014202;
    11'b00011000110: data <= 32'hb7053edd;
    11'b00011000111: data <= 32'hb240b9ea;
    11'b00011001000: data <= 32'h388ebec5;
    11'b00011001001: data <= 32'h39b8b9bb;
    11'b00011001010: data <= 32'h36b83181;
    11'b00011001011: data <= 32'h3b4bb401;
    11'b00011001100: data <= 32'h4010baf8;
    11'b00011001101: data <= 32'h3f9eb745;
    11'b00011001110: data <= 32'hb2b034f2;
    11'b00011001111: data <= 32'hc0952fbe;
    11'b00011010000: data <= 32'hc03db9fb;
    11'b00011010001: data <= 32'hb5e8bc4f;
    11'b00011010010: data <= 32'h3730ba60;
    11'b00011010011: data <= 32'hb60aba78;
    11'b00011010100: data <= 32'hbc3ebbc9;
    11'b00011010101: data <= 32'hb5b7ac09;
    11'b00011010110: data <= 32'h389b3f7d;
    11'b00011010111: data <= 32'h32f741a2;
    11'b00011011000: data <= 32'hbb373e0a;
    11'b00011011001: data <= 32'hbcc7b76d;
    11'b00011011010: data <= 32'hb753b9fd;
    11'b00011011011: data <= 32'h33713776;
    11'b00011011100: data <= 32'h38c43b70;
    11'b00011011101: data <= 32'h3d69b0c9;
    11'b00011011110: data <= 32'h409fbc0c;
    11'b00011011111: data <= 32'h4017b394;
    11'b00011100000: data <= 32'h32ad3c22;
    11'b00011100001: data <= 32'hbd4d3b34;
    11'b00011100010: data <= 32'hbb38b812;
    11'b00011100011: data <= 32'h371fbe30;
    11'b00011100100: data <= 32'h3806be69;
    11'b00011100101: data <= 32'hba1dbdd6;
    11'b00011100110: data <= 32'hbcedbd6f;
    11'b00011100111: data <= 32'ha2f6b80f;
    11'b00011101000: data <= 32'h3c473c35;
    11'b00011101001: data <= 32'h33923f1e;
    11'b00011101010: data <= 32'hbe663aa5;
    11'b00011101011: data <= 32'hc082b5c5;
    11'b00011101100: data <= 32'hbd4aac19;
    11'b00011101101: data <= 32'hb33b3c47;
    11'b00011101110: data <= 32'h34753c02;
    11'b00011101111: data <= 32'h3a9cb62c;
    11'b00011110000: data <= 32'h3e75bb64;
    11'b00011110001: data <= 32'h3e94383a;
    11'b00011110010: data <= 32'h384d405d;
    11'b00011110011: data <= 32'hb5f43f42;
    11'b00011110100: data <= 32'h2b9bb0a2;
    11'b00011110101: data <= 32'h3ae9be09;
    11'b00011110110: data <= 32'h3711bdea;
    11'b00011110111: data <= 32'hb9b9bcb0;
    11'b00011111000: data <= 32'hb8d6bd1f;
    11'b00011111001: data <= 32'h3c17bc39;
    11'b00011111010: data <= 32'h3f8dad42;
    11'b00011111011: data <= 32'h367538ee;
    11'b00011111100: data <= 32'hbfb23347;
    11'b00011111101: data <= 32'hc12bb575;
    11'b00011111110: data <= 32'hbdbf2c07;
    11'b00011111111: data <= 32'hb6793a0d;
    11'b00100000000: data <= 32'hb62a3422;
    11'b00100000001: data <= 32'hb591bbf5;
    11'b00100000010: data <= 32'h36e8bafd;
    11'b00100000011: data <= 32'h3c363cbe;
    11'b00100000100: data <= 32'h396341d9;
    11'b00100000101: data <= 32'h28c84086;
    11'b00100000110: data <= 32'h30e53129;
    11'b00100000111: data <= 32'h3814bb3e;
    11'b00100001000: data <= 32'h2e24b728;
    11'b00100001001: data <= 32'hb7e3b07d;
    11'b00100001010: data <= 32'h3413bada;
    11'b00100001011: data <= 32'h4010bdba;
    11'b00100001100: data <= 32'h4114bab1;
    11'b00100001101: data <= 32'h39952f2c;
    11'b00100001110: data <= 32'hbe3d32cf;
    11'b00100001111: data <= 32'hbf88b309;
    11'b00100010000: data <= 32'hb991b386;
    11'b00100010001: data <= 32'hb32ab01a;
    11'b00100010010: data <= 32'hbc1fba75;
    11'b00100010011: data <= 32'hbdbebeb9;
    11'b00100010100: data <= 32'hb6aebc25;
    11'b00100010101: data <= 32'h3a433cb3;
    11'b00100010110: data <= 32'h399f415d;
    11'b00100010111: data <= 32'hb22e3f9c;
    11'b00100011000: data <= 32'hb8ab332c;
    11'b00100011001: data <= 32'hb69aac8e;
    11'b00100011010: data <= 32'hb7453ae6;
    11'b00100011011: data <= 32'hb6fb3b72;
    11'b00100011100: data <= 32'h38feb7ab;
    11'b00100011101: data <= 32'h4086be2b;
    11'b00100011110: data <= 32'h4123babd;
    11'b00100011111: data <= 32'h3b94386f;
    11'b00100100000: data <= 32'hb97e3aeb;
    11'b00100100001: data <= 32'hb8632e1e;
    11'b00100100010: data <= 32'h36bcb85d;
    11'b00100100011: data <= 32'h2f85ba9c;
    11'b00100100100: data <= 32'hbd72bda7;
    11'b00100100101: data <= 32'hbf45c000;
    11'b00100100110: data <= 32'hb5fabd75;
    11'b00100100111: data <= 32'h3c7c36d6;
    11'b00100101000: data <= 32'h3a583e28;
    11'b00100101001: data <= 32'hb99f3b7e;
    11'b00100101010: data <= 32'hbe0128d5;
    11'b00100101011: data <= 32'hbcef384f;
    11'b00100101100: data <= 32'hbb283eaa;
    11'b00100101101: data <= 32'hb98d3d45;
    11'b00100101110: data <= 32'h3093b83c;
    11'b00100101111: data <= 32'h3de4be0a;
    11'b00100110000: data <= 32'h3fa3b485;
    11'b00100110001: data <= 32'h3bf73e1f;
    11'b00100110010: data <= 32'h31cb3eed;
    11'b00100110011: data <= 32'h38d837af;
    11'b00100110100: data <= 32'h3cadb814;
    11'b00100110101: data <= 32'h3460b9bf;
    11'b00100110110: data <= 32'hbd65bc33;
    11'b00100110111: data <= 32'hbda0becf;
    11'b00100111000: data <= 32'h376dbe9f;
    11'b00100111001: data <= 32'h3f87b8ee;
    11'b00100111010: data <= 32'h3c093229;
    11'b00100111011: data <= 32'hbbd59fbc;
    11'b00100111100: data <= 32'hbf45b218;
    11'b00100111101: data <= 32'hbd29396f;
    11'b00100111110: data <= 32'hbb313e4c;
    11'b00100111111: data <= 32'hbc8c3a68;
    11'b00101000000: data <= 32'hbb8fbc41;
    11'b00101000001: data <= 32'h2fabbe1b;
    11'b00101000010: data <= 32'h3bcc348e;
    11'b00101000011: data <= 32'h3ade4076;
    11'b00101000100: data <= 32'h38a54045;
    11'b00101000101: data <= 32'h3b67394c;
    11'b00101000110: data <= 32'h3c4aad39;
    11'b00101000111: data <= 32'h26ff33a0;
    11'b00101001000: data <= 32'hbccd3067;
    11'b00101001001: data <= 32'hb95dbb8d;
    11'b00101001010: data <= 32'h3d9ebef9;
    11'b00101001011: data <= 32'h4101bd5c;
    11'b00101001100: data <= 32'h3ce9b853;
    11'b00101001101: data <= 32'hb9edb4fa;
    11'b00101001110: data <= 32'hbcb3b270;
    11'b00101001111: data <= 32'hb6913740;
    11'b00101010000: data <= 32'hb67d3abe;
    11'b00101010001: data <= 32'hbdfab16c;
    11'b00101010010: data <= 32'hbff3bee8;
    11'b00101010011: data <= 32'hbbacbea3;
    11'b00101010100: data <= 32'h362c35a3;
    11'b00101010101: data <= 32'h39be400f;
    11'b00101010110: data <= 32'h36953ea1;
    11'b00101010111: data <= 32'h35dd371b;
    11'b00101011000: data <= 32'h346937a8;
    11'b00101011001: data <= 32'hb8033dfa;
    11'b00101011010: data <= 32'hbc9b3dbe;
    11'b00101011011: data <= 32'hb44eb332;
    11'b00101011100: data <= 32'h3ea6be96;
    11'b00101011101: data <= 32'h40e1bd90;
    11'b00101011110: data <= 32'h3cf2b4bf;
    11'b00101011111: data <= 32'haf9131bb;
    11'b00101100000: data <= 32'h2ec02d43;
    11'b00101100001: data <= 32'h3b6d31ca;
    11'b00101100010: data <= 32'h34aa30fa;
    11'b00101100011: data <= 32'hbe5aba4d;
    11'b00101100100: data <= 32'hc0cabfef;
    11'b00101100101: data <= 32'hbc85bf2d;
    11'b00101100110: data <= 32'h382fb1a4;
    11'b00101100111: data <= 32'h3a073b84;
    11'b00101101000: data <= 32'ha97337ad;
    11'b00101101001: data <= 32'hb802ae80;
    11'b00101101010: data <= 32'hb8523aa6;
    11'b00101101011: data <= 32'hbb3c409f;
    11'b00101101100: data <= 32'hbd13401b;
    11'b00101101101: data <= 32'hb889a868;
    11'b00101101110: data <= 32'h3b63be1e;
    11'b00101101111: data <= 32'h3e57bb24;
    11'b00101110000: data <= 32'h3b7838c1;
    11'b00101110001: data <= 32'h37b53c11;
    11'b00101110010: data <= 32'h3d0d372d;
    11'b00101110011: data <= 32'h3fb02ffe;
    11'b00101110100: data <= 32'h39d12fad;
    11'b00101110101: data <= 32'hbdd2b798;
    11'b00101110110: data <= 32'hc017be10;
    11'b00101110111: data <= 32'hb68bbf04;
    11'b00101111000: data <= 32'h3ce7bb9d;
    11'b00101111001: data <= 32'h3badb675;
    11'b00101111010: data <= 32'hb5dfb9c7;
    11'b00101111011: data <= 32'hbb5cb929;
    11'b00101111100: data <= 32'hb9253a89;
    11'b00101111101: data <= 32'hba30408e;
    11'b00101111110: data <= 32'hbda93ebb;
    11'b00101111111: data <= 32'hbd95b7a3;
    11'b00110000000: data <= 32'hb6b7be22;
    11'b00110000001: data <= 32'h362fb4f8;
    11'b00110000010: data <= 32'h373a3d6f;
    11'b00110000011: data <= 32'h398f3dd9;
    11'b00110000100: data <= 32'h3e8c383d;
    11'b00110000101: data <= 32'h400134d1;
    11'b00110000110: data <= 32'h38e53ab2;
    11'b00110000111: data <= 32'hbd213991;
    11'b00110001000: data <= 32'hbd47b7fc;
    11'b00110001001: data <= 32'h387ebdeb;
    11'b00110001010: data <= 32'h3f87bdd9;
    11'b00110001011: data <= 32'h3c71bcc0;
    11'b00110001100: data <= 32'hb559bcf2;
    11'b00110001101: data <= 32'hb7dfbaaa;
    11'b00110001110: data <= 32'h32ca385d;
    11'b00110001111: data <= 32'ha8b83e4c;
    11'b00110010000: data <= 32'hbda039bb;
    11'b00110010001: data <= 32'hc069bca8;
    11'b00110010010: data <= 32'hbe2dbe7f;
    11'b00110010011: data <= 32'hb71bad45;
    11'b00110010100: data <= 32'h2d6d3d62;
    11'b00110010101: data <= 32'h373b3c11;
    11'b00110010110: data <= 32'h3c7b2df5;
    11'b00110010111: data <= 32'h3cfd380f;
    11'b00110011000: data <= 32'h2d023f69;
    11'b00110011001: data <= 32'hbcd94012;
    11'b00110011010: data <= 32'hba6337c4;
    11'b00110011011: data <= 32'h3bd8bc71;
    11'b00110011100: data <= 32'h3f6fbd9f;
    11'b00110011101: data <= 32'h3b73bbf8;
    11'b00110011110: data <= 32'ha969baa0;
    11'b00110011111: data <= 32'h3865b898;
    11'b00110100000: data <= 32'h3e5a342f;
    11'b00110100001: data <= 32'h3b873a70;
    11'b00110100010: data <= 32'hbcc2a8d1;
    11'b00110100011: data <= 32'hc0f4bde2;
    11'b00110100100: data <= 32'hbf1abe6d;
    11'b00110100101: data <= 32'hb6e6b4f8;
    11'b00110100110: data <= 32'h2b0b37cc;
    11'b00110100111: data <= 32'ha402b224;
    11'b00110101000: data <= 32'h3282b9ea;
    11'b00110101001: data <= 32'h3532382f;
    11'b00110101010: data <= 32'hb61d4103;
    11'b00110101011: data <= 32'hbcdb4170;
    11'b00110101100: data <= 32'hbaa63abf;
    11'b00110101101: data <= 32'h3773bb0a;
    11'b00110101110: data <= 32'h3be0bb0c;
    11'b00110101111: data <= 32'h3586ad46;
    11'b00110110000: data <= 32'h329c2d56;
    11'b00110110001: data <= 32'h3e1bb0d4;
    11'b00110110010: data <= 32'h414f300c;
    11'b00110110011: data <= 32'h3e573856;
    11'b00110110100: data <= 32'hbb282be3;
    11'b00110110101: data <= 32'hc028bc01;
    11'b00110110110: data <= 32'hbc37bd33;
    11'b00110110111: data <= 32'h34edb9da;
    11'b00110111000: data <= 32'h34e7b94f;
    11'b00110111001: data <= 32'hb646bde6;
    11'b00110111010: data <= 32'hb674be1e;
    11'b00110111011: data <= 32'h253b34c8;
    11'b00110111100: data <= 32'hb45140cf;
    11'b00110111101: data <= 32'hbc7d40bc;
    11'b00110111110: data <= 32'hbd41367e;
    11'b00110111111: data <= 32'hb969bb3e;
    11'b00111000000: data <= 32'hb4c2b434;
    11'b00111000001: data <= 32'hb69f3aae;
    11'b00111000010: data <= 32'h314d39b6;
    11'b00111000011: data <= 32'h3f3fa7d7;
    11'b00111000100: data <= 32'h418e2e6f;
    11'b00111000101: data <= 32'h3e163b72;
    11'b00111000110: data <= 32'hb9b13c19;
    11'b00111000111: data <= 32'hbd4a2e06;
    11'b00111001000: data <= 32'h2900b9d5;
    11'b00111001001: data <= 32'h3c84bb9b;
    11'b00111001010: data <= 32'h3817bd5b;
    11'b00111001011: data <= 32'hb831c01b;
    11'b00111001100: data <= 32'hb475bf47;
    11'b00111001101: data <= 32'h3952a5c2;
    11'b00111001110: data <= 32'h383f3ead;
    11'b00111001111: data <= 32'hba7f3d3b;
    11'b00111010000: data <= 32'hbf39b6c8;
    11'b00111010001: data <= 32'hbeb3bc3d;
    11'b00111010010: data <= 32'hbcda2e2f;
    11'b00111010011: data <= 32'hbb7f3c64;
    11'b00111010100: data <= 32'hb18e37af;
    11'b00111010101: data <= 32'h3d07b818;
    11'b00111010110: data <= 32'h3fd4234d;
    11'b00111010111: data <= 32'h3aff3e77;
    11'b00111011000: data <= 32'hb9a34072;
    11'b00111011001: data <= 32'hb9963cb9;
    11'b00111011010: data <= 32'h39a9b0e6;
    11'b00111011011: data <= 32'h3d47b9fe;
    11'b00111011100: data <= 32'h34fcbc66;
    11'b00111011101: data <= 32'hb80abe74;
    11'b00111011110: data <= 32'h36e1bdf3;
    11'b00111011111: data <= 32'h3f8eb40c;
    11'b00111100000: data <= 32'h3e7b3a8b;
    11'b00111100001: data <= 32'hb5903545;
    11'b00111100010: data <= 32'hbf8abb8d;
    11'b00111100011: data <= 32'hbf64bc30;
    11'b00111100100: data <= 32'hbcd12f66;
    11'b00111100101: data <= 32'hbb8c3889;
    11'b00111100110: data <= 32'hb8e1b888;
    11'b00111100111: data <= 32'h3466bdd4;
    11'b00111101000: data <= 32'h3ab2b3e2;
    11'b00111101001: data <= 32'h328c4014;
    11'b00111101010: data <= 32'hb9e541ac;
    11'b00111101011: data <= 32'hb81b3e4e;
    11'b00111101100: data <= 32'h381a2f0c;
    11'b00111101101: data <= 32'h38f2b314;
    11'b00111101110: data <= 32'hb617b030;
    11'b00111101111: data <= 32'hb865b847;
    11'b00111110000: data <= 32'h3c97baef;
    11'b00111110001: data <= 32'h41c1b565;
    11'b00111110010: data <= 32'h40aa35e6;
    11'b00111110011: data <= 32'h28cd2f9b;
    11'b00111110100: data <= 32'hbdc5b94b;
    11'b00111110101: data <= 32'hbc4bb934;
    11'b00111110110: data <= 32'hb54f9ead;
    11'b00111110111: data <= 32'hb826b4d8;
    11'b00111111000: data <= 32'hbb67bf0d;
    11'b00111111001: data <= 32'hb7d6c0b0;
    11'b00111111010: data <= 32'h3390b8eb;
    11'b00111111011: data <= 32'h2f2e3f67;
    11'b00111111100: data <= 32'hb8a440de;
    11'b00111111101: data <= 32'hb99e3c2a;
    11'b00111111110: data <= 32'hb555aae5;
    11'b00111111111: data <= 32'hb88c3568;
    11'b01000000000: data <= 32'hbd0c3b5d;
    11'b01000000001: data <= 32'hba443602;
    11'b01000000010: data <= 32'h3d3ab839;
    11'b01000000011: data <= 32'h41e5b65e;
    11'b01000000100: data <= 32'h406d37ab;
    11'b01000000101: data <= 32'h300c3a33;
    11'b01000000110: data <= 32'hb9da352f;
    11'b01000000111: data <= 32'h30582b31;
    11'b01000001000: data <= 32'h3a00204d;
    11'b01000001001: data <= 32'hada6ba89;
    11'b01000001010: data <= 32'hbc40c097;
    11'b01000001011: data <= 32'hb8f8c13f;
    11'b01000001100: data <= 32'h388bbb25;
    11'b01000001101: data <= 32'h3a473c8d;
    11'b01000001110: data <= 32'hb04d3d15;
    11'b01000001111: data <= 32'hbb72a69e;
    11'b01000010000: data <= 32'hbc8eb6e8;
    11'b01000010001: data <= 32'hbdc4396f;
    11'b01000010010: data <= 32'hbf463daa;
    11'b01000010011: data <= 32'hbc8b3752;
    11'b01000010100: data <= 32'h39fbbade;
    11'b01000010101: data <= 32'h4014b8db;
    11'b01000010110: data <= 32'h3d6d3b13;
    11'b01000010111: data <= 32'had163f03;
    11'b01000011000: data <= 32'hb07e3d78;
    11'b01000011001: data <= 32'h3c1239aa;
    11'b01000011010: data <= 32'h3d063483;
    11'b01000011011: data <= 32'haf4db857;
    11'b01000011100: data <= 32'hbc95bf1f;
    11'b01000011101: data <= 32'hb252c03d;
    11'b01000011110: data <= 32'h3e31bb77;
    11'b01000011111: data <= 32'h3f4c353c;
    11'b01000100000: data <= 32'h37072e37;
    11'b01000100001: data <= 32'hbb0fbae4;
    11'b01000100010: data <= 32'hbcf8b8ed;
    11'b01000100011: data <= 32'hbd7e3a34;
    11'b01000100100: data <= 32'hbecc3cac;
    11'b01000100101: data <= 32'hbdabb541;
    11'b01000100110: data <= 32'hb241bef9;
    11'b01000100111: data <= 32'h39ecbbfd;
    11'b01000101000: data <= 32'h36023c89;
    11'b01000101001: data <= 32'hb5404088;
    11'b01000101010: data <= 32'h2e263edf;
    11'b01000101011: data <= 32'h3c653b2e;
    11'b01000101100: data <= 32'h3aab399d;
    11'b01000101101: data <= 32'hb9d6365b;
    11'b01000101110: data <= 32'hbd52b856;
    11'b01000101111: data <= 32'h34fcbccc;
    11'b01000110000: data <= 32'h40d1ba4d;
    11'b01000110001: data <= 32'h4103b0c4;
    11'b01000110010: data <= 32'h3a6cb61d;
    11'b01000110011: data <= 32'hb7ebbb02;
    11'b01000110100: data <= 32'hb7aeb51c;
    11'b01000110101: data <= 32'hb5c73a5a;
    11'b01000110110: data <= 32'hbc003841;
    11'b01000110111: data <= 32'hbe02bd7e;
    11'b01000111000: data <= 32'hbbbbc138;
    11'b01000111001: data <= 32'hafabbd93;
    11'b01000111010: data <= 32'ha81f3b90;
    11'b01000111011: data <= 32'hb4d13f6b;
    11'b01000111100: data <= 32'h28dd3c43;
    11'b01000111101: data <= 32'h380b37e9;
    11'b01000111110: data <= 32'hb1b93c2c;
    11'b01000111111: data <= 32'hbe613dc4;
    11'b01001000000: data <= 32'hbe8938ed;
    11'b01001000001: data <= 32'h36b8b840;
    11'b01001000010: data <= 32'h40e7b97d;
    11'b01001000011: data <= 32'h4095b0d5;
    11'b01001000100: data <= 32'h39921fc7;
    11'b01001000101: data <= 32'h2684adc8;
    11'b01001000110: data <= 32'h39be35eb;
    11'b01001000111: data <= 32'h3ba43b4d;
    11'b01001001000: data <= 32'hb3742f52;
    11'b01001001001: data <= 32'hbdcabf6e;
    11'b01001001010: data <= 32'hbcc0c1a4;
    11'b01001001011: data <= 32'hac0ebe1b;
    11'b01001001100: data <= 32'h36943634;
    11'b01001001101: data <= 32'h2f433998;
    11'b01001001110: data <= 32'hac13b315;
    11'b01001001111: data <= 32'hb132b2f5;
    11'b01001010000: data <= 32'hbbe43cb2;
    11'b01001010001: data <= 32'hc0394003;
    11'b01001010010: data <= 32'hbf943bd2;
    11'b01001010011: data <= 32'ha64ab8d1;
    11'b01001010100: data <= 32'h3e2dbaba;
    11'b01001010101: data <= 32'h3cef2f77;
    11'b01001010110: data <= 32'h31653a80;
    11'b01001010111: data <= 32'h36593af0;
    11'b01001011000: data <= 32'h3e9c3c05;
    11'b01001011001: data <= 32'h3ef93c99;
    11'b01001011010: data <= 32'h276d351b;
    11'b01001011011: data <= 32'hbdc8bd5c;
    11'b01001011100: data <= 32'hbb33c048;
    11'b01001011101: data <= 32'h39babd13;
    11'b01001011110: data <= 32'h3d5eb28b;
    11'b01001011111: data <= 32'h397db821;
    11'b01001100000: data <= 32'h91d5bd5d;
    11'b01001100001: data <= 32'hb4a0b9b9;
    11'b01001100010: data <= 32'hbb473c9d;
    11'b01001100011: data <= 32'hbf653f8b;
    11'b01001100100: data <= 32'hbfa836a5;
    11'b01001100101: data <= 32'hba17bd67;
    11'b01001100110: data <= 32'h32c2bcf1;
    11'b01001100111: data <= 32'ha80934f8;
    11'b01001101000: data <= 32'hb6a63d38;
    11'b01001101001: data <= 32'h37ca3ccf;
    11'b01001101010: data <= 32'h3f673c5a;
    11'b01001101011: data <= 32'h3e433d6c;
    11'b01001101100: data <= 32'hb6b63c4c;
    11'b01001101101: data <= 32'hbe83acc0;
    11'b01001101110: data <= 32'hb79fbb8d;
    11'b01001101111: data <= 32'h3e10ba30;
    11'b01001110000: data <= 32'h3fffb811;
    11'b01001110001: data <= 32'h3bd6bc6a;
    11'b01001110010: data <= 32'h3341be7d;
    11'b01001110011: data <= 32'h351db8f6;
    11'b01001110100: data <= 32'h2ff23c9d;
    11'b01001110101: data <= 32'hbb1f3d6b;
    11'b01001110110: data <= 32'hbe98b845;
    11'b01001110111: data <= 32'hbd5dc05d;
    11'b01001111000: data <= 32'hb9fbbe5e;
    11'b01001111001: data <= 32'hb9ce334a;
    11'b01001111010: data <= 32'hb9073c0a;
    11'b01001111011: data <= 32'h36343843;
    11'b01001111100: data <= 32'h3d81373e;
    11'b01001111101: data <= 32'h39723d72;
    11'b01001111110: data <= 32'hbcf13fad;
    11'b01001111111: data <= 32'hbfab3cb1;
    11'b01010000000: data <= 32'hb4fb2727;
    11'b01010000001: data <= 32'h3e8fb648;
    11'b01010000010: data <= 32'h3f15b70c;
    11'b01010000011: data <= 32'h3964bab7;
    11'b01010000100: data <= 32'h370cbbfa;
    11'b01010000101: data <= 32'h3d489860;
    11'b01010000110: data <= 32'h3e163d1a;
    11'b01010000111: data <= 32'h32143b65;
    11'b01010001000: data <= 32'hbd20bc45;
    11'b01010001001: data <= 32'hbdd8c0c4;
    11'b01010001010: data <= 32'hba8fbe40;
    11'b01010001011: data <= 32'hb7a7abcd;
    11'b01010001100: data <= 32'hb50e2913;
    11'b01010001101: data <= 32'h34b9baa1;
    11'b01010001110: data <= 32'h39dcb896;
    11'b01010001111: data <= 32'hb0a03c9f;
    11'b01010010000: data <= 32'hbeff40b6;
    11'b01010010001: data <= 32'hc01d3ea7;
    11'b01010010010: data <= 32'hb83f3201;
    11'b01010010011: data <= 32'h3b32b67e;
    11'b01010010100: data <= 32'h392cb19e;
    11'b01010010101: data <= 32'hb11cadc5;
    11'b01010010110: data <= 32'h376eab16;
    11'b01010010111: data <= 32'h40373912;
    11'b01010011000: data <= 32'h40e03dbb;
    11'b01010011001: data <= 32'h39b93b9b;
    11'b01010011010: data <= 32'hbc60b995;
    11'b01010011011: data <= 32'hbca3be99;
    11'b01010011100: data <= 32'hafa4bc11;
    11'b01010011101: data <= 32'h3669b4ec;
    11'b01010011110: data <= 32'h3405bc11;
    11'b01010011111: data <= 32'h3507c028;
    11'b01010100000: data <= 32'h379abd74;
    11'b01010100001: data <= 32'hb2413b41;
    11'b01010100010: data <= 32'hbdcc4065;
    11'b01010100011: data <= 32'hbf463cca;
    11'b01010100100: data <= 32'hbb7bb78d;
    11'b01010100101: data <= 32'hb451ba39;
    11'b01010100110: data <= 32'hb9fd28b7;
    11'b01010100111: data <= 32'hbc3e37cc;
    11'b01010101000: data <= 32'h3499362b;
    11'b01010101001: data <= 32'h407e3996;
    11'b01010101010: data <= 32'h40be3dad;
    11'b01010101011: data <= 32'h36553d97;
    11'b01010101100: data <= 32'hbce83678;
    11'b01010101101: data <= 32'hb9d7b53c;
    11'b01010101110: data <= 32'h39cfb20d;
    11'b01010101111: data <= 32'h3c8eb4fd;
    11'b01010110000: data <= 32'h3858be1a;
    11'b01010110001: data <= 32'h35dec0f8;
    11'b01010110010: data <= 32'h3a7abdc2;
    11'b01010110011: data <= 32'h396c3a97;
    11'b01010110100: data <= 32'hb6013ea8;
    11'b01010110101: data <= 32'hbcdc3383;
    11'b01010110110: data <= 32'hbcc4bd6e;
    11'b01010110111: data <= 32'hbc87bc93;
    11'b01010111000: data <= 32'hbe582d80;
    11'b01010111001: data <= 32'hbdf636da;
    11'b01010111010: data <= 32'h2c2fb02d;
    11'b01010111011: data <= 32'h3f0fa87d;
    11'b01010111100: data <= 32'h3e023c65;
    11'b01010111101: data <= 32'hb7203fa1;
    11'b01010111110: data <= 32'hbe1e3e2a;
    11'b01010111111: data <= 32'hb7873a69;
    11'b01011000000: data <= 32'h3c30373f;
    11'b01011000001: data <= 32'h3c38aceb;
    11'b01011000010: data <= 32'h312bbcfb;
    11'b01011000011: data <= 32'h3472bf9f;
    11'b01011000100: data <= 32'h3deabaa6;
    11'b01011000101: data <= 32'h3fd23ba1;
    11'b01011000110: data <= 32'h3af43cac;
    11'b01011000111: data <= 32'hb863b759;
    11'b01011001000: data <= 32'hbc66bec8;
    11'b01011001001: data <= 32'hbcb4bc41;
    11'b01011001010: data <= 32'hbda72c4c;
    11'b01011001011: data <= 32'hbcebb328;
    11'b01011001100: data <= 32'ha862bd76;
    11'b01011001101: data <= 32'h3c50bce8;
    11'b01011001110: data <= 32'h38683887;
    11'b01011001111: data <= 32'hbc584030;
    11'b01011010000: data <= 32'hbe933ff5;
    11'b01011010001: data <= 32'hb7503c44;
    11'b01011010010: data <= 32'h38d73857;
    11'b01011010011: data <= 32'h2bcf331d;
    11'b01011010100: data <= 32'hbaa7b77f;
    11'b01011010101: data <= 32'ha8ecbaf8;
    11'b01011010110: data <= 32'h3ff1ad3f;
    11'b01011010111: data <= 32'h41a23c6e;
    11'b01011011000: data <= 32'h3e1c3c01;
    11'b01011011001: data <= 32'hb290b5d8;
    11'b01011011010: data <= 32'hb9d0bc61;
    11'b01011011011: data <= 32'hb74ab5f2;
    11'b01011011100: data <= 32'hb7a4312f;
    11'b01011011101: data <= 32'hb891bbe0;
    11'b01011011110: data <= 32'h9838c11b;
    11'b01011011111: data <= 32'h3953c059;
    11'b01011100000: data <= 32'h33f12f02;
    11'b01011100001: data <= 32'hbb6a3f4b;
    11'b01011100010: data <= 32'hbd1f3e04;
    11'b01011100011: data <= 32'hb83d362e;
    11'b01011100100: data <= 32'hb4282f17;
    11'b01011100101: data <= 32'hbd1036ab;
    11'b01011100110: data <= 32'hbfa4335c;
    11'b01011100111: data <= 32'hb781b28f;
    11'b01011101000: data <= 32'h3fe33030;
    11'b01011101001: data <= 32'h41753bff;
    11'b01011101010: data <= 32'h3ce63c8d;
    11'b01011101011: data <= 32'hb5b436e4;
    11'b01011101100: data <= 32'hb4ec30e2;
    11'b01011101101: data <= 32'h37be3931;
    11'b01011101110: data <= 32'h374f3732;
    11'b01011101111: data <= 32'hb016bd37;
    11'b01011110000: data <= 32'ha1fec1e0;
    11'b01011110001: data <= 32'h39c0c09d;
    11'b01011110010: data <= 32'h3a8d9a7a;
    11'b01011110011: data <= 32'h2bcd3d1f;
    11'b01011110100: data <= 32'hb7b33779;
    11'b01011110101: data <= 32'hb773b954;
    11'b01011110110: data <= 32'hbb3bb672;
    11'b01011110111: data <= 32'hc02a37fa;
    11'b01011111000: data <= 32'hc0e036b0;
    11'b01011111001: data <= 32'hba31b6d6;
    11'b01011111010: data <= 32'h3dd2b803;
    11'b01011111011: data <= 32'h3f3337e2;
    11'b01011111100: data <= 32'h33f43d3f;
    11'b01011111101: data <= 32'hba5b3d4c;
    11'b01011111110: data <= 32'ha8a33d0d;
    11'b01011111111: data <= 32'h3c123db7;
    11'b01100000000: data <= 32'h393d3a96;
    11'b01100000001: data <= 32'hb644bbab;
    11'b01100000010: data <= 32'hb441c09f;
    11'b01100000011: data <= 32'h3c34be65;
    11'b01100000100: data <= 32'h3f5733b6;
    11'b01100000101: data <= 32'h3d233a47;
    11'b01100000110: data <= 32'h35bbb698;
    11'b01100000111: data <= 32'hb1cfbd16;
    11'b01100001000: data <= 32'hbacdb74b;
    11'b01100001001: data <= 32'hbf8338f1;
    11'b01100001010: data <= 32'hc03d2de2;
    11'b01100001011: data <= 32'hba53bd90;
    11'b01100001100: data <= 32'h3a2ebea8;
    11'b01100001101: data <= 32'h3981b392;
    11'b01100001110: data <= 32'hb92b3d07;
    11'b01100001111: data <= 32'hbc393e92;
    11'b01100010000: data <= 32'h2d763e08;
    11'b01100010001: data <= 32'h3b143e0b;
    11'b01100010010: data <= 32'habdb3c54;
    11'b01100010011: data <= 32'hbd61b1c0;
    11'b01100010100: data <= 32'hba52bc8f;
    11'b01100010101: data <= 32'h3d20b8e8;
    11'b01100010110: data <= 32'h4113386d;
    11'b01100010111: data <= 32'h3fbe384e;
    11'b01100011000: data <= 32'h39f9b8db;
    11'b01100011001: data <= 32'h328ebba1;
    11'b01100011010: data <= 32'haf3731cb;
    11'b01100011011: data <= 32'hbaa13b5d;
    11'b01100011100: data <= 32'hbd01b5e7;
    11'b01100011101: data <= 32'hb8c9c0ca;
    11'b01100011110: data <= 32'h34e8c13b;
    11'b01100011111: data <= 32'h2f86ba4c;
    11'b01100100000: data <= 32'hba313b56;
    11'b01100100001: data <= 32'hba263c7a;
    11'b01100100010: data <= 32'h32bb39e7;
    11'b01100100011: data <= 32'h35533b3e;
    11'b01100100100: data <= 32'hbcc03c82;
    11'b01100100101: data <= 32'hc0de3869;
    11'b01100100110: data <= 32'hbd6fb34b;
    11'b01100100111: data <= 32'h3c94aef3;
    11'b01100101000: data <= 32'h40c6385e;
    11'b01100101001: data <= 32'h3e4237f0;
    11'b01100101010: data <= 32'h3774b022;
    11'b01100101011: data <= 32'h37f92ce7;
    11'b01100101100: data <= 32'h3ac93cdc;
    11'b01100101101: data <= 32'h35453d86;
    11'b01100101110: data <= 32'hb823b824;
    11'b01100101111: data <= 32'hb7afc165;
    11'b01100110000: data <= 32'h32a2c168;
    11'b01100110001: data <= 32'h35efba90;
    11'b01100110010: data <= 32'ha577376a;
    11'b01100110011: data <= 32'h28e42be6;
    11'b01100110100: data <= 32'h3793b81f;
    11'b01100110101: data <= 32'hae662efe;
    11'b01100110110: data <= 32'hbf9d3c3e;
    11'b01100110111: data <= 32'hc1e23ae8;
    11'b01100111000: data <= 32'hbe8db073;
    11'b01100111001: data <= 32'h3964b7cb;
    11'b01100111010: data <= 32'h3dbb2a25;
    11'b01100111011: data <= 32'h36913754;
    11'b01100111100: data <= 32'hb3993829;
    11'b01100111101: data <= 32'h38e43c44;
    11'b01100111110: data <= 32'h3dec4000;
    11'b01100111111: data <= 32'h3aa13f23;
    11'b01101000000: data <= 32'hb812b17e;
    11'b01101000001: data <= 32'hb99cc012;
    11'b01101000010: data <= 32'h3540bf5e;
    11'b01101000011: data <= 32'h3c77b566;
    11'b01101000100: data <= 32'h3c413000;
    11'b01101000101: data <= 32'h3b3cbb2d;
    11'b01101000110: data <= 32'h3abcbda5;
    11'b01101000111: data <= 32'h1a84b369;
    11'b01101001000: data <= 32'hbe9f3c78;
    11'b01101001001: data <= 32'hc10139e5;
    11'b01101001010: data <= 32'hbdcfba85;
    11'b01101001011: data <= 32'h305ebdf7;
    11'b01101001100: data <= 32'h340eb9c0;
    11'b01101001101: data <= 32'hba1c345a;
    11'b01101001110: data <= 32'hba6339ed;
    11'b01101001111: data <= 32'h39253d0c;
    11'b01101010000: data <= 32'h3e1f3ffd;
    11'b01101010001: data <= 32'h368e3f8f;
    11'b01101010010: data <= 32'hbd2037c0;
    11'b01101010011: data <= 32'hbd0dba71;
    11'b01101010100: data <= 32'h364ab8ba;
    11'b01101010101: data <= 32'h3eb8347f;
    11'b01101010110: data <= 32'h3e9e9f26;
    11'b01101010111: data <= 32'h3cfbbd06;
    11'b01101011000: data <= 32'h3c84bd98;
    11'b01101011001: data <= 32'h3932326c;
    11'b01101011010: data <= 32'hb86c3dca;
    11'b01101011011: data <= 32'hbd8d3768;
    11'b01101011100: data <= 32'hbba5be93;
    11'b01101011101: data <= 32'hb241c0be;
    11'b01101011110: data <= 32'hb771bd07;
    11'b01101011111: data <= 32'hbcd1a740;
    11'b01101100000: data <= 32'hb9f1344f;
    11'b01101100001: data <= 32'h3a363716;
    11'b01101100010: data <= 32'h3cb43cb1;
    11'b01101100011: data <= 32'hb8183e94;
    11'b01101100100: data <= 32'hc0933c48;
    11'b01101100101: data <= 32'hbf6333a8;
    11'b01101100110: data <= 32'h33ac3376;
    11'b01101100111: data <= 32'h3e283846;
    11'b01101101000: data <= 32'h3cf3a836;
    11'b01101101001: data <= 32'h3a40bbd7;
    11'b01101101010: data <= 32'h3ca8b8c9;
    11'b01101101011: data <= 32'h3dde3c8b;
    11'b01101101100: data <= 32'h39c93fc8;
    11'b01101101101: data <= 32'hb5523613;
    11'b01101101110: data <= 32'hb866bfaa;
    11'b01101101111: data <= 32'hb3fcc0d4;
    11'b01101110000: data <= 32'hb692bc96;
    11'b01101110001: data <= 32'hb9a6b440;
    11'b01101110010: data <= 32'haaf7b943;
    11'b01101110011: data <= 32'h3c5abb55;
    11'b01101110100: data <= 32'h3acc2bf0;
    11'b01101110101: data <= 32'hbca63d16;
    11'b01101110110: data <= 32'hc1823d3c;
    11'b01101110111: data <= 32'hc00d3829;
    11'b01101111000: data <= 32'hac263045;
    11'b01101111001: data <= 32'h398a31df;
    11'b01101111010: data <= 32'ha307afb8;
    11'b01101111011: data <= 32'hb328b787;
    11'b01101111100: data <= 32'h3bb334b6;
    11'b01101111101: data <= 32'h40013f8a;
    11'b01101111110: data <= 32'h3d9f4095;
    11'b01101111111: data <= 32'ha5f138e5;
    11'b01110000000: data <= 32'hb8b5bd59;
    11'b01110000001: data <= 32'hb159bddd;
    11'b01110000010: data <= 32'h317ab625;
    11'b01110000011: data <= 32'h33f9b4b6;
    11'b01110000100: data <= 32'h3a2fbe05;
    11'b01110000101: data <= 32'h3dc3bff3;
    11'b01110000110: data <= 32'h3b24b8ca;
    11'b01110000111: data <= 32'hbbc33c70;
    11'b01110001000: data <= 32'hc07b3ccc;
    11'b01110001001: data <= 32'hbe5d2607;
    11'b01110001010: data <= 32'hb4f6b9aa;
    11'b01110001011: data <= 32'hb5f0b848;
    11'b01110001100: data <= 32'hbd6cb530;
    11'b01110001101: data <= 32'hbc7ab3b5;
    11'b01110001110: data <= 32'h39ee3825;
    11'b01110001111: data <= 32'h40163f4b;
    11'b01110010000: data <= 32'h3cb24060;
    11'b01110010001: data <= 32'hb8ce3c04;
    11'b01110010010: data <= 32'hbc54b307;
    11'b01110010011: data <= 32'hb081aac2;
    11'b01110010100: data <= 32'h3992389f;
    11'b01110010101: data <= 32'h3ab9b0ae;
    11'b01110010110: data <= 32'h3c4bbf56;
    11'b01110010111: data <= 32'h3e45c056;
    11'b01110011000: data <= 32'h3d41b650;
    11'b01110011001: data <= 32'h26cf3d61;
    11'b01110011010: data <= 32'hbbca3bc7;
    11'b01110011011: data <= 32'hba00b9d5;
    11'b01110011100: data <= 32'hb579be3d;
    11'b01110011101: data <= 32'hbc29bc30;
    11'b01110011110: data <= 32'hbffdb81b;
    11'b01110011111: data <= 32'hbd4cb845;
    11'b01110100000: data <= 32'h39fcb29e;
    11'b01110100001: data <= 32'h3ef03aea;
    11'b01110100010: data <= 32'h35bb3e72;
    11'b01110100011: data <= 32'hbe323d20;
    11'b01110100100: data <= 32'hbe973a15;
    11'b01110100101: data <= 32'hb3533bd4;
    11'b01110100110: data <= 32'h397c3c82;
    11'b01110100111: data <= 32'h3805a048;
    11'b01110101000: data <= 32'h37efbe60;
    11'b01110101001: data <= 32'h3d31bdfe;
    11'b01110101010: data <= 32'h3f4e3742;
    11'b01110101011: data <= 32'h3ce83f4b;
    11'b01110101100: data <= 32'h34ad3ae4;
    11'b01110101101: data <= 32'ha46abc56;
    11'b01110101110: data <= 32'hb231bea9;
    11'b01110101111: data <= 32'hbc09bac7;
    11'b01110110000: data <= 32'hbe9cb7bc;
    11'b01110110001: data <= 32'hba10bcb2;
    11'b01110110010: data <= 32'h3c21bdf1;
    11'b01110110011: data <= 32'h3da3b74b;
    11'b01110110100: data <= 32'hb5573b19;
    11'b01110110101: data <= 32'hc0203d1f;
    11'b01110110110: data <= 32'hbf0c3c32;
    11'b01110110111: data <= 32'hb4f73c38;
    11'b01110111000: data <= 32'h2e343b81;
    11'b01110111001: data <= 32'hb958aa67;
    11'b01110111010: data <= 32'hb9acbc6c;
    11'b01110111011: data <= 32'h39e1b8cf;
    11'b01110111100: data <= 32'h40303cee;
    11'b01110111101: data <= 32'h3f9b4042;
    11'b01110111110: data <= 32'h3a663b56;
    11'b01110111111: data <= 32'h30d7b9d7;
    11'b01111000000: data <= 32'ha88eba5c;
    11'b01111000001: data <= 32'hb75d2e82;
    11'b01111000010: data <= 32'hb9d5b0f2;
    11'b01111000011: data <= 32'h2d30bef4;
    11'b01111000100: data <= 32'h3d76c112;
    11'b01111000101: data <= 32'h3d49bd54;
    11'b01111000110: data <= 32'hb54e3790;
    11'b01111000111: data <= 32'hbe803c3b;
    11'b01111001000: data <= 32'hbca538b4;
    11'b01111001001: data <= 32'hb2d2347d;
    11'b01111001010: data <= 32'hb9703380;
    11'b01111001011: data <= 32'hbfeeb3e0;
    11'b01111001100: data <= 32'hbf57ba4f;
    11'b01111001101: data <= 32'h330db324;
    11'b01111001110: data <= 32'h3fef3cfe;
    11'b01111001111: data <= 32'h3ed03f8c;
    11'b01111010000: data <= 32'h352a3bf1;
    11'b01111010001: data <= 32'hb4ab2ebd;
    11'b01111010010: data <= 32'h987f38af;
    11'b01111010011: data <= 32'h2f683d37;
    11'b01111010100: data <= 32'ha4f6351f;
    11'b01111010101: data <= 32'h3751bf85;
    11'b01111010110: data <= 32'h3d8cc17d;
    11'b01111010111: data <= 32'h3dd8bd0c;
    11'b01111011000: data <= 32'h365538ea;
    11'b01111011001: data <= 32'hb6573a7e;
    11'b01111011010: data <= 32'hacf5b202;
    11'b01111011011: data <= 32'h2ebdb938;
    11'b01111011100: data <= 32'hbc88b591;
    11'b01111011101: data <= 32'hc14bb5d6;
    11'b01111011110: data <= 32'hc06ababe;
    11'b01111011111: data <= 32'h2d8bb992;
    11'b01111100000: data <= 32'h3e87355d;
    11'b01111100001: data <= 32'h3b0d3c4d;
    11'b01111100010: data <= 32'hb9613b42;
    11'b01111100011: data <= 32'hbb543ac8;
    11'b01111100100: data <= 32'haa2f3e8e;
    11'b01111100101: data <= 32'h34c9401b;
    11'b01111100110: data <= 32'hb017392e;
    11'b01111100111: data <= 32'hac0ebe47;
    11'b01111101000: data <= 32'h3b37c029;
    11'b01111101001: data <= 32'h3e73b66f;
    11'b01111101010: data <= 32'h3d603c88;
    11'b01111101011: data <= 32'h3b1f396c;
    11'b01111101100: data <= 32'h3b17b992;
    11'b01111101101: data <= 32'h37e2bbb4;
    11'b01111101110: data <= 32'hbc01b2ed;
    11'b01111101111: data <= 32'hc0a4b0c8;
    11'b01111110000: data <= 32'hbeabbc8d;
    11'b01111110001: data <= 32'h3624bede;
    11'b01111110010: data <= 32'h3d2cbc00;
    11'b01111110011: data <= 32'h2c8e2e3f;
    11'b01111110100: data <= 32'hbd7538f9;
    11'b01111110101: data <= 32'hbc6d3c05;
    11'b01111110110: data <= 32'h25883efa;
    11'b01111110111: data <= 32'h27533fbc;
    11'b01111111000: data <= 32'hbc2a390a;
    11'b01111111001: data <= 32'hbd1abc45;
    11'b01111111010: data <= 32'h2cb5bc60;
    11'b01111111011: data <= 32'h3e3e3840;
    11'b01111111100: data <= 32'h3f6e3e17;
    11'b01111111101: data <= 32'h3dbe38ed;
    11'b01111111110: data <= 32'h3cafb907;
    11'b01111111111: data <= 32'h39c4b57b;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    