
module memory_rom_40(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbc543c9d;
    11'b00000000001: data <= 32'hb89a3996;
    11'b00000000010: data <= 32'h393cb933;
    11'b00000000011: data <= 32'h3f08b929;
    11'b00000000100: data <= 32'h3d773c36;
    11'b00000000101: data <= 32'hac0d40b3;
    11'b00000000110: data <= 32'hb86a3f14;
    11'b00000000111: data <= 32'h37853477;
    11'b00000001000: data <= 32'h3ce2b8a8;
    11'b00000001001: data <= 32'h35e6baef;
    11'b00000001010: data <= 32'hb9fcbd60;
    11'b00000001011: data <= 32'hb007be98;
    11'b00000001100: data <= 32'h3eb2bb5e;
    11'b00000001101: data <= 32'h404c345d;
    11'b00000001110: data <= 32'h371a36c6;
    11'b00000001111: data <= 32'hbe21b810;
    11'b00000010000: data <= 32'hbfc6bad1;
    11'b00000010001: data <= 32'hbd312d79;
    11'b00000010010: data <= 32'hbbdb39df;
    11'b00000010011: data <= 32'hbba2b43f;
    11'b00000010100: data <= 32'hb579be6e;
    11'b00000010101: data <= 32'h386bbc03;
    11'b00000010110: data <= 32'h38a13d63;
    11'b00000010111: data <= 32'hb1a141af;
    11'b00000011000: data <= 32'hb5b7401f;
    11'b00000011001: data <= 32'h35bf376c;
    11'b00000011010: data <= 32'h38c6ad2c;
    11'b00000011011: data <= 32'hb55d30d9;
    11'b00000011100: data <= 32'hbb34b0bd;
    11'b00000011101: data <= 32'h3730bb1f;
    11'b00000011110: data <= 32'h4119bb4a;
    11'b00000011111: data <= 32'h4197b15e;
    11'b00000100000: data <= 32'h3a6230b6;
    11'b00000100001: data <= 32'hbc51b4cd;
    11'b00000100010: data <= 32'hbc5fb758;
    11'b00000100011: data <= 32'hb4912b1a;
    11'b00000100100: data <= 32'hb6700fd3;
    11'b00000100101: data <= 32'hbcadbd70;
    11'b00000100110: data <= 32'hbc67c0ed;
    11'b00000100111: data <= 32'haf89bd94;
    11'b00000101000: data <= 32'h36803c69;
    11'b00000101001: data <= 32'ha95b40b0;
    11'b00000101010: data <= 32'hb7bd3d89;
    11'b00000101011: data <= 32'hb601309d;
    11'b00000101100: data <= 32'hb8083616;
    11'b00000101101: data <= 32'hbcd53cd8;
    11'b00000101110: data <= 32'hbccb3ad7;
    11'b00000101111: data <= 32'h3818b72a;
    11'b00000110000: data <= 32'h4107bb6c;
    11'b00000110001: data <= 32'h411aadfd;
    11'b00000110010: data <= 32'h3a0f39c4;
    11'b00000110011: data <= 32'hb72a38f9;
    11'b00000110100: data <= 32'h30803410;
    11'b00000110101: data <= 32'h3b5930db;
    11'b00000110110: data <= 32'h3159b653;
    11'b00000110111: data <= 32'hbcf0bf1b;
    11'b00000111000: data <= 32'hbd02c149;
    11'b00000111001: data <= 32'h30a7be5c;
    11'b00000111010: data <= 32'h3c1e36e5;
    11'b00000111011: data <= 32'h36b13c8b;
    11'b00000111100: data <= 32'hb90d31a0;
    11'b00000111101: data <= 32'hbc43b670;
    11'b00000111110: data <= 32'hbd1538f8;
    11'b00000111111: data <= 32'hbec43edd;
    11'b00001000000: data <= 32'hbe113c0b;
    11'b00001000001: data <= 32'hab43b9c7;
    11'b00001000010: data <= 32'h3e1dbc98;
    11'b00001000011: data <= 32'h3e2f339f;
    11'b00001000100: data <= 32'h36003e69;
    11'b00001000101: data <= 32'h26fe3e56;
    11'b00001000110: data <= 32'h3c193ae7;
    11'b00001000111: data <= 32'h3e0f36de;
    11'b00001001000: data <= 32'h333fac5f;
    11'b00001001001: data <= 32'hbd3bbca1;
    11'b00001001010: data <= 32'hbb1ebff4;
    11'b00001001011: data <= 32'h3c31bde0;
    11'b00001001100: data <= 32'h400ab464;
    11'b00001001101: data <= 32'h3bdfa9e9;
    11'b00001001110: data <= 32'hb867ba25;
    11'b00001001111: data <= 32'hbc61b9ac;
    11'b00001010000: data <= 32'hbc57395b;
    11'b00001010001: data <= 32'hbdb73e09;
    11'b00001010010: data <= 32'hbea834ba;
    11'b00001010011: data <= 32'hbb6ebe4c;
    11'b00001010100: data <= 32'h3256be3e;
    11'b00001010101: data <= 32'h370236e8;
    11'b00001010110: data <= 32'ha6674013;
    11'b00001010111: data <= 32'h31b63f51;
    11'b00001011000: data <= 32'h3c7d3b70;
    11'b00001011001: data <= 32'h3ca439fa;
    11'b00001011010: data <= 32'hb5983abb;
    11'b00001011011: data <= 32'hbe1630ca;
    11'b00001011100: data <= 32'hb739bb59;
    11'b00001011101: data <= 32'h3f53bc9f;
    11'b00001011110: data <= 32'h413fb92a;
    11'b00001011111: data <= 32'h3d0fb831;
    11'b00001100000: data <= 32'hb346bad2;
    11'b00001100001: data <= 32'hb546b78e;
    11'b00001100010: data <= 32'h270f3993;
    11'b00001100011: data <= 32'hb8733b84;
    11'b00001100100: data <= 32'hbe4bb968;
    11'b00001100101: data <= 32'hbe64c0c8;
    11'b00001100110: data <= 32'hb952bfb0;
    11'b00001100111: data <= 32'haa4d3435;
    11'b00001101000: data <= 32'had423e63;
    11'b00001101001: data <= 32'h2e1f3c43;
    11'b00001101010: data <= 32'h38933588;
    11'b00001101011: data <= 32'h32c63b51;
    11'b00001101100: data <= 32'hbcb93f33;
    11'b00001101101: data <= 32'hbf4e3d59;
    11'b00001101110: data <= 32'hb5d8b09d;
    11'b00001101111: data <= 32'h3f4cbb8e;
    11'b00001110000: data <= 32'h409cb8bf;
    11'b00001110001: data <= 32'h3bf9b0c0;
    11'b00001110010: data <= 32'h3056af50;
    11'b00001110011: data <= 32'h3a6c3203;
    11'b00001110100: data <= 32'h3da03aa3;
    11'b00001110101: data <= 32'h35b3388c;
    11'b00001110110: data <= 32'hbd84bc63;
    11'b00001110111: data <= 32'hbefbc106;
    11'b00001111000: data <= 32'hb8ddbfbb;
    11'b00001111001: data <= 32'h35b6b198;
    11'b00001111010: data <= 32'h34dd37ba;
    11'b00001111011: data <= 32'h19b4b4f5;
    11'b00001111100: data <= 32'haa84b85e;
    11'b00001111101: data <= 32'hb8433afb;
    11'b00001111110: data <= 32'hbe80408e;
    11'b00001111111: data <= 32'hc0043ed1;
    11'b00010000000: data <= 32'hb9eeb161;
    11'b00010000001: data <= 32'h3b65bc3f;
    11'b00010000010: data <= 32'h3c94b525;
    11'b00010000011: data <= 32'h346a390a;
    11'b00010000100: data <= 32'h350c3a63;
    11'b00010000101: data <= 32'h3e933a2f;
    11'b00010000110: data <= 32'h40703c16;
    11'b00010000111: data <= 32'h399639ff;
    11'b00010001000: data <= 32'hbd40b86a;
    11'b00010001001: data <= 32'hbdbfbee3;
    11'b00010001010: data <= 32'h312ebdf7;
    11'b00010001011: data <= 32'h3d11b8ab;
    11'b00010001100: data <= 32'h3ad1b927;
    11'b00010001101: data <= 32'h29b5bde5;
    11'b00010001110: data <= 32'hb1a7bcaa;
    11'b00010001111: data <= 32'hb68439f5;
    11'b00010010000: data <= 32'hbd00403a;
    11'b00010010001: data <= 32'hbf783c93;
    11'b00010010010: data <= 32'hbd4ebb43;
    11'b00010010011: data <= 32'hb582bdcf;
    11'b00010010100: data <= 32'hb1f3aff7;
    11'b00010010101: data <= 32'hb76d3c75;
    11'b00010010110: data <= 32'h34123c5a;
    11'b00010010111: data <= 32'h3f133a0c;
    11'b00010011000: data <= 32'h40153c60;
    11'b00010011001: data <= 32'h34503d94;
    11'b00010011010: data <= 32'hbdf73985;
    11'b00010011011: data <= 32'hbc14b6ee;
    11'b00010011100: data <= 32'h3ba3ba8f;
    11'b00010011101: data <= 32'h3f98b9b1;
    11'b00010011110: data <= 32'h3c4dbc8c;
    11'b00010011111: data <= 32'h316ebf07;
    11'b00010100000: data <= 32'h35b0bc77;
    11'b00010100001: data <= 32'h391c39b7;
    11'b00010100010: data <= 32'hb17d3e52;
    11'b00010100011: data <= 32'hbda73254;
    11'b00010100100: data <= 32'hbeeabeef;
    11'b00010100101: data <= 32'hbcd7bf1d;
    11'b00010100110: data <= 32'hbb24b09b;
    11'b00010100111: data <= 32'hba073af7;
    11'b00010101000: data <= 32'h2d683637;
    11'b00010101001: data <= 32'h3d0ea3a4;
    11'b00010101010: data <= 32'h3c9b3b42;
    11'b00010101011: data <= 32'hb8674026;
    11'b00010101100: data <= 32'hbf1d3f7a;
    11'b00010101101: data <= 32'hbaa238a1;
    11'b00010101110: data <= 32'h3c6eb550;
    11'b00010101111: data <= 32'h3e91b848;
    11'b00010110000: data <= 32'h392bba78;
    11'b00010110001: data <= 32'h3275bc72;
    11'b00010110010: data <= 32'h3cd8b7ee;
    11'b00010110011: data <= 32'h40013ab6;
    11'b00010110100: data <= 32'h3beb3c94;
    11'b00010110101: data <= 32'hbb3bb590;
    11'b00010110110: data <= 32'hbedbbfab;
    11'b00010110111: data <= 32'hbcc9bea1;
    11'b00010111000: data <= 32'hb8ecb489;
    11'b00010111001: data <= 32'hb71925ad;
    11'b00010111010: data <= 32'ha4edbbb9;
    11'b00010111011: data <= 32'h38e0bca4;
    11'b00010111100: data <= 32'h3511382e;
    11'b00010111101: data <= 32'hbc3940b7;
    11'b00010111110: data <= 32'hbf74408c;
    11'b00010111111: data <= 32'hbb9139be;
    11'b00011000000: data <= 32'h374eb53d;
    11'b00011000001: data <= 32'h3812b397;
    11'b00011000010: data <= 32'hb533a67d;
    11'b00011000011: data <= 32'h25d3b0a4;
    11'b00011000100: data <= 32'h3f5330a4;
    11'b00011000101: data <= 32'h41b23bbe;
    11'b00011000110: data <= 32'h3e1c3c70;
    11'b00011000111: data <= 32'hb956a80f;
    11'b00011001000: data <= 32'hbd6bbca5;
    11'b00011001001: data <= 32'hb708bbd5;
    11'b00011001010: data <= 32'h34fdb544;
    11'b00011001011: data <= 32'h30b2baf4;
    11'b00011001100: data <= 32'ha2dac053;
    11'b00011001101: data <= 32'h34ffc003;
    11'b00011001110: data <= 32'h3387319d;
    11'b00011001111: data <= 32'hb9d14039;
    11'b00011010000: data <= 32'hbe083ef4;
    11'b00011010001: data <= 32'hbcb4948a;
    11'b00011010010: data <= 32'hb88bb9e5;
    11'b00011010011: data <= 32'hbad8a566;
    11'b00011010100: data <= 32'hbd4638b7;
    11'b00011010101: data <= 32'hb4d5353b;
    11'b00011010110: data <= 32'h3f6231fb;
    11'b00011010111: data <= 32'h41683ade;
    11'b00011011000: data <= 32'h3ca23dad;
    11'b00011011001: data <= 32'hbaa63bb4;
    11'b00011011010: data <= 32'hbb623102;
    11'b00011011011: data <= 32'h3731a86c;
    11'b00011011100: data <= 32'h3c65b0e9;
    11'b00011011101: data <= 32'h3707bce4;
    11'b00011011110: data <= 32'ha805c0fb;
    11'b00011011111: data <= 32'h3852c01f;
    11'b00011100000: data <= 32'h3c262ddb;
    11'b00011100001: data <= 32'h35ef3e3c;
    11'b00011100010: data <= 32'hba3139cb;
    11'b00011100011: data <= 32'hbcfbbba4;
    11'b00011100100: data <= 32'hbd14bc8b;
    11'b00011100101: data <= 32'hbe782c47;
    11'b00011100110: data <= 32'hbf0738eb;
    11'b00011100111: data <= 32'hb895b05c;
    11'b00011101000: data <= 32'h3d3bb8b5;
    11'b00011101001: data <= 32'h3f153663;
    11'b00011101010: data <= 32'h33bb3f00;
    11'b00011101011: data <= 32'hbcc23fd4;
    11'b00011101100: data <= 32'hb93d3cee;
    11'b00011101101: data <= 32'h3ab03930;
    11'b00011101110: data <= 32'h3c46319c;
    11'b00011101111: data <= 32'h25bdbac1;
    11'b00011110000: data <= 32'hb40dbf4d;
    11'b00011110001: data <= 32'h3c2cbd83;
    11'b00011110010: data <= 32'h4067346c;
    11'b00011110011: data <= 32'h3e683c46;
    11'b00011110100: data <= 32'ha777a5cd;
    11'b00011110101: data <= 32'hbc1bbd6b;
    11'b00011110110: data <= 32'hbcbdbc31;
    11'b00011110111: data <= 32'hbd6130f0;
    11'b00011111000: data <= 32'hbdb92ef9;
    11'b00011111001: data <= 32'hb91bbd21;
    11'b00011111010: data <= 32'h38edbf36;
    11'b00011111011: data <= 32'h3a20b401;
    11'b00011111100: data <= 32'hb7843f22;
    11'b00011111101: data <= 32'hbd4f4089;
    11'b00011111110: data <= 32'hb89c3d9a;
    11'b00011111111: data <= 32'h38183980;
    11'b00100000000: data <= 32'h30bd3783;
    11'b00100000001: data <= 32'hbc0da791;
    11'b00100000010: data <= 32'hb9b6b9c0;
    11'b00100000011: data <= 32'h3d85b85f;
    11'b00100000100: data <= 32'h41de379d;
    11'b00100000101: data <= 32'h40613afa;
    11'b00100000110: data <= 32'h34bca35a;
    11'b00100000111: data <= 32'hb901ba89;
    11'b00100001000: data <= 32'hb64ab50f;
    11'b00100001001: data <= 32'hb4ee3657;
    11'b00100001010: data <= 32'hb963b79a;
    11'b00100001011: data <= 32'hb869c0b4;
    11'b00100001100: data <= 32'h3216c170;
    11'b00100001101: data <= 32'h365fb9e7;
    11'b00100001110: data <= 32'hb5dc3dca;
    11'b00100001111: data <= 32'hbb843ec1;
    11'b00100010000: data <= 32'hb83338d1;
    11'b00100010001: data <= 32'hb21a30a8;
    11'b00100010010: data <= 32'hbc4c38d9;
    11'b00100010011: data <= 32'hc031397b;
    11'b00100010100: data <= 32'hbce92395;
    11'b00100010101: data <= 32'h3d07b460;
    11'b00100010110: data <= 32'h417835c7;
    11'b00100010111: data <= 32'h3f173b58;
    11'b00100011000: data <= 32'h293a3936;
    11'b00100011001: data <= 32'hb424358f;
    11'b00100011010: data <= 32'h389b39d5;
    11'b00100011011: data <= 32'h39b83a6c;
    11'b00100011100: data <= 32'hb0bfb92f;
    11'b00100011101: data <= 32'hb85ec13a;
    11'b00100011110: data <= 32'h31c1c185;
    11'b00100011111: data <= 32'h3af9ba3c;
    11'b00100100000: data <= 32'h38823b79;
    11'b00100100001: data <= 32'hae8d38d8;
    11'b00100100010: data <= 32'hb54bb87f;
    11'b00100100011: data <= 32'hb963b7b3;
    11'b00100100100: data <= 32'hbf11392b;
    11'b00100100101: data <= 32'hc11c3b5a;
    11'b00100100110: data <= 32'hbe0bb008;
    11'b00100100111: data <= 32'h39cfbaea;
    11'b00100101000: data <= 32'h3ef4b21a;
    11'b00100101001: data <= 32'h395f3bbd;
    11'b00100101010: data <= 32'hb8423d94;
    11'b00100101011: data <= 32'hab113d61;
    11'b00100101100: data <= 32'h3c923de1;
    11'b00100101101: data <= 32'h3bfb3ccf;
    11'b00100101110: data <= 32'hb5d2b39b;
    11'b00100101111: data <= 32'hbab9bf92;
    11'b00100110000: data <= 32'h3660bfb2;
    11'b00100110001: data <= 32'h3f0bb66d;
    11'b00100110010: data <= 32'h3ed23820;
    11'b00100110011: data <= 32'h39d8b4c4;
    11'b00100110100: data <= 32'h2415bd0e;
    11'b00100110101: data <= 32'hb81eb8e2;
    11'b00100110110: data <= 32'hbdc33a3f;
    11'b00100110111: data <= 32'hc03a3985;
    11'b00100111000: data <= 32'hbdabbbdc;
    11'b00100111001: data <= 32'h2e9ebfe9;
    11'b00100111010: data <= 32'h38c4bb98;
    11'b00100111011: data <= 32'hb54d3a94;
    11'b00100111100: data <= 32'hbb373e5d;
    11'b00100111101: data <= 32'h298c3dd9;
    11'b00100111110: data <= 32'h3c543dc1;
    11'b00100111111: data <= 32'h36083d87;
    11'b00101000000: data <= 32'hbd223828;
    11'b00101000001: data <= 32'hbdaeb952;
    11'b00101000010: data <= 32'h3824ba87;
    11'b00101000011: data <= 32'h40ae2926;
    11'b00101000100: data <= 32'h407d3539;
    11'b00101000101: data <= 32'h3c20b84c;
    11'b00101000110: data <= 32'h35b7bc24;
    11'b00101000111: data <= 32'h33bea2c5;
    11'b00101001000: data <= 32'hb4c63c90;
    11'b00101001001: data <= 32'hbc6a359a;
    11'b00101001010: data <= 32'hbc57bf79;
    11'b00101001011: data <= 32'hb4a8c1b2;
    11'b00101001100: data <= 32'h9552bdd4;
    11'b00101001101: data <= 32'hb85e37cb;
    11'b00101001110: data <= 32'hb9613c10;
    11'b00101001111: data <= 32'h327b3896;
    11'b00101010000: data <= 32'h391f3964;
    11'b00101010001: data <= 32'hb91a3d25;
    11'b00101010010: data <= 32'hc0a33cbf;
    11'b00101010011: data <= 32'hbff9347b;
    11'b00101010100: data <= 32'h356fb2fa;
    11'b00101010101: data <= 32'h403a2f27;
    11'b00101010110: data <= 32'h3f00348a;
    11'b00101010111: data <= 32'h38bdb080;
    11'b00101011000: data <= 32'h3824ae89;
    11'b00101011001: data <= 32'h3ca13bda;
    11'b00101011010: data <= 32'h3b593e8f;
    11'b00101011011: data <= 32'hb4063489;
    11'b00101011100: data <= 32'hbaeec025;
    11'b00101011101: data <= 32'hb5d0c1a5;
    11'b00101011110: data <= 32'h326fbd70;
    11'b00101011111: data <= 32'h30293090;
    11'b00101100000: data <= 32'h2e8ba4f2;
    11'b00101100001: data <= 32'h3819ba26;
    11'b00101100010: data <= 32'h34f3b463;
    11'b00101100011: data <= 32'hbcf93c5e;
    11'b00101100100: data <= 32'hc1763dd1;
    11'b00101100101: data <= 32'hc05f367d;
    11'b00101100110: data <= 32'hac55b840;
    11'b00101100111: data <= 32'h3c9db5b4;
    11'b00101101000: data <= 32'h37c9329c;
    11'b00101101001: data <= 32'hb49e369e;
    11'b00101101010: data <= 32'h37a03a45;
    11'b00101101011: data <= 32'h3ef13ec3;
    11'b00101101100: data <= 32'h3dd74001;
    11'b00101101101: data <= 32'hb16538f6;
    11'b00101101110: data <= 32'hbc32bd7b;
    11'b00101101111: data <= 32'hb44cbf5e;
    11'b00101110000: data <= 32'h3afcb98f;
    11'b00101110001: data <= 32'h3c88a814;
    11'b00101110010: data <= 32'h3b52bb58;
    11'b00101110011: data <= 32'h3afbbee4;
    11'b00101110100: data <= 32'h3726b9c3;
    11'b00101110101: data <= 32'hbb5d3c55;
    11'b00101110110: data <= 32'hc0563d59;
    11'b00101110111: data <= 32'hbf5ab2de;
    11'b00101111000: data <= 32'hb757bdea;
    11'b00101111001: data <= 32'h2669bc63;
    11'b00101111010: data <= 32'hba191d1a;
    11'b00101111011: data <= 32'hbbee38a0;
    11'b00101111100: data <= 32'h366b3b16;
    11'b00101111101: data <= 32'h3f123e42;
    11'b00101111110: data <= 32'h3c5a3fe2;
    11'b00101111111: data <= 32'hbb293cae;
    11'b00110000000: data <= 32'hbe6ab12d;
    11'b00110000001: data <= 32'hb394b7f4;
    11'b00110000010: data <= 32'h3d7f2dda;
    11'b00110000011: data <= 32'h3e8da50a;
    11'b00110000100: data <= 32'h3c99bced;
    11'b00110000101: data <= 32'h3c39bf03;
    11'b00110000110: data <= 32'h3c1fb587;
    11'b00110000111: data <= 32'h327b3d9c;
    11'b00110001000: data <= 32'hbb783c6a;
    11'b00110001001: data <= 32'hbca4bbdc;
    11'b00110001010: data <= 32'hb90bc096;
    11'b00110001011: data <= 32'hb90abe41;
    11'b00110001100: data <= 32'hbcfcb347;
    11'b00110001101: data <= 32'hbc103041;
    11'b00110001110: data <= 32'h37f42198;
    11'b00110001111: data <= 32'h3dc438c8;
    11'b00110010000: data <= 32'h331e3e2a;
    11'b00110010001: data <= 32'hbf6c3e68;
    11'b00110010010: data <= 32'hc0503a9b;
    11'b00110010011: data <= 32'hb5d73610;
    11'b00110010100: data <= 32'h3cee3737;
    11'b00110010101: data <= 32'h3c9a27da;
    11'b00110010110: data <= 32'h3849bb9f;
    11'b00110010111: data <= 32'h3b45bbfb;
    11'b00110011000: data <= 32'h3eda386c;
    11'b00110011001: data <= 32'h3dcc3f95;
    11'b00110011010: data <= 32'h326b3c21;
    11'b00110011011: data <= 32'hb8f9bcea;
    11'b00110011100: data <= 32'hb89ac08a;
    11'b00110011101: data <= 32'hb852bd4a;
    11'b00110011110: data <= 32'hba34b4d6;
    11'b00110011111: data <= 32'hb5d8b976;
    11'b00110100000: data <= 32'h3a73bd6a;
    11'b00110100001: data <= 32'h3c95b90c;
    11'b00110100010: data <= 32'hb6283c04;
    11'b00110100011: data <= 32'hc0873ed6;
    11'b00110100100: data <= 32'hc07b3c37;
    11'b00110100101: data <= 32'hb86234c1;
    11'b00110100110: data <= 32'h377a308b;
    11'b00110100111: data <= 32'hb037a8ff;
    11'b00110101000: data <= 32'hb8f2b770;
    11'b00110101001: data <= 32'h381bb0bb;
    11'b00110101010: data <= 32'h40353d03;
    11'b00110101011: data <= 32'h402a405e;
    11'b00110101100: data <= 32'h38503cc7;
    11'b00110101101: data <= 32'hb8d6b98d;
    11'b00110101110: data <= 32'hb744bd19;
    11'b00110101111: data <= 32'h29a4b666;
    11'b00110110000: data <= 32'h30f4afdf;
    11'b00110110001: data <= 32'h36dbbd84;
    11'b00110110010: data <= 32'h3c81c0c8;
    11'b00110110011: data <= 32'h3ca4bd6a;
    11'b00110110100: data <= 32'hb2573a08;
    11'b00110110101: data <= 32'hbec43e27;
    11'b00110110110: data <= 32'hbea03844;
    11'b00110110111: data <= 32'hb8c8b855;
    11'b00110111000: data <= 32'hb741b87f;
    11'b00110111001: data <= 32'hbdd6b33b;
    11'b00110111010: data <= 32'hbe76b347;
    11'b00110111011: data <= 32'h310d2b76;
    11'b00110111100: data <= 32'h401b3c81;
    11'b00110111101: data <= 32'h3f443fcf;
    11'b00110111110: data <= 32'ha9a13db6;
    11'b00110111111: data <= 32'hbc6234f3;
    11'b00111000000: data <= 32'hb6bd30a7;
    11'b00111000001: data <= 32'h3898398d;
    11'b00111000010: data <= 32'h39d83279;
    11'b00111000011: data <= 32'h395dbe54;
    11'b00111000100: data <= 32'h3c98c10f;
    11'b00111000101: data <= 32'h3ddbbca0;
    11'b00111000110: data <= 32'h39d23bd1;
    11'b00111000111: data <= 32'hb63c3d37;
    11'b00111001000: data <= 32'hb955b34f;
    11'b00111001001: data <= 32'hb6e4bd94;
    11'b00111001010: data <= 32'hbbc8bc29;
    11'b00111001011: data <= 32'hc01db571;
    11'b00111001100: data <= 32'hbf6bb6fc;
    11'b00111001101: data <= 32'h2f91b911;
    11'b00111001110: data <= 32'h3edf2e9d;
    11'b00111001111: data <= 32'h3bdf3cde;
    11'b00111010000: data <= 32'hbc0a3e07;
    11'b00111010001: data <= 32'hbea43c91;
    11'b00111010010: data <= 32'hb7813c8f;
    11'b00111010011: data <= 32'h38f93d38;
    11'b00111010100: data <= 32'h368436ea;
    11'b00111010101: data <= 32'h23f4bd1d;
    11'b00111010110: data <= 32'h39bdbf52;
    11'b00111010111: data <= 32'h3f2db494;
    11'b00111011000: data <= 32'h3f393de4;
    11'b00111011001: data <= 32'h3aeb3cbc;
    11'b00111011010: data <= 32'h310ab8f5;
    11'b00111011011: data <= 32'hb0ccbe0e;
    11'b00111011100: data <= 32'hbab4ba32;
    11'b00111011101: data <= 32'hbea5b12e;
    11'b00111011110: data <= 32'hbd13bb52;
    11'b00111011111: data <= 32'h36a4bf4a;
    11'b00111100000: data <= 32'h3d94bcfa;
    11'b00111100001: data <= 32'h345535e1;
    11'b00111100010: data <= 32'hbe2b3d62;
    11'b00111100011: data <= 32'hbef13d35;
    11'b00111100100: data <= 32'hb6f93c9d;
    11'b00111100101: data <= 32'h31633c6c;
    11'b00111100110: data <= 32'hb99b366a;
    11'b00111100111: data <= 32'hbd02ba36;
    11'b00111101000: data <= 32'h9ce0bb49;
    11'b00111101001: data <= 32'h3f883824;
    11'b00111101010: data <= 32'h40b33f15;
    11'b00111101011: data <= 32'h3d443cad;
    11'b00111101100: data <= 32'h3553b5da;
    11'b00111101101: data <= 32'h2a09b981;
    11'b00111101110: data <= 32'hb3cd3409;
    11'b00111101111: data <= 32'hb991358a;
    11'b00111110000: data <= 32'hb656bd26;
    11'b00111110001: data <= 32'h3a0fc181;
    11'b00111110010: data <= 32'h3d17c030;
    11'b00111110011: data <= 32'h32b1ada3;
    11'b00111110100: data <= 32'hbc8a3c37;
    11'b00111110101: data <= 32'hbc413a1f;
    11'b00111110110: data <= 32'hb15034f9;
    11'b00111110111: data <= 32'hb6b535a9;
    11'b00111111000: data <= 32'hbfa431fc;
    11'b00111111001: data <= 32'hc0c8b70b;
    11'b00111111010: data <= 32'hb8e0b7db;
    11'b00111111011: data <= 32'h3ea8386e;
    11'b00111111100: data <= 32'h401b3de4;
    11'b00111111101: data <= 32'h3a143c69;
    11'b00111111110: data <= 32'hb15c34e0;
    11'b00111111111: data <= 32'h2bd738d8;
    11'b01000000000: data <= 32'h35af3dfe;
    11'b01000000001: data <= 32'h2b6b3bab;
    11'b01000000010: data <= 32'h1c63bd1f;
    11'b01000000011: data <= 32'h39f0c1b4;
    11'b01000000100: data <= 32'h3d3bbfd0;
    11'b01000000101: data <= 32'h3a7d2e50;
    11'b01000000110: data <= 32'h28433a8b;
    11'b01000000111: data <= 32'h2d48a9d3;
    11'b01000001000: data <= 32'h3512b97d;
    11'b01000001001: data <= 32'hb98bb460;
    11'b01000001010: data <= 32'hc0e92d59;
    11'b01000001011: data <= 32'hc16eb6b2;
    11'b01000001100: data <= 32'hb9e1baff;
    11'b01000001101: data <= 32'h3d30b53d;
    11'b01000001110: data <= 32'h3cbb38b3;
    11'b01000001111: data <= 32'hb5163acc;
    11'b01000010000: data <= 32'hbaea3ae5;
    11'b01000010001: data <= 32'h1ac13e2a;
    11'b01000010010: data <= 32'h38c14073;
    11'b01000010011: data <= 32'h255f3d4f;
    11'b01000010100: data <= 32'hb801bb47;
    11'b01000010101: data <= 32'h31afc03c;
    11'b01000010110: data <= 32'h3d35bc04;
    11'b01000010111: data <= 32'h3e5f39a4;
    11'b01000011000: data <= 32'h3ce239c2;
    11'b01000011001: data <= 32'h3c36b8c0;
    11'b01000011010: data <= 32'h3a53bc45;
    11'b01000011011: data <= 32'hb73ab149;
    11'b01000011100: data <= 32'hc00f35ec;
    11'b01000011101: data <= 32'hc02cb895;
    11'b01000011110: data <= 32'hb5bbbf08;
    11'b01000011111: data <= 32'h3bfdbe66;
    11'b01000100000: data <= 32'h3577b6df;
    11'b01000100001: data <= 32'hbc5b3720;
    11'b01000100010: data <= 32'hbc6a3b01;
    11'b01000100011: data <= 32'h2f6e3e1a;
    11'b01000100100: data <= 32'h3716400c;
    11'b01000100101: data <= 32'hba3b3d06;
    11'b01000100110: data <= 32'hbebab6ca;
    11'b01000100111: data <= 32'hb9cabc5f;
    11'b01000101000: data <= 32'h3c6f2408;
    11'b01000101001: data <= 32'h3fce3caf;
    11'b01000101010: data <= 32'h3e94393d;
    11'b01000101011: data <= 32'h3d12b8eb;
    11'b01000101100: data <= 32'h3bfeb85e;
    11'b01000101101: data <= 32'h309b3a1c;
    11'b01000101110: data <= 32'hbbd63c3b;
    11'b01000101111: data <= 32'hbc18b919;
    11'b01000110000: data <= 32'h30dec0f1;
    11'b01000110001: data <= 32'h3ad3c0d8;
    11'b01000110010: data <= 32'h283fbbc0;
    11'b01000110011: data <= 32'hbbd82d63;
    11'b01000110100: data <= 32'hb85a34f5;
    11'b01000110101: data <= 32'h387338ec;
    11'b01000110110: data <= 32'h31a73c75;
    11'b01000110111: data <= 32'hbefe3b14;
    11'b01000111000: data <= 32'hc196ad89;
    11'b01000111001: data <= 32'hbdcdb746;
    11'b01000111010: data <= 32'h3a1d3584;
    11'b01000111011: data <= 32'h3e613c03;
    11'b01000111100: data <= 32'h3c2236f9;
    11'b01000111101: data <= 32'h3934b44a;
    11'b01000111110: data <= 32'h3b0737e0;
    11'b01000111111: data <= 32'h39db3fec;
    11'b01001000000: data <= 32'ha8773f4d;
    11'b01001000001: data <= 32'hb569b73a;
    11'b01001000010: data <= 32'h3499c0f2;
    11'b01001000011: data <= 32'h3a17c079;
    11'b01001000100: data <= 32'h3512b9ac;
    11'b01001000101: data <= 32'had28aac6;
    11'b01001000110: data <= 32'h388bb7d5;
    11'b01001000111: data <= 32'h3ce0b860;
    11'b01001001000: data <= 32'h300b32e7;
    11'b01001001001: data <= 32'hc05638e7;
    11'b01001001010: data <= 32'hc22c27bc;
    11'b01001001011: data <= 32'hbe35b845;
    11'b01001001100: data <= 32'h3733b419;
    11'b01001001101: data <= 32'h39cc3141;
    11'b01001001110: data <= 32'hb204a1fd;
    11'b01001001111: data <= 32'hb4c42772;
    11'b01001010000: data <= 32'h39243d1b;
    11'b01001010001: data <= 32'h3c244162;
    11'b01001010010: data <= 32'h32dc4070;
    11'b01001010011: data <= 32'hb86cad4d;
    11'b01001010100: data <= 32'hb2bcbee6;
    11'b01001010101: data <= 32'h387dbca8;
    11'b01001010110: data <= 32'h3a802fe3;
    11'b01001010111: data <= 32'h3b762694;
    11'b01001011000: data <= 32'h3e25bc50;
    11'b01001011001: data <= 32'h3f14bcc7;
    11'b01001011010: data <= 32'h36b426c4;
    11'b01001011011: data <= 32'hbed63a75;
    11'b01001011100: data <= 32'hc0b52b5e;
    11'b01001011101: data <= 32'hbbdbbc75;
    11'b01001011110: data <= 32'h350cbd53;
    11'b01001011111: data <= 32'hb08ebade;
    11'b01001100000: data <= 32'hbcd3b84f;
    11'b01001100001: data <= 32'hbab8abfd;
    11'b01001100010: data <= 32'h39173cd4;
    11'b01001100011: data <= 32'h3c2e40d3;
    11'b01001100100: data <= 32'hb4733fff;
    11'b01001100101: data <= 32'hbe12342d;
    11'b01001100110: data <= 32'hbc77b974;
    11'b01001100111: data <= 32'h32ab2d85;
    11'b01001101000: data <= 32'h3c103b22;
    11'b01001101001: data <= 32'h3d202e9e;
    11'b01001101010: data <= 32'h3ecebcf1;
    11'b01001101011: data <= 32'h3f85bbd6;
    11'b01001101100: data <= 32'h3b4239c2;
    11'b01001101101: data <= 32'hb9223df6;
    11'b01001101110: data <= 32'hbc52319b;
    11'b01001101111: data <= 32'hb18cbe86;
    11'b01001110000: data <= 32'h3550c01e;
    11'b01001110001: data <= 32'hb882bd7f;
    11'b01001110010: data <= 32'hbd9bbadf;
    11'b01001110011: data <= 32'hb846b884;
    11'b01001110100: data <= 32'h3c38346d;
    11'b01001110101: data <= 32'h3bc23d42;
    11'b01001110110: data <= 32'hbc133d5f;
    11'b01001110111: data <= 32'hc10636cd;
    11'b01001111000: data <= 32'hbf5f2a1f;
    11'b01001111001: data <= 32'hb0de39b8;
    11'b01001111010: data <= 32'h39613c00;
    11'b01001111011: data <= 32'h3924ac7d;
    11'b01001111100: data <= 32'h3b64bc52;
    11'b01001111101: data <= 32'h3e02b22e;
    11'b01001111110: data <= 32'h3d483f37;
    11'b01001111111: data <= 32'h3604408c;
    11'b01010000000: data <= 32'hae6a36d9;
    11'b01010000001: data <= 32'h3424be64;
    11'b01010000010: data <= 32'h3508bf59;
    11'b01010000011: data <= 32'hb768bbe5;
    11'b01010000100: data <= 32'hba2cba3b;
    11'b01010000101: data <= 32'h36cebccf;
    11'b01010000110: data <= 32'h3efabb90;
    11'b01010000111: data <= 32'h3c1e302d;
    11'b01010001000: data <= 32'hbd6f3a0e;
    11'b01010001001: data <= 32'hc18536fd;
    11'b01010001010: data <= 32'hbf67306e;
    11'b01010001011: data <= 32'hb4c43668;
    11'b01010001100: data <= 32'habd63565;
    11'b01010001101: data <= 32'hb90bb85d;
    11'b01010001110: data <= 32'hb4b9bb6a;
    11'b01010001111: data <= 32'h3b8f378a;
    11'b01010010000: data <= 32'h3df840ec;
    11'b01010010001: data <= 32'h3a384138;
    11'b01010010010: data <= 32'ha3a03976;
    11'b01010010011: data <= 32'ha83bbb9c;
    11'b01010010100: data <= 32'h2e3ab9b7;
    11'b01010010101: data <= 32'hb0522e29;
    11'b01010010110: data <= 32'h2d91b625;
    11'b01010010111: data <= 32'h3d53be90;
    11'b01010011000: data <= 32'h408bbee9;
    11'b01010011001: data <= 32'h3d0eb5e5;
    11'b01010011010: data <= 32'hbbb939b3;
    11'b01010011011: data <= 32'hbfed375a;
    11'b01010011100: data <= 32'hbc38b431;
    11'b01010011101: data <= 32'hb041b7cf;
    11'b01010011110: data <= 32'hba2bb8e5;
    11'b01010011111: data <= 32'hbf15bc53;
    11'b01010100000: data <= 32'hbc9dbc0f;
    11'b01010100001: data <= 32'h395a36e4;
    11'b01010100010: data <= 32'h3ddf4046;
    11'b01010100011: data <= 32'h377c4065;
    11'b01010100100: data <= 32'hba1b3a0a;
    11'b01010100101: data <= 32'hbac5abf0;
    11'b01010100110: data <= 32'hb492392f;
    11'b01010100111: data <= 32'h255f3cbd;
    11'b01010101000: data <= 32'h36d4a18e;
    11'b01010101001: data <= 32'h3dd8bef1;
    11'b01010101010: data <= 32'h4076bec5;
    11'b01010101011: data <= 32'h3e142d4b;
    11'b01010101100: data <= 32'ha9163d1c;
    11'b01010101101: data <= 32'hb8d238ec;
    11'b01010101110: data <= 32'h2c99b984;
    11'b01010101111: data <= 32'h325abcad;
    11'b01010110000: data <= 32'hbc6bbc63;
    11'b01010110001: data <= 32'hc047bd2f;
    11'b01010110010: data <= 32'hbc75bd55;
    11'b01010110011: data <= 32'h3b81b604;
    11'b01010110100: data <= 32'h3db63b94;
    11'b01010110101: data <= 32'hb0ea3cee;
    11'b01010110110: data <= 32'hbeb638c0;
    11'b01010110111: data <= 32'hbe2c387a;
    11'b01010111000: data <= 32'hb8ae3dca;
    11'b01010111001: data <= 32'hb22b3e56;
    11'b01010111010: data <= 32'haf319004;
    11'b01010111011: data <= 32'h38d3be68;
    11'b01010111100: data <= 32'h3e44bc2f;
    11'b01010111101: data <= 32'h3e713c37;
    11'b01010111110: data <= 32'h3ad8400d;
    11'b01010111111: data <= 32'h385b3ac1;
    11'b01011000000: data <= 32'h3a8fb9db;
    11'b01011000001: data <= 32'h3670bc13;
    11'b01011000010: data <= 32'hbc07b927;
    11'b01011000011: data <= 32'hbeaabbb4;
    11'b01011000100: data <= 32'hb4c7bea9;
    11'b01011000101: data <= 32'h3e55bde0;
    11'b01011000110: data <= 32'h3df8b663;
    11'b01011000111: data <= 32'hb82b34f9;
    11'b01011001000: data <= 32'hbfe1358d;
    11'b01011001001: data <= 32'hbe00390c;
    11'b01011001010: data <= 32'hb8273d36;
    11'b01011001011: data <= 32'hb9373c65;
    11'b01011001100: data <= 32'hbd09b69c;
    11'b01011001101: data <= 32'hba29bde4;
    11'b01011001110: data <= 32'h394eb655;
    11'b01011001111: data <= 32'h3df73eeb;
    11'b01011010000: data <= 32'h3cdb40a8;
    11'b01011010001: data <= 32'h3a7c3b76;
    11'b01011010010: data <= 32'h39f3b522;
    11'b01011010011: data <= 32'h3469a329;
    11'b01011010100: data <= 32'hb9b338a8;
    11'b01011010101: data <= 32'hbaddb328;
    11'b01011010110: data <= 32'h38cfbf2d;
    11'b01011010111: data <= 32'h402ec060;
    11'b01011011000: data <= 32'h3e6cbc59;
    11'b01011011001: data <= 32'hb51d21fe;
    11'b01011011010: data <= 32'hbd2f33bc;
    11'b01011011011: data <= 32'hb89d3436;
    11'b01011011100: data <= 32'ha60b37f3;
    11'b01011011101: data <= 32'hbc2e31ea;
    11'b01011011110: data <= 32'hc0a4bb81;
    11'b01011011111: data <= 32'hbf4bbdf0;
    11'b01011100000: data <= 32'h2e2eb499;
    11'b01011100001: data <= 32'h3d313e00;
    11'b01011100010: data <= 32'h3b6a3f39;
    11'b01011100011: data <= 32'h31883997;
    11'b01011100100: data <= 32'h94663420;
    11'b01011100101: data <= 32'hae273d0c;
    11'b01011100110: data <= 32'hb8273f7a;
    11'b01011100111: data <= 32'hb69a378b;
    11'b01011101000: data <= 32'h3a80beb7;
    11'b01011101001: data <= 32'h3fdcc051;
    11'b01011101010: data <= 32'h3e5bba2b;
    11'b01011101011: data <= 32'h34fb377e;
    11'b01011101100: data <= 32'h9e0935fc;
    11'b01011101101: data <= 32'h3a02b189;
    11'b01011101110: data <= 32'h3939b3ed;
    11'b01011101111: data <= 32'hbc89b5e7;
    11'b01011110000: data <= 32'hc15dbc63;
    11'b01011110001: data <= 32'hbfc5be4b;
    11'b01011110010: data <= 32'h32e0ba96;
    11'b01011110011: data <= 32'h3cd63665;
    11'b01011110100: data <= 32'h3505392a;
    11'b01011110101: data <= 32'hba2231bc;
    11'b01011110110: data <= 32'hb9fe38e0;
    11'b01011110111: data <= 32'hb5d64016;
    11'b01011111000: data <= 32'hb86840e6;
    11'b01011111001: data <= 32'hb9b1396b;
    11'b01011111010: data <= 32'h2a02bddc;
    11'b01011111011: data <= 32'h3c7bbe1d;
    11'b01011111100: data <= 32'h3d493216;
    11'b01011111101: data <= 32'h3b5b3cfc;
    11'b01011111110: data <= 32'h3c7438b9;
    11'b01011111111: data <= 32'h3ecfb5a1;
    11'b01100000000: data <= 32'h3c64b4d9;
    11'b01100000001: data <= 32'hbb61a12e;
    11'b01100000010: data <= 32'hc073b8db;
    11'b01100000011: data <= 32'hbcacbe3e;
    11'b01100000100: data <= 32'h3ae3be7c;
    11'b01100000101: data <= 32'h3d14bb49;
    11'b01100000110: data <= 32'hb0cfb7f6;
    11'b01100000111: data <= 32'hbce9b5a7;
    11'b01100001000: data <= 32'hba66383b;
    11'b01100001001: data <= 32'hb1863fa9;
    11'b01100001010: data <= 32'hb98b4015;
    11'b01100001011: data <= 32'hbe4434c6;
    11'b01100001100: data <= 32'hbd21bd51;
    11'b01100001101: data <= 32'ha416ba80;
    11'b01100001110: data <= 32'h3b083c04;
    11'b01100001111: data <= 32'h3c5b3e8f;
    11'b01100010000: data <= 32'h3d9438ab;
    11'b01100010001: data <= 32'h3ef5b312;
    11'b01100010010: data <= 32'h3c3136c6;
    11'b01100010011: data <= 32'hb8e03ca8;
    11'b01100010100: data <= 32'hbd8135d8;
    11'b01100010101: data <= 32'hb134bd5d;
    11'b01100010110: data <= 32'h3dd3c03d;
    11'b01100010111: data <= 32'h3d46be72;
    11'b01100011000: data <= 32'hb218bb97;
    11'b01100011001: data <= 32'hba85b8b0;
    11'b01100011010: data <= 32'h2c202fba;
    11'b01100011011: data <= 32'h385e3c5a;
    11'b01100011100: data <= 32'hb9d33c37;
    11'b01100011101: data <= 32'hc0c5b4e4;
    11'b01100011110: data <= 32'hc0b1bd36;
    11'b01100011111: data <= 32'hba2ab802;
    11'b01100100000: data <= 32'h38083c10;
    11'b01100100001: data <= 32'h39d93cbf;
    11'b01100100010: data <= 32'h3a0230a5;
    11'b01100100011: data <= 32'h3bae1a32;
    11'b01100100100: data <= 32'h38ec3dc7;
    11'b01100100101: data <= 32'hb65b40eb;
    11'b01100100110: data <= 32'hba1f3d1c;
    11'b01100100111: data <= 32'h3458bbf3;
    11'b01100101000: data <= 32'h3da6bff2;
    11'b01100101001: data <= 32'h3c7fbd34;
    11'b01100101010: data <= 32'h2e59b800;
    11'b01100101011: data <= 32'h32deb6c7;
    11'b01100101100: data <= 32'h3d96b533;
    11'b01100101101: data <= 32'h3dd832c8;
    11'b01100101110: data <= 32'hb85634c6;
    11'b01100101111: data <= 32'hc138b87a;
    11'b01100110000: data <= 32'hc0f5bcfd;
    11'b01100110001: data <= 32'hb9a3b9bd;
    11'b01100110010: data <= 32'h367731a5;
    11'b01100110011: data <= 32'h2ebc2702;
    11'b01100110100: data <= 32'hb4a1b904;
    11'b01100110101: data <= 32'h289529e0;
    11'b01100110110: data <= 32'h33bc4020;
    11'b01100110111: data <= 32'hb51f4220;
    11'b01100111000: data <= 32'hba2f3e53;
    11'b01100111001: data <= 32'hb379b9c3;
    11'b01100111010: data <= 32'h38a6bd51;
    11'b01100111011: data <= 32'h38cfb434;
    11'b01100111100: data <= 32'h360136ca;
    11'b01100111101: data <= 32'h3c9aae84;
    11'b01100111110: data <= 32'h40c4b8a4;
    11'b01100111111: data <= 32'h401aae92;
    11'b01101000000: data <= 32'hb3013666;
    11'b01101000001: data <= 32'hc037ae94;
    11'b01101000010: data <= 32'hbe99bbee;
    11'b01101000011: data <= 32'h2ad0bcaf;
    11'b01101000100: data <= 32'h3879bb77;
    11'b01101000101: data <= 32'hb695bca4;
    11'b01101000110: data <= 32'hbbd4bd64;
    11'b01101000111: data <= 32'hb440b255;
    11'b01101001000: data <= 32'h360f3f77;
    11'b01101001001: data <= 32'hb3c8413e;
    11'b01101001010: data <= 32'hbd233c86;
    11'b01101001011: data <= 32'hbd64b944;
    11'b01101001100: data <= 32'hb8d2b898;
    11'b01101001101: data <= 32'hac4839ff;
    11'b01101001110: data <= 32'h35533c3c;
    11'b01101001111: data <= 32'h3d5fa817;
    11'b01101010000: data <= 32'h40d2b91b;
    11'b01101010001: data <= 32'h3fe934a5;
    11'b01101010010: data <= 32'h2a873d64;
    11'b01101010011: data <= 32'hbce73b4b;
    11'b01101010100: data <= 32'hb786b82a;
    11'b01101010101: data <= 32'h3b04bda9;
    11'b01101010110: data <= 32'h399dbe19;
    11'b01101010111: data <= 32'hb8dfbe83;
    11'b01101011000: data <= 32'hbb0fbe72;
    11'b01101011001: data <= 32'h35d1b8d3;
    11'b01101011010: data <= 32'h3c823c06;
    11'b01101011011: data <= 32'ha4613df3;
    11'b01101011100: data <= 32'hbf44350d;
    11'b01101011101: data <= 32'hc090b9e6;
    11'b01101011110: data <= 32'hbd96b051;
    11'b01101011111: data <= 32'hb83c3c3e;
    11'b01101100000: data <= 32'hac833acb;
    11'b01101100001: data <= 32'h3948b7b5;
    11'b01101100010: data <= 32'h3e0eb962;
    11'b01101100011: data <= 32'h3d713c05;
    11'b01101100100: data <= 32'h30ee40ff;
    11'b01101100101: data <= 32'hb8173f87;
    11'b01101100110: data <= 32'h33e0a83b;
    11'b01101100111: data <= 32'h3c58bcbd;
    11'b01101101000: data <= 32'h3828bca8;
    11'b01101101001: data <= 32'hb887bc60;
    11'b01101101010: data <= 32'hb166bd36;
    11'b01101101011: data <= 32'h3e26bb96;
    11'b01101101100: data <= 32'h40392a26;
    11'b01101101101: data <= 32'h35aa377c;
    11'b01101101110: data <= 32'hbf96b25a;
    11'b01101101111: data <= 32'hc0b4b9c5;
    11'b01101110000: data <= 32'hbd1eafe6;
    11'b01101110001: data <= 32'hb8413857;
    11'b01101110010: data <= 32'hb8f2b064;
    11'b01101110011: data <= 32'hb72dbd50;
    11'b01101110100: data <= 32'h3591bacb;
    11'b01101110101: data <= 32'h39ca3dc0;
    11'b01101110110: data <= 32'h313f420f;
    11'b01101110111: data <= 32'hb50a4056;
    11'b01101111000: data <= 32'h2c153256;
    11'b01101111001: data <= 32'h371eb894;
    11'b01101111010: data <= 32'hacb2ac29;
    11'b01101111011: data <= 32'hb84429ff;
    11'b01101111100: data <= 32'h3861b9ce;
    11'b01101111101: data <= 32'h40e2bc75;
    11'b01101111110: data <= 32'h4170b71c;
    11'b01101111111: data <= 32'h398a33f3;
    11'b01110000000: data <= 32'hbd9829e7;
    11'b01110000001: data <= 32'hbddcb693;
    11'b01110000010: data <= 32'hb55bb526;
    11'b01110000011: data <= 32'hb082b51c;
    11'b01110000100: data <= 32'hbc24bcf1;
    11'b01110000101: data <= 32'hbd2ac033;
    11'b01110000110: data <= 32'hb44ebca8;
    11'b01110000111: data <= 32'h39023cd3;
    11'b01110001000: data <= 32'h3455410f;
    11'b01110001001: data <= 32'hb8903e42;
    11'b01110001010: data <= 32'hba3d2aee;
    11'b01110001011: data <= 32'hb91a2d61;
    11'b01110001100: data <= 32'hba893c54;
    11'b01110001101: data <= 32'hb9993bea;
    11'b01110001110: data <= 32'h3952b66f;
    11'b01110001111: data <= 32'h40d5bcb1;
    11'b01110010000: data <= 32'h4110b4c4;
    11'b01110010001: data <= 32'h3a5e3b45;
    11'b01110010010: data <= 32'hb8d33b8a;
    11'b01110010011: data <= 32'hb14130cf;
    11'b01110010100: data <= 32'h3a49b655;
    11'b01110010101: data <= 32'h344cba61;
    11'b01110010110: data <= 32'hbcd2be9d;
    11'b01110010111: data <= 32'hbdb5c096;
    11'b01110011000: data <= 32'h2b7abdd0;
    11'b01110011001: data <= 32'h3cef369b;
    11'b01110011010: data <= 32'h38b63d24;
    11'b01110011011: data <= 32'hbb30377d;
    11'b01110011100: data <= 32'hbe42b4c1;
    11'b01110011101: data <= 32'hbd8a3791;
    11'b01110011110: data <= 32'hbd073e71;
    11'b01110011111: data <= 32'hbc2b3c5d;
    11'b01110100000: data <= 32'h25f4b97b;
    11'b01110100001: data <= 32'h3db0bd29;
    11'b01110100010: data <= 32'h3ea0322a;
    11'b01110100011: data <= 32'h390d3f83;
    11'b01110100100: data <= 32'h299d3f74;
    11'b01110100101: data <= 32'h3a0d3945;
    11'b01110100110: data <= 32'h3d45b157;
    11'b01110100111: data <= 32'h347eb729;
    11'b01110101000: data <= 32'hbce8bc25;
    11'b01110101001: data <= 32'hbb98bf0b;
    11'b01110101010: data <= 32'h3c1abe31;
    11'b01110101011: data <= 32'h4054b783;
    11'b01110101100: data <= 32'h3c0f2cbe;
    11'b01110101101: data <= 32'hbb66b611;
    11'b01110101110: data <= 32'hbe75b808;
    11'b01110101111: data <= 32'hbccc3836;
    11'b01110110000: data <= 32'hbc513d55;
    11'b01110110001: data <= 32'hbd7d355f;
    11'b01110110010: data <= 32'hbc0abddd;
    11'b01110110011: data <= 32'h2cf1be2e;
    11'b01110110100: data <= 32'h39773830;
    11'b01110110101: data <= 32'h364440b6;
    11'b01110110110: data <= 32'h34204031;
    11'b01110110111: data <= 32'h3a893a11;
    11'b01110111000: data <= 32'h3b773454;
    11'b01110111001: data <= 32'hb34538ae;
    11'b01110111010: data <= 32'hbd243446;
    11'b01110111011: data <= 32'hb5f4bad4;
    11'b01110111100: data <= 32'h3f67bdc8;
    11'b01110111101: data <= 32'h4176bba4;
    11'b01110111110: data <= 32'h3d16b636;
    11'b01110111111: data <= 32'hb86cb6b0;
    11'b01111000000: data <= 32'hba36b4e6;
    11'b01111000001: data <= 32'haee336c6;
    11'b01111000010: data <= 32'hb6053921;
    11'b01111000011: data <= 32'hbe0fb942;
    11'b01111000100: data <= 32'hbf4dc06a;
    11'b01111000101: data <= 32'hba3dbf4e;
    11'b01111000110: data <= 32'h346735de;
    11'b01111000111: data <= 32'h35a13f8e;
    11'b01111001000: data <= 32'h2dc63d75;
    11'b01111001001: data <= 32'h31643548;
    11'b01111001010: data <= 32'ha44a394a;
    11'b01111001011: data <= 32'hbb973ec6;
    11'b01111001100: data <= 32'hbdda3dc7;
    11'b01111001101: data <= 32'hb356b252;
    11'b01111001110: data <= 32'h3f5bbd49;
    11'b01111001111: data <= 32'h40dfbb0a;
    11'b01111010000: data <= 32'h3c832b58;
    11'b01111010001: data <= 32'h99523506;
    11'b01111010010: data <= 32'h37b63356;
    11'b01111010011: data <= 32'h3cf73657;
    11'b01111010100: data <= 32'h361831ee;
    11'b01111010101: data <= 32'hbde1bc4b;
    11'b01111010110: data <= 32'hc006c0a5;
    11'b01111010111: data <= 32'hb973bfa7;
    11'b01111011000: data <= 32'h3979b2bb;
    11'b01111011001: data <= 32'h3907397b;
    11'b01111011010: data <= 32'hb1582a08;
    11'b01111011011: data <= 32'hb869b601;
    11'b01111011100: data <= 32'hb9f23a7d;
    11'b01111011101: data <= 32'hbd594083;
    11'b01111011110: data <= 32'hbea03f26;
    11'b01111011111: data <= 32'hb988b3e4;
    11'b01111100000: data <= 32'h3b0fbd7c;
    11'b01111100001: data <= 32'h3d6cb78e;
    11'b01111100010: data <= 32'h38e73b66;
    11'b01111100011: data <= 32'h36413cc6;
    11'b01111100100: data <= 32'h3db139ad;
    11'b01111100101: data <= 32'h400d383c;
    11'b01111100110: data <= 32'h394d365a;
    11'b01111100111: data <= 32'hbd92b7da;
    11'b01111101000: data <= 32'hbe7abe6e;
    11'b01111101001: data <= 32'h30e7beb2;
    11'b01111101010: data <= 32'h3e31baad;
    11'b01111101011: data <= 32'h3c29b84c;
    11'b01111101100: data <= 32'hb3afbc41;
    11'b01111101101: data <= 32'hb98fbb18;
    11'b01111101110: data <= 32'hb8b539de;
    11'b01111101111: data <= 32'hbc07401e;
    11'b01111110000: data <= 32'hbeba3cc5;
    11'b01111110001: data <= 32'hbde3bb74;
    11'b01111110010: data <= 32'hb771be77;
    11'b01111110011: data <= 32'h2f2bb04b;
    11'b01111110100: data <= 32'h28d03dd2;
    11'b01111110101: data <= 32'h370b3dce;
    11'b01111110110: data <= 32'h3e3d3986;
    11'b01111110111: data <= 32'h3f5239a5;
    11'b01111111000: data <= 32'h348b3cc7;
    11'b01111111001: data <= 32'hbdbf3a7a;
    11'b01111111010: data <= 32'hbc43b6e7;
    11'b01111111011: data <= 32'h3bf1bcdc;
    11'b01111111100: data <= 32'h4043bc7f;
    11'b01111111101: data <= 32'h3cd9bc46;
    11'b01111111110: data <= 32'had33bd48;
    11'b01111111111: data <= 32'hac36badd;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    