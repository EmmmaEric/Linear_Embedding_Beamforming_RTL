
module memory_rom_12(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbb173d45;
    11'b00000000001: data <= 32'hb6fb39b4;
    11'b00000000010: data <= 32'h38dfba52;
    11'b00000000011: data <= 32'h3eb0bacd;
    11'b00000000100: data <= 32'h3ddc3b77;
    11'b00000000101: data <= 32'h335540b7;
    11'b00000000110: data <= 32'hb4683f12;
    11'b00000000111: data <= 32'h386c3086;
    11'b00000001000: data <= 32'h3c76ba2e;
    11'b00000001001: data <= 32'h3190bb55;
    11'b00000001010: data <= 32'hbba9bcf7;
    11'b00000001011: data <= 32'hb4b6be75;
    11'b00000001100: data <= 32'h3e61bc73;
    11'b00000001101: data <= 32'h4046995a;
    11'b00000001110: data <= 32'h36593577;
    11'b00000001111: data <= 32'hbe9cb4f7;
    11'b00000010000: data <= 32'hc00db856;
    11'b00000010001: data <= 32'hbcf23525;
    11'b00000010010: data <= 32'hbaea3ae4;
    11'b00000010011: data <= 32'hbbdcb23e;
    11'b00000010100: data <= 32'hb849be49;
    11'b00000010101: data <= 32'h36febbf8;
    11'b00000010110: data <= 32'h3a163d6b;
    11'b00000010111: data <= 32'h32de41b5;
    11'b00000011000: data <= 32'ha9904008;
    11'b00000011001: data <= 32'h372b3593;
    11'b00000011010: data <= 32'h3878b122;
    11'b00000011011: data <= 32'hb5ba32c0;
    11'b00000011100: data <= 32'hbb35aa28;
    11'b00000011101: data <= 32'h3680bbdf;
    11'b00000011110: data <= 32'h40eabd0b;
    11'b00000011111: data <= 32'h4163b84b;
    11'b00000100000: data <= 32'h39a128a4;
    11'b00000100001: data <= 32'hbca0b0f0;
    11'b00000100010: data <= 32'hbc73b493;
    11'b00000100011: data <= 32'hb3fd2f5a;
    11'b00000100100: data <= 32'hb6f2274b;
    11'b00000100101: data <= 32'hbd8fbcf8;
    11'b00000100110: data <= 32'hbdadc092;
    11'b00000100111: data <= 32'hb437bd16;
    11'b00000101000: data <= 32'h389a3c86;
    11'b00000101001: data <= 32'h346040a8;
    11'b00000101010: data <= 32'hb4a53d7d;
    11'b00000101011: data <= 32'hb58b3184;
    11'b00000101100: data <= 32'hb75d37e3;
    11'b00000101101: data <= 32'hbc2c3d96;
    11'b00000101110: data <= 32'hbc1b3bbc;
    11'b00000101111: data <= 32'h3845b8aa;
    11'b00000110000: data <= 32'h40d0bd1e;
    11'b00000110001: data <= 32'h40edb690;
    11'b00000110010: data <= 32'h3a2f3909;
    11'b00000110011: data <= 32'hb5d0394f;
    11'b00000110100: data <= 32'h332732dd;
    11'b00000110101: data <= 32'h3b762021;
    11'b00000110110: data <= 32'h28aeb73f;
    11'b00000110111: data <= 32'hbe20be89;
    11'b00000111000: data <= 32'hbe55c0de;
    11'b00000111001: data <= 32'ha218be12;
    11'b00000111010: data <= 32'h3c61358f;
    11'b00000111011: data <= 32'h383b3c36;
    11'b00000111100: data <= 32'hb920330e;
    11'b00000111101: data <= 32'hbc79b347;
    11'b00000111110: data <= 32'hbcaf3af2;
    11'b00000111111: data <= 32'hbdbc3fd7;
    11'b00001000000: data <= 32'hbd4b3c95;
    11'b00001000001: data <= 32'hadb2ba3b;
    11'b00001000010: data <= 32'h3d8ebd58;
    11'b00001000011: data <= 32'h3e252de0;
    11'b00001000100: data <= 32'h38833e45;
    11'b00001000101: data <= 32'h34733e21;
    11'b00001000110: data <= 32'h3cbe3958;
    11'b00001000111: data <= 32'h3e283223;
    11'b00001001000: data <= 32'h300daffc;
    11'b00001001001: data <= 32'hbe03bc02;
    11'b00001001010: data <= 32'hbc6abf6c;
    11'b00001001011: data <= 32'h3b46be45;
    11'b00001001100: data <= 32'h3fd3b837;
    11'b00001001101: data <= 32'h3b20b26b;
    11'b00001001110: data <= 32'hb9adb997;
    11'b00001001111: data <= 32'hbcbbb802;
    11'b00001010000: data <= 32'hbbc43b1c;
    11'b00001010001: data <= 32'hbcdb3ec9;
    11'b00001010010: data <= 32'hbe6d3723;
    11'b00001010011: data <= 32'hbc6cbdec;
    11'b00001010100: data <= 32'h21adbe14;
    11'b00001010101: data <= 32'h37f13768;
    11'b00001010110: data <= 32'h343a4019;
    11'b00001010111: data <= 32'h37923ef5;
    11'b00001011000: data <= 32'h3d1b39c8;
    11'b00001011001: data <= 32'h3ce038a9;
    11'b00001011010: data <= 32'hb4d83b14;
    11'b00001011011: data <= 32'hbdfb352c;
    11'b00001011100: data <= 32'hb7dfbb20;
    11'b00001011101: data <= 32'h3ee8bda4;
    11'b00001011110: data <= 32'h40f6bbff;
    11'b00001011111: data <= 32'h3c5eb9a0;
    11'b00001100000: data <= 32'hb62dba7d;
    11'b00001100001: data <= 32'hb5e9b610;
    11'b00001100010: data <= 32'h304e39d7;
    11'b00001100011: data <= 32'hb76e3bdc;
    11'b00001100100: data <= 32'hbeccb839;
    11'b00001100101: data <= 32'hbfa1c056;
    11'b00001100110: data <= 32'hbb17beef;
    11'b00001100111: data <= 32'h221535c6;
    11'b00001101000: data <= 32'h30d83e6a;
    11'b00001101001: data <= 32'h343c3bef;
    11'b00001101010: data <= 32'h3903340a;
    11'b00001101011: data <= 32'h34db3b6c;
    11'b00001101100: data <= 32'hbbb33fe9;
    11'b00001101101: data <= 32'hbe653e21;
    11'b00001101110: data <= 32'hb4a7b143;
    11'b00001101111: data <= 32'h3ef1bcdd;
    11'b00001110000: data <= 32'h4054bb26;
    11'b00001110001: data <= 32'h3b34b468;
    11'b00001110010: data <= 32'h2f92b033;
    11'b00001110011: data <= 32'h3af72da7;
    11'b00001110100: data <= 32'h3e083912;
    11'b00001110101: data <= 32'h359a3792;
    11'b00001110110: data <= 32'hbe60bbae;
    11'b00001110111: data <= 32'hc024c082;
    11'b00001111000: data <= 32'hba86bf0d;
    11'b00001111001: data <= 32'h35adb130;
    11'b00001111010: data <= 32'h35a736bf;
    11'b00001111011: data <= 32'haaf0b585;
    11'b00001111100: data <= 32'hb036b802;
    11'b00001111101: data <= 32'hb6d73c1d;
    11'b00001111110: data <= 32'hbd42410b;
    11'b00001111111: data <= 32'hbee73f9f;
    11'b00010000000: data <= 32'hb981b09b;
    11'b00010000001: data <= 32'h3a76bcc1;
    11'b00010000010: data <= 32'h3c42b6e7;
    11'b00010000011: data <= 32'h356a38e4;
    11'b00010000100: data <= 32'h377f39dd;
    11'b00010000101: data <= 32'h3f32382d;
    11'b00010000110: data <= 32'h40a43993;
    11'b00010000111: data <= 32'h399138ed;
    11'b00010001000: data <= 32'hbdc8b699;
    11'b00010001001: data <= 32'hbe85be17;
    11'b00010001010: data <= 32'h25c0bde3;
    11'b00010001011: data <= 32'h3cbbb9e9;
    11'b00010001100: data <= 32'h39a3ba4e;
    11'b00010001101: data <= 32'hb258bdf0;
    11'b00010001110: data <= 32'hb56bbc46;
    11'b00010001111: data <= 32'hb4e23b23;
    11'b00010010000: data <= 32'hbbbf4094;
    11'b00010010001: data <= 32'hbec73d45;
    11'b00010010010: data <= 32'hbda4ba3d;
    11'b00010010011: data <= 32'hb829bd72;
    11'b00010010100: data <= 32'hb28fa56d;
    11'b00010010101: data <= 32'hb4a13cc7;
    11'b00010010110: data <= 32'h37843c0a;
    11'b00010010111: data <= 32'h3fa837af;
    11'b00010011000: data <= 32'h40483a81;
    11'b00010011001: data <= 32'h35ed3d63;
    11'b00010011010: data <= 32'hbda93ad8;
    11'b00010011011: data <= 32'hbc05b53c;
    11'b00010011100: data <= 32'h3b3bbbaf;
    11'b00010011101: data <= 32'h3f12bbdf;
    11'b00010011110: data <= 32'h3ab6bd3b;
    11'b00010011111: data <= 32'haebbbf12;
    11'b00010100000: data <= 32'h3312bc60;
    11'b00010100001: data <= 32'h39e73987;
    11'b00010100010: data <= 32'h19653e53;
    11'b00010100011: data <= 32'hbdb03505;
    11'b00010100100: data <= 32'hbfd6be10;
    11'b00010100101: data <= 32'hbdb4be23;
    11'b00010100110: data <= 32'hbb1e2bef;
    11'b00010100111: data <= 32'hb8cb3bcc;
    11'b00010101000: data <= 32'h32163542;
    11'b00010101001: data <= 32'h3d21b22a;
    11'b00010101010: data <= 32'h3cec3a61;
    11'b00010101011: data <= 32'hb51e4058;
    11'b00010101100: data <= 32'hbdfe4022;
    11'b00010101101: data <= 32'hb94938ff;
    11'b00010101110: data <= 32'h3c70b829;
    11'b00010101111: data <= 32'h3e17ba2d;
    11'b00010110000: data <= 32'h3788bb40;
    11'b00010110001: data <= 32'h2b19bc85;
    11'b00010110010: data <= 32'h3cc2b8fc;
    11'b00010110011: data <= 32'h403638b0;
    11'b00010110100: data <= 32'h3c3f3bbc;
    11'b00010110101: data <= 32'hbc1bb49a;
    11'b00010110110: data <= 32'hbfebbeb6;
    11'b00010110111: data <= 32'hbd8bbdaa;
    11'b00010111000: data <= 32'hb90ab098;
    11'b00010111001: data <= 32'hb6e62b91;
    11'b00010111010: data <= 32'hb063bbfe;
    11'b00010111011: data <= 32'h3741bcce;
    11'b00010111100: data <= 32'h35c13898;
    11'b00010111101: data <= 32'hba0a4114;
    11'b00010111110: data <= 32'hbe0d40f1;
    11'b00010111111: data <= 32'hba2f3a27;
    11'b00011000000: data <= 32'h3708b699;
    11'b00011000001: data <= 32'h3705b4a0;
    11'b00011000010: data <= 32'hb591265c;
    11'b00011000011: data <= 32'h2badb10c;
    11'b00011000100: data <= 32'h3fadaed1;
    11'b00011000101: data <= 32'h41e93893;
    11'b00011000110: data <= 32'h3e493ae5;
    11'b00011000111: data <= 32'hb9fa22c3;
    11'b00011001000: data <= 32'hbdfcbbcc;
    11'b00011001001: data <= 32'hb831bb07;
    11'b00011001010: data <= 32'h3455b5d3;
    11'b00011001011: data <= 32'h9e61bb79;
    11'b00011001100: data <= 32'hb544c05b;
    11'b00011001101: data <= 32'h28cebfe2;
    11'b00011001110: data <= 32'h33f33416;
    11'b00011001111: data <= 32'hb743407a;
    11'b00011010000: data <= 32'hbd063f81;
    11'b00011010001: data <= 32'hbc902e5b;
    11'b00011010010: data <= 32'hb946b91b;
    11'b00011010011: data <= 32'hbafb30d1;
    11'b00011010100: data <= 32'hbcd93a3d;
    11'b00011010101: data <= 32'hb16a3561;
    11'b00011010110: data <= 32'h3fc1ad5f;
    11'b00011010111: data <= 32'h419137e6;
    11'b00011011000: data <= 32'h3d043d01;
    11'b00011011001: data <= 32'hb9ea3c2d;
    11'b00011011010: data <= 32'hbacb3428;
    11'b00011011011: data <= 32'h37f7aec5;
    11'b00011011100: data <= 32'h3c36b55f;
    11'b00011011101: data <= 32'h32a6bd56;
    11'b00011011110: data <= 32'hb651c0f9;
    11'b00011011111: data <= 32'h3475c01b;
    11'b00011100000: data <= 32'h3c3428f2;
    11'b00011100001: data <= 32'h385f3e07;
    11'b00011100010: data <= 32'hb9ae3a13;
    11'b00011100011: data <= 32'hbd87ba7f;
    11'b00011100100: data <= 32'hbdb1bb34;
    11'b00011100101: data <= 32'hbe6935bb;
    11'b00011100110: data <= 32'hbe853acf;
    11'b00011100111: data <= 32'hb816aea8;
    11'b00011101000: data <= 32'h3d19ba29;
    11'b00011101001: data <= 32'h3f263299;
    11'b00011101010: data <= 32'h36a73efd;
    11'b00011101011: data <= 32'hbb51402f;
    11'b00011101100: data <= 32'hb68d3d17;
    11'b00011101101: data <= 32'h3bbe37e9;
    11'b00011101110: data <= 32'h3c31a120;
    11'b00011101111: data <= 32'hb0e8bb17;
    11'b00011110000: data <= 32'hb7ddbf2a;
    11'b00011110001: data <= 32'h3b48bddf;
    11'b00011110010: data <= 32'h407c249c;
    11'b00011110011: data <= 32'h3eb43a90;
    11'b00011110100: data <= 32'haef6ad29;
    11'b00011110101: data <= 32'hbcf2bcda;
    11'b00011110110: data <= 32'hbd48ba80;
    11'b00011110111: data <= 32'hbd413634;
    11'b00011111000: data <= 32'hbd923457;
    11'b00011111001: data <= 32'hba2ebcf8;
    11'b00011111010: data <= 32'h363abf69;
    11'b00011111011: data <= 32'h399fb41b;
    11'b00011111100: data <= 32'hb4183f9e;
    11'b00011111101: data <= 32'hbbdf40d6;
    11'b00011111110: data <= 32'hb5063dab;
    11'b00011111111: data <= 32'h390138b1;
    11'b00100000000: data <= 32'h313d3707;
    11'b00100000001: data <= 32'hbc2c2dd3;
    11'b00100000010: data <= 32'hb9ffb911;
    11'b00100000011: data <= 32'h3d90b9c9;
    11'b00100000100: data <= 32'h41fd2d27;
    11'b00100000101: data <= 32'h406e384d;
    11'b00100000110: data <= 32'h32c4ae4d;
    11'b00100000111: data <= 32'hb9f7b9c6;
    11'b00100001000: data <= 32'hb69cb2e0;
    11'b00100001001: data <= 32'hb420370e;
    11'b00100001010: data <= 32'hba13b726;
    11'b00100001011: data <= 32'hbafec0a1;
    11'b00100001100: data <= 32'hb193c15b;
    11'b00100001101: data <= 32'h3491b960;
    11'b00100001110: data <= 32'hb1d33e33;
    11'b00100001111: data <= 32'hb9813f18;
    11'b00100010000: data <= 32'hb68938fe;
    11'b00100010001: data <= 32'hb1b331d1;
    11'b00100010010: data <= 32'hbc1e3a4b;
    11'b00100010011: data <= 32'hbff23bbe;
    11'b00100010100: data <= 32'hbc8230d4;
    11'b00100010101: data <= 32'h3d40b759;
    11'b00100010110: data <= 32'h418aa055;
    11'b00100010111: data <= 32'h3f3c3952;
    11'b00100011000: data <= 32'h2d2738fe;
    11'b00100011001: data <= 32'hb1bb3619;
    11'b00100011010: data <= 32'h39b2393c;
    11'b00100011011: data <= 32'h3a5f394f;
    11'b00100011100: data <= 32'hb4b6b9a6;
    11'b00100011101: data <= 32'hbb5dc122;
    11'b00100011110: data <= 32'hb1a0c16b;
    11'b00100011111: data <= 32'h3a2bba62;
    11'b00100100000: data <= 32'h39593b02;
    11'b00100100001: data <= 32'ha92e3886;
    11'b00100100010: data <= 32'hb6b5b84f;
    11'b00100100011: data <= 32'hba1cb553;
    11'b00100100100: data <= 32'hbece3b97;
    11'b00100100101: data <= 32'hc0ca3d08;
    11'b00100100110: data <= 32'hbdbb27ba;
    11'b00100100111: data <= 32'h396ebbcb;
    11'b00100101000: data <= 32'h3ec3b63b;
    11'b00100101001: data <= 32'h39ef3b41;
    11'b00100101010: data <= 32'hb5713dd8;
    11'b00100101011: data <= 32'h324d3d53;
    11'b00100101100: data <= 32'h3d843d26;
    11'b00100101101: data <= 32'h3c713c0c;
    11'b00100101110: data <= 32'hb764b419;
    11'b00100101111: data <= 32'hbc5ebf31;
    11'b00100110000: data <= 32'h322bbfb5;
    11'b00100110001: data <= 32'h3ee6b8b8;
    11'b00100110010: data <= 32'h3eea3435;
    11'b00100110011: data <= 32'h3907b740;
    11'b00100110100: data <= 32'hb229bd09;
    11'b00100110101: data <= 32'hb8f8b761;
    11'b00100110110: data <= 32'hbd653c1e;
    11'b00100110111: data <= 32'hc0003b87;
    11'b00100111000: data <= 32'hbdfbbacc;
    11'b00100111001: data <= 32'hb037bfe8;
    11'b00100111010: data <= 32'h3719bb8f;
    11'b00100111011: data <= 32'hb3e63b72;
    11'b00100111100: data <= 32'hb92d3ed6;
    11'b00100111101: data <= 32'h35143db1;
    11'b00100111110: data <= 32'h3d2d3d12;
    11'b00100111111: data <= 32'h38063d37;
    11'b00101000000: data <= 32'hbd05393d;
    11'b00101000001: data <= 32'hbdd4b7e4;
    11'b00101000010: data <= 32'h37fdbafc;
    11'b00101000011: data <= 32'h40bbb45c;
    11'b00101000100: data <= 32'h4071a4b4;
    11'b00101000101: data <= 32'h3b17b9c2;
    11'b00101000110: data <= 32'h3234bc3f;
    11'b00101000111: data <= 32'h339a24f0;
    11'b00101001000: data <= 32'hb1383cc5;
    11'b00101001001: data <= 32'hbc4d36d7;
    11'b00101001010: data <= 32'hbd56bf1f;
    11'b00101001011: data <= 32'hb95dc187;
    11'b00101001100: data <= 32'hb2cebd62;
    11'b00101001101: data <= 32'hb7c33900;
    11'b00101001110: data <= 32'hb7f23c5b;
    11'b00101001111: data <= 32'h35363821;
    11'b00101010000: data <= 32'h39bb38cc;
    11'b00101010001: data <= 32'hb8323d96;
    11'b00101010010: data <= 32'hc0543df6;
    11'b00101010011: data <= 32'hbf733826;
    11'b00101010100: data <= 32'h36a3b47e;
    11'b00101010101: data <= 32'h4047b1e3;
    11'b00101010110: data <= 32'h3ee125b8;
    11'b00101010111: data <= 32'h383db3a8;
    11'b00101011000: data <= 32'h3835b0d7;
    11'b00101011001: data <= 32'h3d413ad2;
    11'b00101011010: data <= 32'h3c6d3deb;
    11'b00101011011: data <= 32'hb45a3329;
    11'b00101011100: data <= 32'hbcafc003;
    11'b00101011101: data <= 32'hb9e3c16f;
    11'b00101011110: data <= 32'h258fbd29;
    11'b00101011111: data <= 32'h309f30e9;
    11'b00101100000: data <= 32'h2eb4aca8;
    11'b00101100001: data <= 32'h3684bacc;
    11'b00101100010: data <= 32'h336cb418;
    11'b00101100011: data <= 32'hbc973d4c;
    11'b00101100100: data <= 32'hc10a3f48;
    11'b00101100101: data <= 32'hc012393a;
    11'b00101100110: data <= 32'hab45b85c;
    11'b00101100111: data <= 32'h3c64b7f3;
    11'b00101101000: data <= 32'h376b310a;
    11'b00101101001: data <= 32'hb3373753;
    11'b00101101010: data <= 32'h393939d2;
    11'b00101101011: data <= 32'h40003dcf;
    11'b00101101100: data <= 32'h3eb63f00;
    11'b00101101101: data <= 32'hb1183875;
    11'b00101101110: data <= 32'hbcfbbd11;
    11'b00101101111: data <= 32'hb79bbf0e;
    11'b00101110000: data <= 32'h3a6cba1c;
    11'b00101110001: data <= 32'h3c6eb29a;
    11'b00101110010: data <= 32'h3a0dbc63;
    11'b00101110011: data <= 32'h38ddbf51;
    11'b00101110100: data <= 32'h34e8b989;
    11'b00101110101: data <= 32'hba833d18;
    11'b00101110110: data <= 32'hbfea3e69;
    11'b00101110111: data <= 32'hbf3da7a9;
    11'b00101111000: data <= 32'hb8f7bdb0;
    11'b00101111001: data <= 32'hb0a5bc2a;
    11'b00101111010: data <= 32'hba483133;
    11'b00101111011: data <= 32'hbaea39cd;
    11'b00101111100: data <= 32'h38e13a9d;
    11'b00101111101: data <= 32'h40013d46;
    11'b00101111110: data <= 32'h3d253f2d;
    11'b00101111111: data <= 32'hba613cf6;
    11'b00110000000: data <= 32'hbe602723;
    11'b00110000001: data <= 32'hb314b741;
    11'b00110000010: data <= 32'h3dadae23;
    11'b00110000011: data <= 32'h3e61b4b6;
    11'b00110000100: data <= 32'h3b75bdc1;
    11'b00110000101: data <= 32'h3a5fbf78;
    11'b00110000110: data <= 32'h3bb9b667;
    11'b00110000111: data <= 32'h35be3da0;
    11'b00110001000: data <= 32'hba753ca8;
    11'b00110001001: data <= 32'hbd29bb2e;
    11'b00110001010: data <= 32'hbb88c060;
    11'b00110001011: data <= 32'hbaebbd8e;
    11'b00110001100: data <= 32'hbd1d14f6;
    11'b00110001101: data <= 32'hbb863449;
    11'b00110001110: data <= 32'h3887ac3f;
    11'b00110001111: data <= 32'h3e0e36cb;
    11'b00110010000: data <= 32'h35b33e22;
    11'b00110010001: data <= 32'hbeae3f5f;
    11'b00110010010: data <= 32'hbfe33c5e;
    11'b00110010011: data <= 32'hb2c93698;
    11'b00110010100: data <= 32'h3d453428;
    11'b00110010101: data <= 32'h3c6cb184;
    11'b00110010110: data <= 32'h3606bc37;
    11'b00110010111: data <= 32'h3a60bc58;
    11'b00110011000: data <= 32'h3f393604;
    11'b00110011001: data <= 32'h3eaf3ebc;
    11'b00110011010: data <= 32'h34833b4d;
    11'b00110011011: data <= 32'hba91bcd8;
    11'b00110011100: data <= 32'hbb22c050;
    11'b00110011101: data <= 32'hb9d3bcaa;
    11'b00110011110: data <= 32'hba7fb17b;
    11'b00110011111: data <= 32'hb6ccb956;
    11'b00110100000: data <= 32'h3929bddf;
    11'b00110100001: data <= 32'h3c16b9c7;
    11'b00110100010: data <= 32'hb51b3c80;
    11'b00110100011: data <= 32'hc014400c;
    11'b00110100100: data <= 32'hc0073d49;
    11'b00110100101: data <= 32'hb6cd3584;
    11'b00110100110: data <= 32'h37c42c81;
    11'b00110100111: data <= 32'hb1c4a7e5;
    11'b00110101000: data <= 32'hb956b61a;
    11'b00110101001: data <= 32'h3890b20c;
    11'b00110101010: data <= 32'h40a33bef;
    11'b00110101011: data <= 32'h40ab3f72;
    11'b00110101100: data <= 32'h38fd3c21;
    11'b00110101101: data <= 32'hb9d2b948;
    11'b00110101110: data <= 32'hb8dfbcb7;
    11'b00110101111: data <= 32'h1bd2b5cf;
    11'b00110110000: data <= 32'h3044b183;
    11'b00110110001: data <= 32'h3396be00;
    11'b00110110010: data <= 32'h3a50c112;
    11'b00110110011: data <= 32'h3b71bdaa;
    11'b00110110100: data <= 32'hb0e13ae7;
    11'b00110110101: data <= 32'hbdf23f0a;
    11'b00110110110: data <= 32'hbe2039a2;
    11'b00110110111: data <= 32'hb918b7a2;
    11'b00110111000: data <= 32'hb877b780;
    11'b00110111001: data <= 32'hbe121afa;
    11'b00110111010: data <= 32'hbe5d1cd1;
    11'b00110111011: data <= 32'h34582aa6;
    11'b00110111100: data <= 32'h407e3ae0;
    11'b00110111101: data <= 32'h400a3eba;
    11'b00110111110: data <= 32'h2d073d86;
    11'b00110111111: data <= 32'hbc2f36eb;
    11'b00111000000: data <= 32'hb57532fb;
    11'b00111000001: data <= 32'h399438e2;
    11'b00111000010: data <= 32'h39e3284a;
    11'b00111000011: data <= 32'h36ddbef9;
    11'b00111000100: data <= 32'h3a5ac154;
    11'b00111000101: data <= 32'h3d23bd08;
    11'b00111000110: data <= 32'h3a913b76;
    11'b00111000111: data <= 32'hb3873d3f;
    11'b00111001000: data <= 32'hb98fb296;
    11'b00111001001: data <= 32'hb910bd52;
    11'b00111001010: data <= 32'hbca0babe;
    11'b00111001011: data <= 32'hc03aa437;
    11'b00111001100: data <= 32'hbf5fb1f0;
    11'b00111001101: data <= 32'h3000b930;
    11'b00111001110: data <= 32'h3ef9ae7f;
    11'b00111001111: data <= 32'h3c4e3c6d;
    11'b00111010000: data <= 32'hbad13e8f;
    11'b00111010001: data <= 32'hbdd13d6c;
    11'b00111010010: data <= 32'hb34e3ccb;
    11'b00111010011: data <= 32'h3a933cc0;
    11'b00111010100: data <= 32'h36dc34db;
    11'b00111010101: data <= 32'hb1a4bd54;
    11'b00111010110: data <= 32'h37f4bf94;
    11'b00111010111: data <= 32'h3f1ab74d;
    11'b00111011000: data <= 32'h3fe93cf1;
    11'b00111011001: data <= 32'h3bd03be6;
    11'b00111011010: data <= 32'h28bab9ab;
    11'b00111011011: data <= 32'hb632bddf;
    11'b00111011100: data <= 32'hbbd2b8ba;
    11'b00111011101: data <= 32'hbebe2d31;
    11'b00111011110: data <= 32'hbd5dba3c;
    11'b00111011111: data <= 32'h32f6bf8c;
    11'b00111100000: data <= 32'h3ccebd7e;
    11'b00111100001: data <= 32'h33e63672;
    11'b00111100010: data <= 32'hbd853e52;
    11'b00111100011: data <= 32'hbdf53e1a;
    11'b00111100100: data <= 32'hb28f3cc9;
    11'b00111100101: data <= 32'h35043c3c;
    11'b00111100110: data <= 32'hb986374d;
    11'b00111100111: data <= 32'hbd5fb902;
    11'b00111101000: data <= 32'ha9edbb05;
    11'b00111101001: data <= 32'h400534dc;
    11'b00111101010: data <= 32'h41203db5;
    11'b00111101011: data <= 32'h3da23b43;
    11'b00111101100: data <= 32'h33c7b755;
    11'b00111101101: data <= 32'hab49b948;
    11'b00111101110: data <= 32'hb3073539;
    11'b00111101111: data <= 32'hb93a367b;
    11'b00111110000: data <= 32'hb86fbd3d;
    11'b00111110001: data <= 32'h3646c1ba;
    11'b00111110010: data <= 32'h3b96c05c;
    11'b00111110011: data <= 32'h3061a692;
    11'b00111110100: data <= 32'hbbff3ce6;
    11'b00111110101: data <= 32'hbb443b0b;
    11'b00111110110: data <= 32'hae153524;
    11'b00111110111: data <= 32'hb69c36c3;
    11'b00111111000: data <= 32'hbfb4373b;
    11'b00111111001: data <= 32'hc0ccaf47;
    11'b00111111010: data <= 32'hb87ab62f;
    11'b00111111011: data <= 32'h3f363599;
    11'b00111111100: data <= 32'h406e3cb2;
    11'b00111111101: data <= 32'h3ac13b99;
    11'b00111111110: data <= 32'hb04a34fc;
    11'b00111111111: data <= 32'h31ab3904;
    11'b01000000000: data <= 32'h38923dcc;
    11'b01000000001: data <= 32'h31773af3;
    11'b01000000010: data <= 32'hb1cbbd80;
    11'b01000000011: data <= 32'h35a8c1e6;
    11'b01000000100: data <= 32'h3c15c013;
    11'b01000000101: data <= 32'h3a4e2b58;
    11'b01000000110: data <= 32'h303d3a57;
    11'b01000000111: data <= 32'h2d85aed2;
    11'b01000001000: data <= 32'h326eb9cb;
    11'b01000001001: data <= 32'hba60b027;
    11'b01000001010: data <= 32'hc0f43724;
    11'b01000001011: data <= 32'hc168ab05;
    11'b01000001100: data <= 32'hb9f4ba2e;
    11'b01000001101: data <= 32'h3d27b7a9;
    11'b01000001110: data <= 32'h3cd3371b;
    11'b01000001111: data <= 32'hb3f33b24;
    11'b01000010000: data <= 32'hb9ae3beb;
    11'b01000010001: data <= 32'h34803e3c;
    11'b01000010010: data <= 32'h3b4a403c;
    11'b01000010011: data <= 32'h314d3ced;
    11'b01000010100: data <= 32'hb91dbb5e;
    11'b01000010101: data <= 32'had4ac040;
    11'b01000010110: data <= 32'h3cc1bc6c;
    11'b01000010111: data <= 32'h3eb53816;
    11'b01000011000: data <= 32'h3d2a37dc;
    11'b01000011001: data <= 32'h3b8eba5a;
    11'b01000011010: data <= 32'h38c7bc99;
    11'b01000011011: data <= 32'hb850a909;
    11'b01000011100: data <= 32'hc0013945;
    11'b01000011101: data <= 32'hc037b549;
    11'b01000011110: data <= 32'hb83abee7;
    11'b01000011111: data <= 32'h3a32bec3;
    11'b01000100000: data <= 32'h32f7b69d;
    11'b01000100001: data <= 32'hbc323909;
    11'b01000100010: data <= 32'hbb5d3c2c;
    11'b01000100011: data <= 32'h36443e13;
    11'b01000100100: data <= 32'h39a63fc1;
    11'b01000100101: data <= 32'hb9493d34;
    11'b01000100110: data <= 32'hbef0b3a2;
    11'b01000100111: data <= 32'hba5ebbc3;
    11'b01000101000: data <= 32'h3cb4adac;
    11'b01000101001: data <= 32'h40373b1b;
    11'b01000101010: data <= 32'h3ec535a8;
    11'b01000101011: data <= 32'h3c99baa1;
    11'b01000101100: data <= 32'h3b25b91d;
    11'b01000101101: data <= 32'h32b43a5a;
    11'b01000101110: data <= 32'hbad33ca1;
    11'b01000101111: data <= 32'hbc58b8aa;
    11'b01000110000: data <= 32'hb134c10a;
    11'b01000110001: data <= 32'h37d8c0f2;
    11'b01000110010: data <= 32'hb100bb1d;
    11'b01000110011: data <= 32'hbbc43408;
    11'b01000110100: data <= 32'hb7113625;
    11'b01000110101: data <= 32'h395d385e;
    11'b01000110110: data <= 32'h34683c64;
    11'b01000110111: data <= 32'hbec23c70;
    11'b01000111000: data <= 32'hc18b3485;
    11'b01000111001: data <= 32'hbd9ab397;
    11'b01000111010: data <= 32'h3b1d3435;
    11'b01000111011: data <= 32'h3ee03a16;
    11'b01000111100: data <= 32'h3c3133b8;
    11'b01000111101: data <= 32'h38d8b5d2;
    11'b01000111110: data <= 32'h3bae36c4;
    11'b01000111111: data <= 32'h3bf63f98;
    11'b01001000000: data <= 32'h321e3f00;
    11'b01001000001: data <= 32'hb682b820;
    11'b01001000010: data <= 32'haa5cc112;
    11'b01001000011: data <= 32'h36ecc089;
    11'b01001000100: data <= 32'h3205b97a;
    11'b01001000101: data <= 32'had45a9e2;
    11'b01001000110: data <= 32'h383fb8c2;
    11'b01001000111: data <= 32'h3c80b995;
    11'b01001001000: data <= 32'h2c8333ce;
    11'b01001001001: data <= 32'hc04a3b70;
    11'b01001001010: data <= 32'hc2113718;
    11'b01001001011: data <= 32'hbe0eb522;
    11'b01001001100: data <= 32'h3779b4d9;
    11'b01001001101: data <= 32'h39b22c30;
    11'b01001001110: data <= 32'hb3231f8b;
    11'b01001001111: data <= 32'hb4232e2e;
    11'b01001010000: data <= 32'h3b003cf2;
    11'b01001010001: data <= 32'h3da34116;
    11'b01001010010: data <= 32'h37a84031;
    11'b01001010011: data <= 32'hb8acaece;
    11'b01001010100: data <= 32'hb6dfbece;
    11'b01001010101: data <= 32'h36b1bcb5;
    11'b01001010110: data <= 32'h3a9f289a;
    11'b01001010111: data <= 32'h3b7fb0f3;
    11'b01001011000: data <= 32'h3d8bbd57;
    11'b01001011001: data <= 32'h3e3bbd9e;
    11'b01001011010: data <= 32'h355928c6;
    11'b01001011011: data <= 32'hbe963c3b;
    11'b01001011100: data <= 32'hc09b3578;
    11'b01001011101: data <= 32'hbc3fbc04;
    11'b01001011110: data <= 32'h3069bd69;
    11'b01001011111: data <= 32'hb50bba67;
    11'b01001100000: data <= 32'hbd2db578;
    11'b01001100001: data <= 32'hba3b2de0;
    11'b01001100010: data <= 32'h3af93ca3;
    11'b01001100011: data <= 32'h3d734085;
    11'b01001100100: data <= 32'hac2a3fdf;
    11'b01001100101: data <= 32'hbdfa368d;
    11'b01001100110: data <= 32'hbc9cb821;
    11'b01001100111: data <= 32'h34792e5f;
    11'b01001101000: data <= 32'h3c9d39dc;
    11'b01001101001: data <= 32'h3d25b0dd;
    11'b01001101010: data <= 32'h3e12be08;
    11'b01001101011: data <= 32'h3ed6bcbd;
    11'b01001101100: data <= 32'h3b913949;
    11'b01001101101: data <= 32'hb78e3e3c;
    11'b01001101110: data <= 32'hbc2433b9;
    11'b01001101111: data <= 32'hb5f7be99;
    11'b01001110000: data <= 32'h244dc022;
    11'b01001110001: data <= 32'hba79bcf1;
    11'b01001110010: data <= 32'hbe0cb90f;
    11'b01001110011: data <= 32'hb849b780;
    11'b01001110100: data <= 32'h3c8c3132;
    11'b01001110101: data <= 32'h3c643cc9;
    11'b01001110110: data <= 32'hbb4c3dda;
    11'b01001110111: data <= 32'hc0e43a04;
    11'b01001111000: data <= 32'hbefb351d;
    11'b01001111001: data <= 32'h25ba3a09;
    11'b01001111010: data <= 32'h3a8a3af3;
    11'b01001111011: data <= 32'h38ecb341;
    11'b01001111100: data <= 32'h3a3fbcdc;
    11'b01001111101: data <= 32'h3df0b54d;
    11'b01001111110: data <= 32'h3e323ea9;
    11'b01001111111: data <= 32'h39464052;
    11'b01010000000: data <= 32'haa4f354d;
    11'b01010000001: data <= 32'h2836beb2;
    11'b01010000010: data <= 32'h2695bf53;
    11'b01010000011: data <= 32'hb914baf9;
    11'b01010000100: data <= 32'hbaddb965;
    11'b01010000101: data <= 32'h3511bd18;
    11'b01010000110: data <= 32'h3e74bca0;
    11'b01010000111: data <= 32'h3bad28cf;
    11'b01010001000: data <= 32'hbd573bba;
    11'b01010001001: data <= 32'hc1593a85;
    11'b01010001010: data <= 32'hbef13663;
    11'b01010001011: data <= 32'hb2113723;
    11'b01010001100: data <= 32'ha89c3521;
    11'b01010001101: data <= 32'hb9c9b7ca;
    11'b01010001110: data <= 32'hb613badd;
    11'b01010001111: data <= 32'h3c45369e;
    11'b01010010000: data <= 32'h3f58408d;
    11'b01010010001: data <= 32'h3c6640d8;
    11'b01010010010: data <= 32'h2adf38a7;
    11'b01010010011: data <= 32'hb151bbbc;
    11'b01010010100: data <= 32'h9eadb96f;
    11'b01010010101: data <= 32'hb00a3021;
    11'b01010010110: data <= 32'h2b64b736;
    11'b01010010111: data <= 32'h3c89bf79;
    11'b01010011000: data <= 32'h4001c002;
    11'b01010011001: data <= 32'h3c78b780;
    11'b01010011010: data <= 32'hbb7a3b01;
    11'b01010011011: data <= 32'hbf9039b1;
    11'b01010011100: data <= 32'hbc1bb056;
    11'b01010011101: data <= 32'hb24eb771;
    11'b01010011110: data <= 32'hbb44b7fc;
    11'b01010011111: data <= 32'hbfb6ba9d;
    11'b01010100000: data <= 32'hbcdcba7c;
    11'b01010100001: data <= 32'h3a7a3671;
    11'b01010100010: data <= 32'h3f0b3fcb;
    11'b01010100011: data <= 32'h39b54024;
    11'b01010100100: data <= 32'hb97b3a62;
    11'b01010100101: data <= 32'hba9b2c10;
    11'b01010100110: data <= 32'hb11d39cc;
    11'b01010100111: data <= 32'h32723c9d;
    11'b01010101000: data <= 32'h370fb12a;
    11'b01010101001: data <= 32'h3cf0bff1;
    11'b01010101010: data <= 32'h3fe2bfca;
    11'b01010101011: data <= 32'h3ddbaa37;
    11'b01010101100: data <= 32'h2de73d25;
    11'b01010101101: data <= 32'hb8053918;
    11'b01010101110: data <= 32'h9c84b9ed;
    11'b01010101111: data <= 32'h9e76bcba;
    11'b01010110000: data <= 32'hbd4bbb4f;
    11'b01010110001: data <= 32'hc09fbbd9;
    11'b01010110010: data <= 32'hbcd5bc99;
    11'b01010110011: data <= 32'h3b9eb755;
    11'b01010110100: data <= 32'h3e163a32;
    11'b01010110101: data <= 32'habd83cf2;
    11'b01010110110: data <= 32'hbe6e3a81;
    11'b01010110111: data <= 32'hbd9c3a68;
    11'b01010111000: data <= 32'hb53a3e33;
    11'b01010111001: data <= 32'h28df3e3c;
    11'b01010111010: data <= 32'haf0cace4;
    11'b01010111011: data <= 32'h3675bed6;
    11'b01010111100: data <= 32'h3dbdbcc4;
    11'b01010111101: data <= 32'h3ef13b29;
    11'b01010111110: data <= 32'h3c713f7d;
    11'b01010111111: data <= 32'h39423967;
    11'b01011000000: data <= 32'h39a0bb1d;
    11'b01011000001: data <= 32'h327ebc2e;
    11'b01011000010: data <= 32'hbc9ab797;
    11'b01011000011: data <= 32'hbf1bb9f2;
    11'b01011000100: data <= 32'hb731be89;
    11'b01011000101: data <= 32'h3da0bea0;
    11'b01011000110: data <= 32'h3d73b875;
    11'b01011000111: data <= 32'hb881368c;
    11'b01011001000: data <= 32'hbfa93913;
    11'b01011001001: data <= 32'hbd5a3aea;
    11'b01011001010: data <= 32'hb4c43d86;
    11'b01011001011: data <= 32'hb8283c91;
    11'b01011001100: data <= 32'hbd4db4c0;
    11'b01011001101: data <= 32'hbb66bd69;
    11'b01011001110: data <= 32'h395fb684;
    11'b01011001111: data <= 32'h3efd3e43;
    11'b01011010000: data <= 32'h3e0f4033;
    11'b01011010001: data <= 32'h3b5c39d3;
    11'b01011010010: data <= 32'h3970b71d;
    11'b01011010011: data <= 32'h339ca217;
    11'b01011010100: data <= 32'hb93f397b;
    11'b01011010101: data <= 32'hbaddb15d;
    11'b01011010110: data <= 32'h3684bfb6;
    11'b01011010111: data <= 32'h3f1dc0e6;
    11'b01011011000: data <= 32'h3d79bcf5;
    11'b01011011001: data <= 32'hb63c2e43;
    11'b01011011010: data <= 32'hbcfa36d3;
    11'b01011011011: data <= 32'hb7c2358a;
    11'b01011011100: data <= 32'h28f23803;
    11'b01011011101: data <= 32'hbc5334f2;
    11'b01011011110: data <= 32'hc0edb913;
    11'b01011011111: data <= 32'hbfcdbcc8;
    11'b01011100000: data <= 32'h30c1b349;
    11'b01011100001: data <= 32'h3e193d63;
    11'b01011100010: data <= 32'h3c8f3e80;
    11'b01011100011: data <= 32'h33da38f5;
    11'b01011100100: data <= 32'h29303465;
    11'b01011100101: data <= 32'h2d603d46;
    11'b01011100110: data <= 32'hb41e3fa4;
    11'b01011100111: data <= 32'hb52336c9;
    11'b01011101000: data <= 32'h38e9bf6f;
    11'b01011101001: data <= 32'h3e9cc0ca;
    11'b01011101010: data <= 32'h3dadbb50;
    11'b01011101011: data <= 32'h355c372a;
    11'b01011101100: data <= 32'h2c37357b;
    11'b01011101101: data <= 32'h39f5b4cd;
    11'b01011101110: data <= 32'h387eb549;
    11'b01011101111: data <= 32'hbd18b28f;
    11'b01011110000: data <= 32'hc1aeb9cd;
    11'b01011110001: data <= 32'hc022bd1d;
    11'b01011110010: data <= 32'h31e9ba6b;
    11'b01011110011: data <= 32'h3d04341c;
    11'b01011110100: data <= 32'h357e38af;
    11'b01011110101: data <= 32'hba0e3487;
    11'b01011110110: data <= 32'hb8ff3a18;
    11'b01011110111: data <= 32'haa1b4042;
    11'b01011111000: data <= 32'hb2a640f1;
    11'b01011111001: data <= 32'hb8de3950;
    11'b01011111010: data <= 32'hb008be15;
    11'b01011111011: data <= 32'h3b64be83;
    11'b01011111100: data <= 32'h3d542cc6;
    11'b01011111101: data <= 32'h3c543c6a;
    11'b01011111110: data <= 32'h3cd535dc;
    11'b01011111111: data <= 32'h3e8eb8f4;
    11'b01100000000: data <= 32'h3bd0b6e8;
    11'b01100000001: data <= 32'hbc07304d;
    11'b01100000010: data <= 32'hc09ab517;
    11'b01100000011: data <= 32'hbd32bda7;
    11'b01100000100: data <= 32'h3977bede;
    11'b01100000101: data <= 32'h3c5dbc34;
    11'b01100000110: data <= 32'hb4afb744;
    11'b01100000111: data <= 32'hbd19b0d1;
    11'b01100001000: data <= 32'hb955398f;
    11'b01100001001: data <= 32'h2fb23fdb;
    11'b01100001010: data <= 32'hb6fd402a;
    11'b01100001011: data <= 32'hbe2736ed;
    11'b01100001100: data <= 32'hbdb1bca5;
    11'b01100001101: data <= 32'hac65b9ea;
    11'b01100001110: data <= 32'h3c2f3b6f;
    11'b01100001111: data <= 32'h3d493dc5;
    11'b01100010000: data <= 32'h3de934fe;
    11'b01100010001: data <= 32'h3ebfb795;
    11'b01100010010: data <= 32'h3c2d3524;
    11'b01100010011: data <= 32'hb8003d04;
    11'b01100010100: data <= 32'hbd3837dd;
    11'b01100010101: data <= 32'hb48ebd84;
    11'b01100010110: data <= 32'h3caec0a1;
    11'b01100010111: data <= 32'h3c15befb;
    11'b01100011000: data <= 32'hb62cbb0e;
    11'b01100011001: data <= 32'hbb00b717;
    11'b01100011010: data <= 32'h305330b3;
    11'b01100011011: data <= 32'h39793c1c;
    11'b01100011100: data <= 32'hb93d3c7e;
    11'b01100011101: data <= 32'hc0eaa35b;
    11'b01100011110: data <= 32'hc0edbba7;
    11'b01100011111: data <= 32'hba00b535;
    11'b01100100000: data <= 32'h39783bc8;
    11'b01100100001: data <= 32'h3b1e3c23;
    11'b01100100010: data <= 32'h3a22a024;
    11'b01100100011: data <= 32'h3babae78;
    11'b01100100100: data <= 32'h3a5c3dac;
    11'b01100100101: data <= 32'hacbf40fd;
    11'b01100100110: data <= 32'hb8863d1c;
    11'b01100100111: data <= 32'h3190bc76;
    11'b01100101000: data <= 32'h3c83c058;
    11'b01100101001: data <= 32'h3b13bd99;
    11'b01100101010: data <= 32'h96f9b7ce;
    11'b01100101011: data <= 32'h321eb75e;
    11'b01100101100: data <= 32'h3d85b820;
    11'b01100101101: data <= 32'h3db82656;
    11'b01100101110: data <= 32'hb8dc35ed;
    11'b01100101111: data <= 32'hc170b2b7;
    11'b01100110000: data <= 32'hc127bb0f;
    11'b01100110001: data <= 32'hb9beb897;
    11'b01100110010: data <= 32'h370b304b;
    11'b01100110011: data <= 32'h2ce1a3e1;
    11'b01100110100: data <= 32'hb610b8b2;
    11'b01100110101: data <= 32'h2cb62efd;
    11'b01100110110: data <= 32'h385a402e;
    11'b01100110111: data <= 32'h2e404223;
    11'b01100111000: data <= 32'hb85f3e4a;
    11'b01100111001: data <= 32'hb4eaba11;
    11'b01100111010: data <= 32'h3677bd84;
    11'b01100111011: data <= 32'h3864b4af;
    11'b01100111100: data <= 32'h370e35cc;
    11'b01100111101: data <= 32'h3cb4b4ff;
    11'b01100111110: data <= 32'h409bbb68;
    11'b01100111111: data <= 32'h3fcdb5bf;
    11'b01101000000: data <= 32'hb4553720;
    11'b01101000001: data <= 32'hc047317a;
    11'b01101000010: data <= 32'hbedaba35;
    11'b01101000011: data <= 32'hab45bcaa;
    11'b01101000100: data <= 32'h3653bbfe;
    11'b01101000101: data <= 32'hb906bc66;
    11'b01101000110: data <= 32'hbc9fbcb3;
    11'b01101000111: data <= 32'hb387ad09;
    11'b01101001000: data <= 32'h39483f79;
    11'b01101001001: data <= 32'h2dce4139;
    11'b01101001010: data <= 32'hbc973cdf;
    11'b01101001011: data <= 32'hbda6b800;
    11'b01101001100: data <= 32'hb91eb6fd;
    11'b01101001101: data <= 32'h2c2e3a62;
    11'b01101001110: data <= 32'h38133bbd;
    11'b01101001111: data <= 32'h3d7eb4a2;
    11'b01101010000: data <= 32'h40a1bbd1;
    11'b01101010001: data <= 32'h3fc62c4a;
    11'b01101010010: data <= 32'h31333d6d;
    11'b01101010011: data <= 32'hbc623c1d;
    11'b01101010100: data <= 32'hb7c0b81f;
    11'b01101010101: data <= 32'h3987be33;
    11'b01101010110: data <= 32'h36c3be6b;
    11'b01101010111: data <= 32'hbb1fbe17;
    11'b01101011000: data <= 32'hbc4cbdcd;
    11'b01101011001: data <= 32'h357eb8b9;
    11'b01101011010: data <= 32'h3d0b3b1c;
    11'b01101011011: data <= 32'h2f5d3dda;
    11'b01101011100: data <= 32'hbf45382a;
    11'b01101011101: data <= 32'hc0b2b689;
    11'b01101011110: data <= 32'hbd612fbe;
    11'b01101011111: data <= 32'hb56a3c9c;
    11'b01101100000: data <= 32'h2c713a63;
    11'b01101100001: data <= 32'h38f0b905;
    11'b01101100010: data <= 32'h3db5bacb;
    11'b01101100011: data <= 32'h3ddf3b21;
    11'b01101100100: data <= 32'h377c40f5;
    11'b01101100101: data <= 32'hb3873f74;
    11'b01101100110: data <= 32'h3472b0f3;
    11'b01101100111: data <= 32'h3b3fbd67;
    11'b01101101000: data <= 32'h34aebcd6;
    11'b01101101001: data <= 32'hb9f6bc02;
    11'b01101101010: data <= 32'hb4c1bd1a;
    11'b01101101011: data <= 32'h3dd2bc8c;
    11'b01101101100: data <= 32'h4024b2f0;
    11'b01101101101: data <= 32'h34ea36ac;
    11'b01101101110: data <= 32'hbfe92ac8;
    11'b01101101111: data <= 32'hc0cfb5ea;
    11'b01101110000: data <= 32'hbce72e5f;
    11'b01101110001: data <= 32'hb6ff38ed;
    11'b01101110010: data <= 32'hb92dae80;
    11'b01101110011: data <= 32'hb8eebd1e;
    11'b01101110100: data <= 32'h343fba93;
    11'b01101110101: data <= 32'h3b7a3db1;
    11'b01101110110: data <= 32'h389a41fc;
    11'b01101110111: data <= 32'h9ef54038;
    11'b01101111000: data <= 32'h2efa2f2c;
    11'b01101111001: data <= 32'h35a8b900;
    11'b01101111010: data <= 32'haf42a606;
    11'b01101111011: data <= 32'hb81c2e8d;
    11'b01101111100: data <= 32'h3818bac5;
    11'b01101111101: data <= 32'h40a2bdd7;
    11'b01101111110: data <= 32'h412aba52;
    11'b01101111111: data <= 32'h38e1317f;
    11'b01110000000: data <= 32'hbdba3381;
    11'b01110000001: data <= 32'hbde0b29b;
    11'b01110000010: data <= 32'hb563b439;
    11'b01110000011: data <= 32'hb2e3b4fd;
    11'b01110000100: data <= 32'hbd01bc79;
    11'b01110000101: data <= 32'hbe40bf95;
    11'b01110000110: data <= 32'hb5e4bc21;
    11'b01110000111: data <= 32'h3a943ccc;
    11'b01110001000: data <= 32'h38cf40f1;
    11'b01110001001: data <= 32'hb5f43e3d;
    11'b01110001010: data <= 32'hba1c301f;
    11'b01110001011: data <= 32'hb8e732e2;
    11'b01110001100: data <= 32'hb93e3ce4;
    11'b01110001101: data <= 32'hb82d3c21;
    11'b01110001110: data <= 32'h3962b88f;
    11'b01110001111: data <= 32'h408abe10;
    11'b01110010000: data <= 32'h40d8b8c7;
    11'b01110010001: data <= 32'h3ab33a9c;
    11'b01110010010: data <= 32'hb7b63bfa;
    11'b01110010011: data <= 32'hae2a3035;
    11'b01110010100: data <= 32'h39ddb831;
    11'b01110010101: data <= 32'h2d74bac5;
    11'b01110010110: data <= 32'hbdf7bdfb;
    11'b01110010111: data <= 32'hbed7c021;
    11'b01110011000: data <= 32'hac57bd89;
    11'b01110011001: data <= 32'h3d3634ca;
    11'b01110011010: data <= 32'h39aa3cc0;
    11'b01110011011: data <= 32'hbb0f3867;
    11'b01110011100: data <= 32'hbe61ac1b;
    11'b01110011101: data <= 32'hbd1f39d4;
    11'b01110011110: data <= 32'hbc033f32;
    11'b01110011111: data <= 32'hbad73ca6;
    11'b01110100000: data <= 32'ha5c7ba14;
    11'b01110100001: data <= 32'h3d0fbddb;
    11'b01110100010: data <= 32'h3e9c2948;
    11'b01110100011: data <= 32'h3adb3f41;
    11'b01110100100: data <= 32'h35153f2f;
    11'b01110100101: data <= 32'h3b0c37b4;
    11'b01110100110: data <= 32'h3d11b5ff;
    11'b01110100111: data <= 32'h3057b7cd;
    11'b01110101000: data <= 32'hbda1bb03;
    11'b01110101001: data <= 32'hbc8abe84;
    11'b01110101010: data <= 32'h3b0dbea1;
    11'b01110101011: data <= 32'h4026b9e2;
    11'b01110101100: data <= 32'h3b69ac3e;
    11'b01110101101: data <= 32'hbc28b413;
    11'b01110101110: data <= 32'hbea6b3aa;
    11'b01110101111: data <= 32'hbc533a00;
    11'b01110110000: data <= 32'hbb113de8;
    11'b01110110001: data <= 32'hbd4c3741;
    11'b01110110010: data <= 32'hbcbbbd73;
    11'b01110110011: data <= 32'hae21bdf6;
    11'b01110110100: data <= 32'h3a2a3832;
    11'b01110110101: data <= 32'h39c1409f;
    11'b01110110110: data <= 32'h388b3fed;
    11'b01110110111: data <= 32'h3b8238a0;
    11'b01110111000: data <= 32'h3b803084;
    11'b01110111001: data <= 32'hb284390a;
    11'b01110111010: data <= 32'hbcfd36a2;
    11'b01110111011: data <= 32'hb69cbacd;
    11'b01110111100: data <= 32'h3ed2bed9;
    11'b01110111101: data <= 32'h4117bd3c;
    11'b01110111110: data <= 32'h3c70b85f;
    11'b01110111111: data <= 32'hb943b54d;
    11'b01111000000: data <= 32'hba47b177;
    11'b01111000001: data <= 32'ha5c1376f;
    11'b01111000010: data <= 32'hb52e395d;
    11'b01111000011: data <= 32'hbe99b805;
    11'b01111000100: data <= 32'hc039bfd2;
    11'b01111000101: data <= 32'hbbc2be84;
    11'b01111000110: data <= 32'h35d836b7;
    11'b01111000111: data <= 32'h38eb3f59;
    11'b01111001000: data <= 32'h34713d22;
    11'b01111001001: data <= 32'h32f23480;
    11'b01111001010: data <= 32'h2b9c39a6;
    11'b01111001011: data <= 32'hb9d93f65;
    11'b01111001100: data <= 32'hbceb3e5a;
    11'b01111001101: data <= 32'hb1abb403;
    11'b01111001110: data <= 32'h3ec8be65;
    11'b01111001111: data <= 32'h4085bcb8;
    11'b01111010000: data <= 32'h3c3aac6e;
    11'b01111010001: data <= 32'h27c534f3;
    11'b01111010010: data <= 32'h387230d7;
    11'b01111010011: data <= 32'h3d2932ef;
    11'b01111010100: data <= 32'h35292eb7;
    11'b01111010101: data <= 32'hbec0bb3e;
    11'b01111010110: data <= 32'hc09ec00f;
    11'b01111010111: data <= 32'hbaf3bef9;
    11'b01111011000: data <= 32'h397db3ba;
    11'b01111011001: data <= 32'h398838b5;
    11'b01111011010: data <= 32'hb234287d;
    11'b01111011011: data <= 32'hb8d5b458;
    11'b01111011100: data <= 32'hb8fa3bed;
    11'b01111011101: data <= 32'hbc1240ec;
    11'b01111011110: data <= 32'hbd7f3fc0;
    11'b01111011111: data <= 32'hb94fb3aa;
    11'b01111100000: data <= 32'h39cfbdf9;
    11'b01111100001: data <= 32'h3d10b8c4;
    11'b01111100010: data <= 32'h39b53af7;
    11'b01111100011: data <= 32'h38ab3c6b;
    11'b01111100100: data <= 32'h3e403779;
    11'b01111100101: data <= 32'h40213358;
    11'b01111100110: data <= 32'h38ec34a0;
    11'b01111100111: data <= 32'hbe14b538;
    11'b01111101000: data <= 32'hbf2dbd90;
    11'b01111101001: data <= 32'h91e5bea9;
    11'b01111101010: data <= 32'h3dbabc15;
    11'b01111101011: data <= 32'h3b26b981;
    11'b01111101100: data <= 32'hb709bc1f;
    11'b01111101101: data <= 32'hba78b9d7;
    11'b01111101110: data <= 32'hb76f3b2b;
    11'b01111101111: data <= 32'hb9cd4068;
    11'b01111110000: data <= 32'hbe113d5f;
    11'b01111110001: data <= 32'hbe46ba4f;
    11'b01111110010: data <= 32'hb934be0a;
    11'b01111110011: data <= 32'h2ef7ac03;
    11'b01111110100: data <= 32'h34133de2;
    11'b01111110101: data <= 32'h39793d55;
    11'b01111110110: data <= 32'h3ebd36d3;
    11'b01111110111: data <= 32'h3f8a374b;
    11'b01111111000: data <= 32'h35d73ca6;
    11'b01111111001: data <= 32'hbd633bc8;
    11'b01111111010: data <= 32'hbc37b55a;
    11'b01111111011: data <= 32'h3b20bd7b;
    11'b01111111100: data <= 32'h3fc7bda8;
    11'b01111111101: data <= 32'h3bcbbcef;
    11'b01111111110: data <= 32'hb4e2bd2c;
    11'b01111111111: data <= 32'hb102ba5a;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    