module adder_tree(
CLK, rst, 
input_a_real1_vmm0, input_a_real2_vmm0,  input_a_real3_vmm0,  input_a_real4_vmm0,  input_a_real5_vmm0,  input_a_real6_vmm0,  input_a_real7_vmm0,  input_a_real8_vmm0,
input_a_imag1_vmm0, input_a_imag2_vmm0,  input_a_imag3_vmm0,  input_a_imag4_vmm0,  input_a_imag5_vmm0,  input_a_imag6_vmm0,  input_a_imag7_vmm0,  input_a_imag8_vmm0,
input_a_real9_vmm0, input_a_real10_vmm0, input_a_real11_vmm0, input_a_real12_vmm0, input_a_real13_vmm0, input_a_real14_vmm0, input_a_real15_vmm0, input_a_real16_vmm0,
input_a_imag9_vmm0, input_a_imag10_vmm0, input_a_imag11_vmm0, input_a_imag12_vmm0, input_a_imag13_vmm0, input_a_imag14_vmm0, input_a_imag15_vmm0, input_a_imag16_vmm0,
input_a_real1_vmm1, input_a_real2_vmm1,  input_a_real3_vmm1,  input_a_real4_vmm1,  input_a_real5_vmm1,  input_a_real6_vmm1,  input_a_real7_vmm1,  input_a_real8_vmm1,
input_a_imag1_vmm1, input_a_imag2_vmm1,  input_a_imag3_vmm1,  input_a_imag4_vmm1,  input_a_imag5_vmm1,  input_a_imag6_vmm1,  input_a_imag7_vmm1,  input_a_imag8_vmm1,
input_a_real9_vmm1, input_a_real10_vmm1, input_a_real11_vmm1, input_a_real12_vmm1, input_a_real13_vmm1, input_a_real14_vmm1, input_a_real15_vmm1, input_a_real16_vmm1,
input_a_imag9_vmm1, input_a_imag10_vmm1, input_a_imag11_vmm1, input_a_imag12_vmm1, input_a_imag13_vmm1, input_a_imag14_vmm1, input_a_imag15_vmm1, input_a_imag16_vmm1,
input_a_real1_vmm2, input_a_real2_vmm2,  input_a_real3_vmm2,  input_a_real4_vmm2,  input_a_real5_vmm2,  input_a_real6_vmm2,  input_a_real7_vmm2,  input_a_real8_vmm2,
input_a_imag1_vmm2, input_a_imag2_vmm2,  input_a_imag3_vmm2,  input_a_imag4_vmm2,  input_a_imag5_vmm2,  input_a_imag6_vmm2,  input_a_imag7_vmm2,  input_a_imag8_vmm2,
input_a_real9_vmm2, input_a_real10_vmm2, input_a_real11_vmm2, input_a_real12_vmm2, input_a_real13_vmm2, input_a_real14_vmm2, input_a_real15_vmm2, input_a_real16_vmm2,
input_a_imag9_vmm2, input_a_imag10_vmm2, input_a_imag11_vmm2, input_a_imag12_vmm2, input_a_imag13_vmm2, input_a_imag14_vmm2, input_a_imag15_vmm2, input_a_imag16_vmm2,
input_a_real1_vmm3, input_a_real2_vmm3,  input_a_real3_vmm3,  input_a_real4_vmm3,  input_a_real5_vmm3,  input_a_real6_vmm3,  input_a_real7_vmm3,  input_a_real8_vmm3,
input_a_imag1_vmm3, input_a_imag2_vmm3,  input_a_imag3_vmm3,  input_a_imag4_vmm3,  input_a_imag5_vmm3,  input_a_imag6_vmm3,  input_a_imag7_vmm3,  input_a_imag8_vmm3,
input_a_real9_vmm3, input_a_real10_vmm3, input_a_real11_vmm3, input_a_real12_vmm3, input_a_real13_vmm3, input_a_real14_vmm3, input_a_real15_vmm3, input_a_real16_vmm3,
input_a_imag9_vmm3, input_a_imag10_vmm3, input_a_imag11_vmm3, input_a_imag12_vmm3, input_a_imag13_vmm3, input_a_imag14_vmm3, input_a_imag15_vmm3, input_a_imag16_vmm3,
output_z_real1_0_level6,
output_z_imag1_0_level6
);

input CLK, rst;
input [15:0] input_a_real1_vmm0, input_a_real2_vmm0,  input_a_real3_vmm0,  input_a_real4_vmm0,  input_a_real5_vmm0,  input_a_real6_vmm0,  input_a_real7_vmm0,  input_a_real8_vmm0;
input [15:0] input_a_imag1_vmm0, input_a_imag2_vmm0,  input_a_imag3_vmm0,  input_a_imag4_vmm0,  input_a_imag5_vmm0,  input_a_imag6_vmm0,  input_a_imag7_vmm0,  input_a_imag8_vmm0;
input [15:0] input_a_real9_vmm0, input_a_real10_vmm0, input_a_real11_vmm0, input_a_real12_vmm0, input_a_real13_vmm0, input_a_real14_vmm0, input_a_real15_vmm0, input_a_real16_vmm0;
input [15:0] input_a_imag9_vmm0, input_a_imag10_vmm0, input_a_imag11_vmm0, input_a_imag12_vmm0, input_a_imag13_vmm0, input_a_imag14_vmm0, input_a_imag15_vmm0, input_a_imag16_vmm0;
wire [15:0] output_z_real1_0_level1, output_z_real2_0_level1,  output_z_real3_0_level1,  output_z_real4_0_level1,  output_z_real5_0_level1,  output_z_real6_0_level1,  output_z_real7_0_level1,  output_z_real8_0_level1;
wire [15:0] output_z_imag1_0_level1, output_z_imag2_0_level1,  output_z_imag3_0_level1,  output_z_imag4_0_level1,  output_z_imag5_0_level1,  output_z_imag6_0_level1,  output_z_imag7_0_level1,  output_z_imag8_0_level1;

input [15:0] input_a_real1_vmm1, input_a_real2_vmm1,  input_a_real3_vmm1,  input_a_real4_vmm1,  input_a_real5_vmm1,  input_a_real6_vmm1,  input_a_real7_vmm1,  input_a_real8_vmm1;
input [15:0] input_a_imag1_vmm1, input_a_imag2_vmm1,  input_a_imag3_vmm1,  input_a_imag4_vmm1,  input_a_imag5_vmm1,  input_a_imag6_vmm1,  input_a_imag7_vmm1,  input_a_imag8_vmm1;
input [15:0] input_a_real9_vmm1, input_a_real10_vmm1, input_a_real11_vmm1, input_a_real12_vmm1, input_a_real13_vmm1, input_a_real14_vmm1, input_a_real15_vmm1, input_a_real16_vmm1;
input [15:0] input_a_imag9_vmm1, input_a_imag10_vmm1, input_a_imag11_vmm1, input_a_imag12_vmm1, input_a_imag13_vmm1, input_a_imag14_vmm1, input_a_imag15_vmm1, input_a_imag16_vmm1;
wire [15:0] output_z_real1_1_level1, output_z_real2_1_level1,  output_z_real3_1_level1,  output_z_real4_1_level1,  output_z_real5_1_level1,  output_z_real6_1_level1,  output_z_real7_1_level1,  output_z_real8_1_level1;
wire [15:0] output_z_imag1_1_level1, output_z_imag2_1_level1,  output_z_imag3_1_level1,  output_z_imag4_1_level1,  output_z_imag5_1_level1,  output_z_imag6_1_level1,  output_z_imag7_1_level1,  output_z_imag8_1_level1;

input [15:0] input_a_real1_vmm2, input_a_real2_vmm2,  input_a_real3_vmm2,  input_a_real4_vmm2,  input_a_real5_vmm2,  input_a_real6_vmm2,  input_a_real7_vmm2,  input_a_real8_vmm2;
input [15:0] input_a_imag1_vmm2, input_a_imag2_vmm2,  input_a_imag3_vmm2,  input_a_imag4_vmm2,  input_a_imag5_vmm2,  input_a_imag6_vmm2,  input_a_imag7_vmm2,  input_a_imag8_vmm2;
input [15:0] input_a_real9_vmm2, input_a_real10_vmm2, input_a_real11_vmm2, input_a_real12_vmm2, input_a_real13_vmm2, input_a_real14_vmm2, input_a_real15_vmm2, input_a_real16_vmm2;
input [15:0] input_a_imag9_vmm2, input_a_imag10_vmm2, input_a_imag11_vmm2, input_a_imag12_vmm2, input_a_imag13_vmm2, input_a_imag14_vmm2, input_a_imag15_vmm2, input_a_imag16_vmm2;
wire [15:0] output_z_real1_2_level1, output_z_real2_2_level1,  output_z_real3_2_level1,  output_z_real4_2_level1,  output_z_real5_2_level1,  output_z_real6_2_level1,  output_z_real7_2_level1,  output_z_real8_2_level1;
wire [15:0] output_z_imag1_2_level1, output_z_imag2_2_level1,  output_z_imag3_2_level1,  output_z_imag4_2_level1,  output_z_imag5_2_level1,  output_z_imag6_2_level1,  output_z_imag7_2_level1,  output_z_imag8_2_level1;

input [15:0] input_a_real1_vmm3, input_a_real2_vmm3,  input_a_real3_vmm3,  input_a_real4_vmm3,  input_a_real5_vmm3,  input_a_real6_vmm3,  input_a_real7_vmm3,  input_a_real8_vmm3;
input [15:0] input_a_imag1_vmm3, input_a_imag2_vmm3,  input_a_imag3_vmm3,  input_a_imag4_vmm3,  input_a_imag5_vmm3,  input_a_imag6_vmm3,  input_a_imag7_vmm3,  input_a_imag8_vmm3;
input [15:0] input_a_real9_vmm3, input_a_real10_vmm3, input_a_real11_vmm3, input_a_real12_vmm3, input_a_real13_vmm3, input_a_real14_vmm3, input_a_real15_vmm3, input_a_real16_vmm3;
input [15:0] input_a_imag9_vmm3, input_a_imag10_vmm3, input_a_imag11_vmm3, input_a_imag12_vmm3, input_a_imag13_vmm3, input_a_imag14_vmm3, input_a_imag15_vmm3, input_a_imag16_vmm3;
wire [15:0] output_z_real1_3_level1, output_z_real2_3_level1,  output_z_real3_3_level1,  output_z_real4_3_level1,  output_z_real5_3_level1,  output_z_real6_3_level1,  output_z_real7_3_level1,  output_z_real8_3_level1;
wire [15:0] output_z_imag1_3_level1, output_z_imag2_3_level1,  output_z_imag3_3_level1,  output_z_imag4_3_level1,  output_z_imag5_3_level1,  output_z_imag6_3_level1,  output_z_imag7_3_level1,  output_z_imag8_3_level1;

complex_adder DUT_ADDER0_1_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real1_vmm0), .input_b_real(input_a_real2_vmm0), .output_z_real(output_z_real1_0_level1),
.input_a_imag(input_a_imag1_vmm0), .input_b_imag(input_a_imag2_vmm0), .output_z_imag(output_z_imag1_0_level1)
);


complex_adder DUT_ADDER0_2_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real3_vmm0), .input_b_real(input_a_real4_vmm0), .output_z_real(output_z_real2_0_level1),
.input_a_imag(input_a_imag3_vmm0), .input_b_imag(input_a_imag4_vmm0), .output_z_imag(output_z_imag2_0_level1)
);


complex_adder DUT_ADDER0_3_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real5_vmm0), .input_b_real(input_a_real6_vmm0), .output_z_real(output_z_real3_0_level1),
.input_a_imag(input_a_imag5_vmm0), .input_b_imag(input_a_imag6_vmm0), .output_z_imag(output_z_imag3_0_level1)
);


complex_adder DUT_ADDER0_4_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real7_vmm0), .input_b_real(input_a_real8_vmm0), .output_z_real(output_z_real4_0_level1),
.input_a_imag(input_a_imag7_vmm0), .input_b_imag(input_a_imag8_vmm0), .output_z_imag(output_z_imag4_0_level1)
);


complex_adder DUT_ADDER0_5_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real9_vmm0), .input_b_real(input_a_real10_vmm0), .output_z_real(output_z_real5_0_level1),
.input_a_imag(input_a_imag9_vmm0), .input_b_imag(input_a_imag10_vmm0), .output_z_imag(output_z_imag5_0_level1)
);


complex_adder DUT_ADDER0_6_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real11_vmm0), .input_b_real(input_a_real12_vmm0), .output_z_real(output_z_real6_0_level1),
.input_a_imag(input_a_imag11_vmm0), .input_b_imag(input_a_imag12_vmm0), .output_z_imag(output_z_imag6_0_level1)
);


complex_adder DUT_ADDER0_7_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real13_vmm0), .input_b_real(input_a_real14_vmm0), .output_z_real(output_z_real7_0_level1),
.input_a_imag(input_a_imag13_vmm0), .input_b_imag(input_a_imag14_vmm0), .output_z_imag(output_z_imag7_0_level1)
);


complex_adder DUT_ADDER0_8_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real15_vmm0), .input_b_real(input_a_real16_vmm0), .output_z_real(output_z_real8_0_level1),
.input_a_imag(input_a_imag15_vmm0), .input_b_imag(input_a_imag16_vmm0), .output_z_imag(output_z_imag8_0_level1)
);


complex_adder DUT_ADDER1_1_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real1_vmm1), .input_b_real(input_a_real2_vmm1), .output_z_real(output_z_real1_1_level1),
.input_a_imag(input_a_imag1_vmm1), .input_b_imag(input_a_imag2_vmm1), .output_z_imag(output_z_imag1_1_level1)
);


complex_adder DUT_ADDER1_2_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real3_vmm1), .input_b_real(input_a_real4_vmm1), .output_z_real(output_z_real2_1_level1),
.input_a_imag(input_a_imag3_vmm1), .input_b_imag(input_a_imag4_vmm1), .output_z_imag(output_z_imag2_1_level1)
);


complex_adder DUT_ADDER1_3_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real5_vmm1), .input_b_real(input_a_real6_vmm1), .output_z_real(output_z_real3_1_level1),
.input_a_imag(input_a_imag5_vmm1), .input_b_imag(input_a_imag6_vmm1), .output_z_imag(output_z_imag3_1_level1)
);


complex_adder DUT_ADDER1_4_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real7_vmm1), .input_b_real(input_a_real8_vmm1), .output_z_real(output_z_real4_1_level1),
.input_a_imag(input_a_imag7_vmm1), .input_b_imag(input_a_imag8_vmm1), .output_z_imag(output_z_imag4_1_level1)
);


complex_adder DUT_ADDER1_5_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real9_vmm1), .input_b_real(input_a_real10_vmm1), .output_z_real(output_z_real5_1_level1),
.input_a_imag(input_a_imag9_vmm1), .input_b_imag(input_a_imag10_vmm1), .output_z_imag(output_z_imag5_1_level1)
);


complex_adder DUT_ADDER1_6_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real11_vmm1), .input_b_real(input_a_real12_vmm1), .output_z_real(output_z_real6_1_level1),
.input_a_imag(input_a_imag11_vmm1), .input_b_imag(input_a_imag12_vmm1), .output_z_imag(output_z_imag6_1_level1)
);


complex_adder DUT_ADDER1_7_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real13_vmm1), .input_b_real(input_a_real14_vmm1), .output_z_real(output_z_real7_1_level1),
.input_a_imag(input_a_imag13_vmm1), .input_b_imag(input_a_imag14_vmm1), .output_z_imag(output_z_imag7_1_level1)
);


complex_adder DUT_ADDER1_8_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real15_vmm1), .input_b_real(input_a_real16_vmm1), .output_z_real(output_z_real8_1_level1),
.input_a_imag(input_a_imag15_vmm1), .input_b_imag(input_a_imag16_vmm1), .output_z_imag(output_z_imag8_1_level1)
);


complex_adder DUT_ADDER2_1_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real1_vmm2), .input_b_real(input_a_real2_vmm2), .output_z_real(output_z_real1_2_level1),
.input_a_imag(input_a_imag1_vmm2), .input_b_imag(input_a_imag2_vmm2), .output_z_imag(output_z_imag1_2_level1)
);


complex_adder DUT_ADDER2_2_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real3_vmm2), .input_b_real(input_a_real4_vmm2), .output_z_real(output_z_real2_2_level1),
.input_a_imag(input_a_imag3_vmm2), .input_b_imag(input_a_imag4_vmm2), .output_z_imag(output_z_imag2_2_level1)
);


complex_adder DUT_ADDER2_3_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real5_vmm2), .input_b_real(input_a_real6_vmm2), .output_z_real(output_z_real3_2_level1),
.input_a_imag(input_a_imag5_vmm2), .input_b_imag(input_a_imag6_vmm2), .output_z_imag(output_z_imag3_2_level1)
);


complex_adder DUT_ADDER2_4_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real7_vmm2), .input_b_real(input_a_real8_vmm2), .output_z_real(output_z_real4_2_level1),
.input_a_imag(input_a_imag7_vmm2), .input_b_imag(input_a_imag8_vmm2), .output_z_imag(output_z_imag4_2_level1)
);


complex_adder DUT_ADDER2_5_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real9_vmm2), .input_b_real(input_a_real10_vmm2), .output_z_real(output_z_real5_2_level1),
.input_a_imag(input_a_imag9_vmm2), .input_b_imag(input_a_imag10_vmm2), .output_z_imag(output_z_imag5_2_level1)
);


complex_adder DUT_ADDER2_6_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real11_vmm2), .input_b_real(input_a_real12_vmm2), .output_z_real(output_z_real6_2_level1),
.input_a_imag(input_a_imag11_vmm2), .input_b_imag(input_a_imag12_vmm2), .output_z_imag(output_z_imag6_2_level1)
);


complex_adder DUT_ADDER2_7_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real13_vmm2), .input_b_real(input_a_real14_vmm2), .output_z_real(output_z_real7_2_level1),
.input_a_imag(input_a_imag13_vmm2), .input_b_imag(input_a_imag14_vmm2), .output_z_imag(output_z_imag7_2_level1)
);


complex_adder DUT_ADDER2_8_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real15_vmm2), .input_b_real(input_a_real16_vmm2), .output_z_real(output_z_real8_2_level1),
.input_a_imag(input_a_imag15_vmm2), .input_b_imag(input_a_imag16_vmm2), .output_z_imag(output_z_imag8_2_level1)
);


complex_adder DUT_ADDER3_1_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real1_vmm3), .input_b_real(input_a_real2_vmm3), .output_z_real(output_z_real1_3_level1),
.input_a_imag(input_a_imag1_vmm3), .input_b_imag(input_a_imag2_vmm3), .output_z_imag(output_z_imag1_3_level1)
);


complex_adder DUT_ADDER3_2_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real3_vmm3), .input_b_real(input_a_real4_vmm3), .output_z_real(output_z_real2_3_level1),
.input_a_imag(input_a_imag3_vmm3), .input_b_imag(input_a_imag4_vmm3), .output_z_imag(output_z_imag2_3_level1)
);


complex_adder DUT_ADDER3_3_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real5_vmm3), .input_b_real(input_a_real6_vmm3), .output_z_real(output_z_real3_3_level1),
.input_a_imag(input_a_imag5_vmm3), .input_b_imag(input_a_imag6_vmm3), .output_z_imag(output_z_imag3_3_level1)
);


complex_adder DUT_ADDER3_4_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real7_vmm3), .input_b_real(input_a_real8_vmm3), .output_z_real(output_z_real4_3_level1),
.input_a_imag(input_a_imag7_vmm3), .input_b_imag(input_a_imag8_vmm3), .output_z_imag(output_z_imag4_3_level1)
);


complex_adder DUT_ADDER3_5_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real9_vmm3), .input_b_real(input_a_real10_vmm3), .output_z_real(output_z_real5_3_level1),
.input_a_imag(input_a_imag9_vmm3), .input_b_imag(input_a_imag10_vmm3), .output_z_imag(output_z_imag5_3_level1)
);


complex_adder DUT_ADDER3_6_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real11_vmm3), .input_b_real(input_a_real12_vmm3), .output_z_real(output_z_real6_3_level1),
.input_a_imag(input_a_imag11_vmm3), .input_b_imag(input_a_imag12_vmm3), .output_z_imag(output_z_imag6_3_level1)
);


complex_adder DUT_ADDER3_7_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real13_vmm3), .input_b_real(input_a_real14_vmm3), .output_z_real(output_z_real7_3_level1),
.input_a_imag(input_a_imag13_vmm3), .input_b_imag(input_a_imag14_vmm3), .output_z_imag(output_z_imag7_3_level1)
);


complex_adder DUT_ADDER3_8_level1(
.CLK(CLK), .rst(rst), 
.input_a_real(input_a_real15_vmm3), .input_b_real(input_a_real16_vmm3), .output_z_real(output_z_real8_3_level1),
.input_a_imag(input_a_imag15_vmm3), .input_b_imag(input_a_imag16_vmm3), .output_z_imag(output_z_imag8_3_level1)
);


wire [15:0] output_z_real1_0_level2, output_z_real2_0_level2,  output_z_real3_0_level2,  output_z_real4_0_level2;
wire [15:0] output_z_imag1_0_level2, output_z_imag2_0_level2,  output_z_imag3_0_level2,  output_z_imag4_0_level2;


wire [15:0] output_z_real1_1_level2, output_z_real2_1_level2,  output_z_real3_1_level2,  output_z_real4_1_level2;
wire [15:0] output_z_imag1_1_level2, output_z_imag2_1_level2,  output_z_imag3_1_level2,  output_z_imag4_1_level2;


wire [15:0] output_z_real1_2_level2, output_z_real2_2_level2,  output_z_real3_2_level2,  output_z_real4_2_level2;
wire [15:0] output_z_imag1_2_level2, output_z_imag2_2_level2,  output_z_imag3_2_level2,  output_z_imag4_2_level2;


wire [15:0] output_z_real1_3_level2, output_z_real2_3_level2,  output_z_real3_3_level2,  output_z_real4_3_level2;
wire [15:0] output_z_imag1_3_level2, output_z_imag2_3_level2,  output_z_imag3_3_level2,  output_z_imag4_3_level2;


complex_adder DUT_ADDER0_1_level2(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real1_0_level1), .input_b_real(output_z_real2_0_level1), .output_z_real(output_z_real1_0_level2),
.input_a_imag(output_z_imag1_0_level1), .input_b_imag(output_z_imag2_0_level1), .output_z_imag(output_z_imag1_0_level2)
);


complex_adder DUT_ADDER0_2_level2(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real3_0_level1), .input_b_real(output_z_real4_0_level1), .output_z_real(output_z_real2_0_level2),
.input_a_imag(output_z_imag3_0_level1), .input_b_imag(output_z_imag4_0_level1), .output_z_imag(output_z_imag2_0_level2)
);


complex_adder DUT_ADDER0_3_level2(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real5_0_level1), .input_b_real(output_z_real6_0_level1), .output_z_real(output_z_real3_0_level2),
.input_a_imag(output_z_imag5_0_level1), .input_b_imag(output_z_imag6_0_level1), .output_z_imag(output_z_imag3_0_level2)
);


complex_adder DUT_ADDER0_4_level2(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real7_0_level1), .input_b_real(output_z_real8_0_level1), .output_z_real(output_z_real4_0_level2),
.input_a_imag(output_z_imag7_0_level1), .input_b_imag(output_z_imag8_0_level1), .output_z_imag(output_z_imag4_0_level2)
);


complex_adder DUT_ADDER1_1_level2(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real1_1_level1), .input_b_real(output_z_real2_1_level1), .output_z_real(output_z_real1_1_level2),
.input_a_imag(output_z_imag1_1_level1), .input_b_imag(output_z_imag2_1_level1), .output_z_imag(output_z_imag1_1_level2)
);


complex_adder DUT_ADDER1_2_level2(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real3_1_level1), .input_b_real(output_z_real4_1_level1), .output_z_real(output_z_real2_1_level2),
.input_a_imag(output_z_imag3_1_level1), .input_b_imag(output_z_imag4_1_level1), .output_z_imag(output_z_imag2_1_level2)
);


complex_adder DUT_ADDER1_3_level2(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real5_1_level1), .input_b_real(output_z_real6_1_level1), .output_z_real(output_z_real3_1_level2),
.input_a_imag(output_z_imag5_1_level1), .input_b_imag(output_z_imag6_1_level1), .output_z_imag(output_z_imag3_1_level2)
);


complex_adder DUT_ADDER1_4_level2(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real7_1_level1), .input_b_real(output_z_real8_1_level1), .output_z_real(output_z_real4_1_level2),
.input_a_imag(output_z_imag7_1_level1), .input_b_imag(output_z_imag8_1_level1), .output_z_imag(output_z_imag4_1_level2)
);


complex_adder DUT_ADDER2_1_level2(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real1_2_level1), .input_b_real(output_z_real2_2_level1), .output_z_real(output_z_real1_2_level2),
.input_a_imag(output_z_imag1_2_level1), .input_b_imag(output_z_imag2_2_level1), .output_z_imag(output_z_imag1_2_level2)
);


complex_adder DUT_ADDER2_2_level2(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real3_2_level1), .input_b_real(output_z_real4_2_level1), .output_z_real(output_z_real2_2_level2),
.input_a_imag(output_z_imag3_2_level1), .input_b_imag(output_z_imag4_2_level1), .output_z_imag(output_z_imag2_2_level2)
);


complex_adder DUT_ADDER2_3_level2(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real5_2_level1), .input_b_real(output_z_real6_2_level1), .output_z_real(output_z_real3_2_level2),
.input_a_imag(output_z_imag5_2_level1), .input_b_imag(output_z_imag6_2_level1), .output_z_imag(output_z_imag3_2_level2)
);


complex_adder DUT_ADDER2_4_level2(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real7_2_level1), .input_b_real(output_z_real8_2_level1), .output_z_real(output_z_real4_2_level2),
.input_a_imag(output_z_imag7_2_level1), .input_b_imag(output_z_imag8_2_level1), .output_z_imag(output_z_imag4_2_level2)
);


complex_adder DUT_ADDER3_1_level2(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real1_3_level1), .input_b_real(output_z_real2_3_level1), .output_z_real(output_z_real1_3_level2),
.input_a_imag(output_z_imag1_3_level1), .input_b_imag(output_z_imag2_3_level1), .output_z_imag(output_z_imag1_3_level2)
);


complex_adder DUT_ADDER3_2_level2(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real3_3_level1), .input_b_real(output_z_real4_3_level1), .output_z_real(output_z_real2_3_level2),
.input_a_imag(output_z_imag3_3_level1), .input_b_imag(output_z_imag4_3_level1), .output_z_imag(output_z_imag2_3_level2)
);


complex_adder DUT_ADDER3_3_level2(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real5_3_level1), .input_b_real(output_z_real6_3_level1), .output_z_real(output_z_real3_3_level2),
.input_a_imag(output_z_imag5_3_level1), .input_b_imag(output_z_imag6_3_level1), .output_z_imag(output_z_imag3_3_level2)
);


complex_adder DUT_ADDER3_4_level2(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real7_3_level1), .input_b_real(output_z_real8_3_level1), .output_z_real(output_z_real4_3_level2),
.input_a_imag(output_z_imag7_3_level1), .input_b_imag(output_z_imag8_3_level1), .output_z_imag(output_z_imag4_3_level2)
);


wire [15:0] output_z_real1_0_level3, output_z_real2_0_level3;
wire [15:0] output_z_imag1_0_level3, output_z_imag2_0_level3;


wire [15:0] output_z_real1_1_level3, output_z_real2_1_level3;
wire [15:0] output_z_imag1_1_level3, output_z_imag2_1_level3;


wire [15:0] output_z_real1_2_level3, output_z_real2_2_level3;
wire [15:0] output_z_imag1_2_level3, output_z_imag2_2_level3;


wire [15:0] output_z_real1_3_level3, output_z_real2_3_level3;
wire [15:0] output_z_imag1_3_level3, output_z_imag2_3_level3;


complex_adder DUT_ADDER0_1_level3(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real1_0_level2), .input_b_real(output_z_real2_0_level2), .output_z_real(output_z_real1_0_level3),
.input_a_imag(output_z_imag1_0_level2), .input_b_imag(output_z_imag2_0_level2), .output_z_imag(output_z_imag1_0_level3)
);


complex_adder DUT_ADDER0_2_level3(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real3_0_level2), .input_b_real(output_z_real4_0_level2), .output_z_real(output_z_real2_0_level3),
.input_a_imag(output_z_imag3_0_level2), .input_b_imag(output_z_imag4_0_level2), .output_z_imag(output_z_imag2_0_level3)
);


complex_adder DUT_ADDER1_1_level3(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real1_1_level2), .input_b_real(output_z_real2_1_level2), .output_z_real(output_z_real1_1_level3),
.input_a_imag(output_z_imag1_1_level2), .input_b_imag(output_z_imag2_1_level2), .output_z_imag(output_z_imag1_1_level3)
);


complex_adder DUT_ADDER1_2_level3(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real3_1_level2), .input_b_real(output_z_real4_1_level2), .output_z_real(output_z_real2_1_level3),
.input_a_imag(output_z_imag3_1_level2), .input_b_imag(output_z_imag4_1_level2), .output_z_imag(output_z_imag2_1_level3)
);


complex_adder DUT_ADDER2_1_level3(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real1_2_level2), .input_b_real(output_z_real2_2_level2), .output_z_real(output_z_real1_2_level3),
.input_a_imag(output_z_imag1_2_level2), .input_b_imag(output_z_imag2_2_level2), .output_z_imag(output_z_imag1_2_level3)
);


complex_adder DUT_ADDER2_2_level3(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real3_2_level2), .input_b_real(output_z_real4_2_level2), .output_z_real(output_z_real2_2_level3),
.input_a_imag(output_z_imag3_2_level2), .input_b_imag(output_z_imag4_2_level2), .output_z_imag(output_z_imag2_2_level3)
);


complex_adder DUT_ADDER3_1_level3(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real1_3_level2), .input_b_real(output_z_real2_3_level2), .output_z_real(output_z_real1_3_level3),
.input_a_imag(output_z_imag1_3_level2), .input_b_imag(output_z_imag2_3_level2), .output_z_imag(output_z_imag1_3_level3)
);


complex_adder DUT_ADDER3_2_level3(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real3_3_level2), .input_b_real(output_z_real4_3_level2), .output_z_real(output_z_real2_3_level3),
.input_a_imag(output_z_imag3_3_level2), .input_b_imag(output_z_imag4_3_level2), .output_z_imag(output_z_imag2_3_level3)
);


wire [15:0] output_z_real1_0_level4;
wire [15:0] output_z_imag1_0_level4;
wire [15:0] output_z_real1_1_level4;
wire [15:0] output_z_imag1_1_level4;
wire [15:0] output_z_real1_2_level4;
wire [15:0] output_z_imag1_2_level4;
wire [15:0] output_z_real1_3_level4;
wire [15:0] output_z_imag1_3_level4;


complex_adder DUT_ADDER0_1_level4(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real1_0_level3), .input_b_real(output_z_real2_0_level3), .output_z_real(output_z_real1_0_level4),
.input_a_imag(output_z_imag1_0_level3), .input_b_imag(output_z_imag2_0_level3), .output_z_imag(output_z_imag1_0_level4)
);


complex_adder DUT_ADDER1_1_level4(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real1_1_level3), .input_b_real(output_z_real2_1_level3), .output_z_real(output_z_real1_1_level4),
.input_a_imag(output_z_imag1_1_level3), .input_b_imag(output_z_imag2_1_level3), .output_z_imag(output_z_imag1_1_level4)
);


complex_adder DUT_ADDER2_1_level4(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real1_2_level3), .input_b_real(output_z_real2_2_level3), .output_z_real(output_z_real1_2_level4),
.input_a_imag(output_z_imag1_2_level3), .input_b_imag(output_z_imag2_2_level3), .output_z_imag(output_z_imag1_2_level4)
);


complex_adder DUT_ADDER3_1_level4(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real1_3_level3), .input_b_real(output_z_real2_3_level3), .output_z_real(output_z_real1_3_level4),
.input_a_imag(output_z_imag1_3_level3), .input_b_imag(output_z_imag2_3_level3), .output_z_imag(output_z_imag1_3_level4)
);

wire [15:0] output_z_real1_0_level5;
wire [15:0] output_z_imag1_0_level5;
wire [15:0] output_z_real1_1_level5;
wire [15:0] output_z_imag1_1_level5;

complex_adder DUT_ADDER0_level5(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real1_0_level4), .input_b_real(output_z_real1_1_level4), .output_z_real(output_z_real1_0_level5),
.input_a_imag(output_z_imag1_0_level4), .input_b_imag(output_z_imag1_1_level4), .output_z_imag(output_z_imag1_0_level5)
);

complex_adder DUT_ADDER1_level5(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real1_2_level4), .input_b_real(output_z_real1_3_level4), .output_z_real(output_z_real1_1_level5),
.input_a_imag(output_z_imag1_2_level4), .input_b_imag(output_z_imag1_3_level4), .output_z_imag(output_z_imag1_1_level5)
);

output [15:0] output_z_real1_0_level6;
output [15:0] output_z_imag1_0_level6;

complex_adder DUT_ADDER0_level6(
.CLK(CLK), .rst(rst), 
.input_a_real(output_z_real1_0_level5), .input_b_real(output_z_real1_1_level5), .output_z_real(output_z_real1_0_level6),
.input_a_imag(output_z_imag1_0_level5), .input_b_imag(output_z_imag1_1_level5), .output_z_imag(output_z_imag1_0_level6)
);

endmodule
