
module memory_rom_36(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbe52add1;
    11'b00000000001: data <= 32'hbb291b46;
    11'b00000000010: data <= 32'h3b6e2dc5;
    11'b00000000011: data <= 32'h3e783b8f;
    11'b00000000100: data <= 32'h2a823ee7;
    11'b00000000101: data <= 32'hbf6a3dcd;
    11'b00000000110: data <= 32'hbed239a3;
    11'b00000000111: data <= 32'h2e423853;
    11'b00000001000: data <= 32'h3cec3882;
    11'b00000001001: data <= 32'h3b2fb478;
    11'b00000001010: data <= 32'h3871bdc1;
    11'b00000001011: data <= 32'h3cc4bc92;
    11'b00000001100: data <= 32'h3f1e39ae;
    11'b00000001101: data <= 32'h3ca23f4e;
    11'b00000001110: data <= 32'haa1c38ca;
    11'b00000001111: data <= 32'hb8b9be0d;
    11'b00000010000: data <= 32'hb8b5c012;
    11'b00000010001: data <= 32'hbb31bb7b;
    11'b00000010010: data <= 32'hbcc4b492;
    11'b00000010011: data <= 32'hb65cbb45;
    11'b00000010100: data <= 32'h3c18bd28;
    11'b00000010101: data <= 32'h3c79b2a2;
    11'b00000010110: data <= 32'hb96e3d41;
    11'b00000010111: data <= 32'hc09a3eb9;
    11'b00000011000: data <= 32'hbf363c28;
    11'b00000011001: data <= 32'haf873892;
    11'b00000011010: data <= 32'h3711367b;
    11'b00000011011: data <= 32'hb561b14d;
    11'b00000011100: data <= 32'hb752ba4e;
    11'b00000011101: data <= 32'h3bddb2ea;
    11'b00000011110: data <= 32'h40ab3d8b;
    11'b00000011111: data <= 32'h3fa34014;
    11'b00000100000: data <= 32'h3636398f;
    11'b00000100001: data <= 32'hb762bc1d;
    11'b00000100010: data <= 32'hb585bc84;
    11'b00000100011: data <= 32'hb338b1bd;
    11'b00000100100: data <= 32'hb41cb50c;
    11'b00000100101: data <= 32'h34d7bf1c;
    11'b00000100110: data <= 32'h3cc5c0d7;
    11'b00000100111: data <= 32'h3bebbbc1;
    11'b00000101000: data <= 32'hb8ca3c1b;
    11'b00000101001: data <= 32'hbf543ddc;
    11'b00000101010: data <= 32'hbd77380e;
    11'b00000101011: data <= 32'hb58fb253;
    11'b00000101100: data <= 32'hb8f8b093;
    11'b00000101101: data <= 32'hbed5b0f9;
    11'b00000101110: data <= 32'hbda9b5fc;
    11'b00000101111: data <= 32'h397e2f40;
    11'b00000110000: data <= 32'h40a63d62;
    11'b00000110001: data <= 32'h3ec63f99;
    11'b00000110010: data <= 32'had0f3c24;
    11'b00000110011: data <= 32'hba1b2a80;
    11'b00000110100: data <= 32'hae603466;
    11'b00000110101: data <= 32'h378d3a6c;
    11'b00000110110: data <= 32'h368fb057;
    11'b00000110111: data <= 32'h38a1c031;
    11'b00000111000: data <= 32'h3cefc14c;
    11'b00000111001: data <= 32'h3d3fbb1f;
    11'b00000111010: data <= 32'h351c3c4c;
    11'b00000111011: data <= 32'hb8dd3c2a;
    11'b00000111100: data <= 32'hb84bb61a;
    11'b00000111101: data <= 32'hb5ffbc4e;
    11'b00000111110: data <= 32'hbd32b899;
    11'b00000111111: data <= 32'hc0cfb27c;
    11'b00001000000: data <= 32'hbef2b82a;
    11'b00001000001: data <= 32'h3844b804;
    11'b00001000010: data <= 32'h3f723728;
    11'b00001000011: data <= 32'h3a5a3d60;
    11'b00001000100: data <= 32'hbc003d3f;
    11'b00001000101: data <= 32'hbcc73c23;
    11'b00001000110: data <= 32'h0f6d3d5f;
    11'b00001000111: data <= 32'h391d3dbe;
    11'b00001001000: data <= 32'h32332f8d;
    11'b00001001001: data <= 32'h2b22bf05;
    11'b00001001010: data <= 32'h3bbbbfcc;
    11'b00001001011: data <= 32'h3f34afbc;
    11'b00001001100: data <= 32'h3dfe3d84;
    11'b00001001101: data <= 32'h394939bc;
    11'b00001001110: data <= 32'h3394bb61;
    11'b00001001111: data <= 32'hb11dbd2b;
    11'b00001010000: data <= 32'hbcdeb665;
    11'b00001010001: data <= 32'hc026b056;
    11'b00001010010: data <= 32'hbd20bc63;
    11'b00001010011: data <= 32'h3902bee1;
    11'b00001010100: data <= 32'h3d4bbab3;
    11'b00001010101: data <= 32'hac1538f6;
    11'b00001010110: data <= 32'hbe583d24;
    11'b00001010111: data <= 32'hbd233d3b;
    11'b00001011000: data <= 32'h21093dd5;
    11'b00001011001: data <= 32'h313f3d77;
    11'b00001011010: data <= 32'hbb033428;
    11'b00001011011: data <= 32'hbc55bc50;
    11'b00001011100: data <= 32'h36e0bb6b;
    11'b00001011101: data <= 32'h4022396d;
    11'b00001011110: data <= 32'h40573e69;
    11'b00001011111: data <= 32'h3cd23904;
    11'b00001100000: data <= 32'h380eb9cc;
    11'b00001100001: data <= 32'h30c6b865;
    11'b00001100010: data <= 32'hb82f378a;
    11'b00001100011: data <= 32'hbc50314c;
    11'b00001100100: data <= 32'hb7acbe9e;
    11'b00001100101: data <= 32'h3a92c184;
    11'b00001100110: data <= 32'h3c30beeb;
    11'b00001100111: data <= 32'hb3ca307d;
    11'b00001101000: data <= 32'hbd203bad;
    11'b00001101001: data <= 32'hba013a06;
    11'b00001101010: data <= 32'h2e87394b;
    11'b00001101011: data <= 32'hb89e39fa;
    11'b00001101100: data <= 32'hc04a33a4;
    11'b00001101101: data <= 32'hc060b868;
    11'b00001101110: data <= 32'haed6b5e1;
    11'b00001101111: data <= 32'h3f9a3a71;
    11'b00001110000: data <= 32'h3fb33d90;
    11'b00001110001: data <= 32'h39f53951;
    11'b00001110010: data <= 32'h319327f6;
    11'b00001110011: data <= 32'h35ed39f5;
    11'b00001110100: data <= 32'h34273e74;
    11'b00001110101: data <= 32'hb2c138ff;
    11'b00001110110: data <= 32'ha878bf1b;
    11'b00001110111: data <= 32'h3a8dc1e5;
    11'b00001111000: data <= 32'h3c60bec4;
    11'b00001111001: data <= 32'h35b63176;
    11'b00001111010: data <= 32'hb1a73851;
    11'b00001111011: data <= 32'h33cdb26a;
    11'b00001111100: data <= 32'h3622b62e;
    11'b00001111101: data <= 32'hbc1930dc;
    11'b00001111110: data <= 32'hc1983292;
    11'b00001111111: data <= 32'hc12bb753;
    11'b00010000000: data <= 32'hb545b967;
    11'b00010000001: data <= 32'h3da528be;
    11'b00010000010: data <= 32'h3bc63968;
    11'b00010000011: data <= 32'hb50238e9;
    11'b00010000100: data <= 32'hb6853a0e;
    11'b00010000101: data <= 32'h37643f0f;
    11'b00010000110: data <= 32'h390c40b7;
    11'b00010000111: data <= 32'hb04e3c02;
    11'b00010001000: data <= 32'hb69fbd80;
    11'b00010001001: data <= 32'h3693c068;
    11'b00010001010: data <= 32'h3d02ba8b;
    11'b00010001011: data <= 32'h3d0738d5;
    11'b00010001100: data <= 32'h3c29338a;
    11'b00010001101: data <= 32'h3ca5bb4f;
    11'b00010001110: data <= 32'h3a37bb03;
    11'b00010001111: data <= 32'hbac3316a;
    11'b00010010000: data <= 32'hc0dc3632;
    11'b00010010001: data <= 32'hc021b9b2;
    11'b00010010010: data <= 32'hb075be68;
    11'b00010010011: data <= 32'h3b2abcc0;
    11'b00010010100: data <= 32'ha82db2f4;
    11'b00010010101: data <= 32'hbca035bd;
    11'b00010010110: data <= 32'hb9533b2d;
    11'b00010010111: data <= 32'h38733f65;
    11'b00010011000: data <= 32'h37574088;
    11'b00010011001: data <= 32'hbb433c5a;
    11'b00010011010: data <= 32'hbdedb9b4;
    11'b00010011011: data <= 32'hb4f0bc39;
    11'b00010011100: data <= 32'h3cfe32fc;
    11'b00010011101: data <= 32'h3f0c3c03;
    11'b00010011110: data <= 32'h3e3e2dc6;
    11'b00010011111: data <= 32'h3dd5bbf7;
    11'b00010100000: data <= 32'h3c52b6ed;
    11'b00010100001: data <= 32'hb0cb3ba2;
    11'b00010100010: data <= 32'hbd503af9;
    11'b00010100011: data <= 32'hbc32bbc8;
    11'b00010100100: data <= 32'h337bc0e2;
    11'b00010100101: data <= 32'h38b7c01f;
    11'b00010100110: data <= 32'hb77fba2b;
    11'b00010100111: data <= 32'hbc9aa4f9;
    11'b00010101000: data <= 32'hb38a350f;
    11'b00010101001: data <= 32'h3a933bbb;
    11'b00010101010: data <= 32'h27253ddd;
    11'b00010101011: data <= 32'hbfd43b2e;
    11'b00010101100: data <= 32'hc124b1a1;
    11'b00010101101: data <= 32'hbbb1b436;
    11'b00010101110: data <= 32'h3bc73928;
    11'b00010101111: data <= 32'h3dd73b56;
    11'b00010110000: data <= 32'h3c21a717;
    11'b00010110001: data <= 32'h3be2b86f;
    11'b00010110010: data <= 32'h3c9f38ff;
    11'b00010110011: data <= 32'h390a4028;
    11'b00010110100: data <= 32'hb4023ded;
    11'b00010110101: data <= 32'hb4edbb76;
    11'b00010110110: data <= 32'h3616c118;
    11'b00010110111: data <= 32'h380bbfe3;
    11'b00010111000: data <= 32'hb1c3b92f;
    11'b00010111001: data <= 32'hb4c1b540;
    11'b00010111010: data <= 32'h39e5b910;
    11'b00010111011: data <= 32'h3d1eb44c;
    11'b00010111100: data <= 32'hb2d638a7;
    11'b00010111101: data <= 32'hc0ff398d;
    11'b00010111110: data <= 32'hc1de24d2;
    11'b00010111111: data <= 32'hbc92b444;
    11'b00011000000: data <= 32'h3865309e;
    11'b00011000001: data <= 32'h38063397;
    11'b00011000010: data <= 32'hb219b44d;
    11'b00011000011: data <= 32'h3036ac6d;
    11'b00011000100: data <= 32'h3c423e0c;
    11'b00011000101: data <= 32'h3c4c419f;
    11'b00011000110: data <= 32'h2f903f7b;
    11'b00011000111: data <= 32'hb66fb860;
    11'b00011001000: data <= 32'h279abf23;
    11'b00011001001: data <= 32'h378ebba5;
    11'b00011001010: data <= 32'h373d27fd;
    11'b00011001011: data <= 32'h3a22b734;
    11'b00011001100: data <= 32'h3ea3bd97;
    11'b00011001101: data <= 32'h3ef2bc25;
    11'b00011001110: data <= 32'h128434cf;
    11'b00011001111: data <= 32'hc0313a52;
    11'b00011010000: data <= 32'hc097aaf5;
    11'b00011010001: data <= 32'hb9eebb42;
    11'b00011010010: data <= 32'h327fbb3f;
    11'b00011010011: data <= 32'hb84eb95d;
    11'b00011010100: data <= 32'hbd30b915;
    11'b00011010101: data <= 32'hb6f5a3fb;
    11'b00011010110: data <= 32'h3c2c3e32;
    11'b00011010111: data <= 32'h3c424142;
    11'b00011011000: data <= 32'hb5bf3f27;
    11'b00011011001: data <= 32'hbd17a81c;
    11'b00011011010: data <= 32'hb9a2b8da;
    11'b00011011011: data <= 32'h351b3548;
    11'b00011011100: data <= 32'h3a9539f3;
    11'b00011011101: data <= 32'h3ce6b748;
    11'b00011011110: data <= 32'h3f97be7a;
    11'b00011011111: data <= 32'h3fb3bb24;
    11'b00011100000: data <= 32'h38a73aeb;
    11'b00011100001: data <= 32'hbbbc3d1c;
    11'b00011100010: data <= 32'hbc30b092;
    11'b00011100011: data <= 32'hab50be4a;
    11'b00011100100: data <= 32'h2b40becc;
    11'b00011100101: data <= 32'hbc60bcca;
    11'b00011100110: data <= 32'hbe60bba6;
    11'b00011100111: data <= 32'hb3feb82d;
    11'b00011101000: data <= 32'h3d2d3919;
    11'b00011101001: data <= 32'h3a873e7a;
    11'b00011101010: data <= 32'hbccf3d32;
    11'b00011101011: data <= 32'hc0873556;
    11'b00011101100: data <= 32'hbd6e34a0;
    11'b00011101101: data <= 32'h297d3c3f;
    11'b00011101110: data <= 32'h38663b6c;
    11'b00011101111: data <= 32'h3952b843;
    11'b00011110000: data <= 32'h3cfcbd72;
    11'b00011110001: data <= 32'h3ee8ac3e;
    11'b00011110010: data <= 32'h3cc23f81;
    11'b00011110011: data <= 32'h32593fa0;
    11'b00011110100: data <= 32'h10fbaa86;
    11'b00011110101: data <= 32'h362bbea4;
    11'b00011110110: data <= 32'h2958be4e;
    11'b00011110111: data <= 32'hbbe0bb76;
    11'b00011111000: data <= 32'hbbf2bc21;
    11'b00011111001: data <= 32'h38b6bd3e;
    11'b00011111010: data <= 32'h3f1fb963;
    11'b00011111011: data <= 32'h395936f1;
    11'b00011111100: data <= 32'hbebc3a3b;
    11'b00011111101: data <= 32'hc12e36de;
    11'b00011111110: data <= 32'hbdbd3748;
    11'b00011111111: data <= 32'hb24f3aad;
    11'b00100000000: data <= 32'hb4503686;
    11'b00100000001: data <= 32'hb900ba6f;
    11'b00100000010: data <= 32'h2e9ebc03;
    11'b00100000011: data <= 32'h3d3c39cd;
    11'b00100000100: data <= 32'h3e084121;
    11'b00100000101: data <= 32'h39cc4076;
    11'b00100000110: data <= 32'h32623293;
    11'b00100000111: data <= 32'h3348bc05;
    11'b00100001000: data <= 32'ha1f7b7fb;
    11'b00100001001: data <= 32'hb8062406;
    11'b00100001010: data <= 32'hab7bbaa4;
    11'b00100001011: data <= 32'h3ddbbfba;
    11'b00100001100: data <= 32'h406bbe59;
    11'b00100001101: data <= 32'h3a76b109;
    11'b00100001110: data <= 32'hbd6e392a;
    11'b00100001111: data <= 32'hbf9535ad;
    11'b00100010000: data <= 32'hba54a4de;
    11'b00100010001: data <= 32'hb38baae9;
    11'b00100010010: data <= 32'hbca5b716;
    11'b00100010011: data <= 32'hbf77bcb3;
    11'b00100010100: data <= 32'hba48bb6b;
    11'b00100010101: data <= 32'h3c183a6f;
    11'b00100010110: data <= 32'h3de040ac;
    11'b00100010111: data <= 32'h36bc3fc4;
    11'b00100011000: data <= 32'hb7a2370b;
    11'b00100011001: data <= 32'hb6e426c0;
    11'b00100011010: data <= 32'hb21e3b51;
    11'b00100011011: data <= 32'hb1123c3b;
    11'b00100011100: data <= 32'h368fb855;
    11'b00100011101: data <= 32'h3eacc031;
    11'b00100011110: data <= 32'h4078be78;
    11'b00100011111: data <= 32'h3c9531cf;
    11'b00100100000: data <= 32'hb5d13c1f;
    11'b00100100001: data <= 32'hb83834d4;
    11'b00100100010: data <= 32'h3327b8f0;
    11'b00100100011: data <= 32'hac5cba9a;
    11'b00100100100: data <= 32'hbe8cbb92;
    11'b00100100101: data <= 32'hc0adbd84;
    11'b00100100110: data <= 32'hbad9bcf3;
    11'b00100100111: data <= 32'h3c8c239f;
    11'b00100101000: data <= 32'h3d023cdf;
    11'b00100101001: data <= 32'hb5313c86;
    11'b00100101010: data <= 32'hbda837b3;
    11'b00100101011: data <= 32'hbc423a98;
    11'b00100101100: data <= 32'hb6563f4b;
    11'b00100101101: data <= 32'hb4933e1c;
    11'b00100101110: data <= 32'ha9e6b721;
    11'b00100101111: data <= 32'h3b64bf6f;
    11'b00100110000: data <= 32'h3ef1bb4c;
    11'b00100110001: data <= 32'h3db83c6d;
    11'b00100110010: data <= 32'h39883e8c;
    11'b00100110011: data <= 32'h399735c6;
    11'b00100110100: data <= 32'h3bd9ba66;
    11'b00100110101: data <= 32'h3028ba46;
    11'b00100110110: data <= 32'hbe1fb8de;
    11'b00100110111: data <= 32'hbf83bcc1;
    11'b00100111000: data <= 32'hb064bedf;
    11'b00100111001: data <= 32'h3e5dbcb8;
    11'b00100111010: data <= 32'h3c67b09b;
    11'b00100111011: data <= 32'hbad83458;
    11'b00100111100: data <= 32'hbf323538;
    11'b00100111101: data <= 32'hbc5c3bcd;
    11'b00100111110: data <= 32'hb69a3f04;
    11'b00100111111: data <= 32'hba9a3ca9;
    11'b00101000000: data <= 32'hbce1b952;
    11'b00101000001: data <= 32'hb638be0f;
    11'b00101000010: data <= 32'h3bb9af10;
    11'b00101000011: data <= 32'h3ddd3f55;
    11'b00101000100: data <= 32'h3cbc3fb6;
    11'b00101000101: data <= 32'h3c4b3709;
    11'b00101000110: data <= 32'h3c16b635;
    11'b00101000111: data <= 32'h310431d8;
    11'b00101001000: data <= 32'hbc4a37f8;
    11'b00101001001: data <= 32'hbbbeb913;
    11'b00101001010: data <= 32'h3a07c011;
    11'b00101001011: data <= 32'h4002c015;
    11'b00101001100: data <= 32'h3c6ebb68;
    11'b00101001101: data <= 32'hb9dcaeba;
    11'b00101001110: data <= 32'hbcd4304a;
    11'b00101001111: data <= 32'hb4e23835;
    11'b00101010000: data <= 32'haf303b63;
    11'b00101010001: data <= 32'hbda03533;
    11'b00101010010: data <= 32'hc0cbbc1f;
    11'b00101010011: data <= 32'hbdebbd65;
    11'b00101010100: data <= 32'h36523049;
    11'b00101010101: data <= 32'h3d123ece;
    11'b00101010110: data <= 32'h3b2f3e15;
    11'b00101010111: data <= 32'h37c735c2;
    11'b00101011000: data <= 32'h368a3567;
    11'b00101011001: data <= 32'ha4913e19;
    11'b00101011010: data <= 32'hb9663eff;
    11'b00101011011: data <= 32'hb5f6a6d9;
    11'b00101011100: data <= 32'h3c31c000;
    11'b00101011101: data <= 32'h3fc0c028;
    11'b00101011110: data <= 32'h3ca8b9a6;
    11'b00101011111: data <= 32'ha7e3322e;
    11'b00101100000: data <= 32'h2d762c1b;
    11'b00101100001: data <= 32'h3b5fae3b;
    11'b00101100010: data <= 32'h36622c05;
    11'b00101100011: data <= 32'hbe98b431;
    11'b00101100100: data <= 32'hc1bbbcb2;
    11'b00101100101: data <= 32'hbecabdac;
    11'b00101100110: data <= 32'h3602b623;
    11'b00101100111: data <= 32'h3c0a394b;
    11'b00101101000: data <= 32'h30ab3804;
    11'b00101101001: data <= 32'hb8072981;
    11'b00101101010: data <= 32'hb4b93b05;
    11'b00101101011: data <= 32'hb21a40d8;
    11'b00101101100: data <= 32'hb8db40ca;
    11'b00101101101: data <= 32'hb8a63404;
    11'b00101101110: data <= 32'h363dbec2;
    11'b00101101111: data <= 32'h3cfcbd81;
    11'b00101110000: data <= 32'h3c5b3388;
    11'b00101110001: data <= 32'h39ff3acb;
    11'b00101110010: data <= 32'h3d2f2f0f;
    11'b00101110011: data <= 32'h3f87b6e8;
    11'b00101110100: data <= 32'h3a9eaf56;
    11'b00101110101: data <= 32'hbdbda455;
    11'b00101110110: data <= 32'hc0d3ba89;
    11'b00101110111: data <= 32'hbbfabe34;
    11'b00101111000: data <= 32'h3acdbd2e;
    11'b00101111001: data <= 32'h3ad3b971;
    11'b00101111010: data <= 32'hb7feb8aa;
    11'b00101111011: data <= 32'hbc4fb635;
    11'b00101111100: data <= 32'hb6b43b16;
    11'b00101111101: data <= 32'hacab40bb;
    11'b00101111110: data <= 32'hba9a402d;
    11'b00101111111: data <= 32'hbde329fa;
    11'b00110000000: data <= 32'hbb28bd5a;
    11'b00110000001: data <= 32'h3392b7d5;
    11'b00110000010: data <= 32'h3a7c3c7d;
    11'b00110000011: data <= 32'h3c433cf7;
    11'b00110000100: data <= 32'h3ebf2da6;
    11'b00110000101: data <= 32'h400ab4eb;
    11'b00110000110: data <= 32'h3b4f389f;
    11'b00110000111: data <= 32'hbbab3c34;
    11'b00110001000: data <= 32'hbdc4a59b;
    11'b00110001001: data <= 32'h2654be1c;
    11'b00110001010: data <= 32'h3d74bfce;
    11'b00110001011: data <= 32'h3a51bded;
    11'b00110001100: data <= 32'hb907bc68;
    11'b00110001101: data <= 32'hb9fbb988;
    11'b00110001110: data <= 32'h350d365d;
    11'b00110001111: data <= 32'h37533dfa;
    11'b00110010000: data <= 32'hbc373c98;
    11'b00110010001: data <= 32'hc0d8b693;
    11'b00110010010: data <= 32'hc003bc82;
    11'b00110010011: data <= 32'hb820a71f;
    11'b00110010100: data <= 32'h371f3cf5;
    11'b00110010101: data <= 32'h39b63b2d;
    11'b00110010110: data <= 32'h3c50b277;
    11'b00110010111: data <= 32'h3d632c5a;
    11'b00110011000: data <= 32'h394f3eb8;
    11'b00110011001: data <= 32'hb84740a5;
    11'b00110011010: data <= 32'hb94a3a68;
    11'b00110011011: data <= 32'h3871bd18;
    11'b00110011100: data <= 32'h3d82bf93;
    11'b00110011101: data <= 32'h394ebd07;
    11'b00110011110: data <= 32'hb440ba4e;
    11'b00110011111: data <= 32'h34c9b9bb;
    11'b00110100000: data <= 32'h3e3eb3bc;
    11'b00110100001: data <= 32'h3cd537ae;
    11'b00110100010: data <= 32'hbc223578;
    11'b00110100011: data <= 32'hc188b939;
    11'b00110100100: data <= 32'hc078bc2e;
    11'b00110100101: data <= 32'hb88fb32d;
    11'b00110100110: data <= 32'h32173734;
    11'b00110100111: data <= 32'hab32b03d;
    11'b00110101000: data <= 32'ha89dba2d;
    11'b00110101001: data <= 32'h371c3500;
    11'b00110101010: data <= 32'h361440dc;
    11'b00110101011: data <= 32'hb59941fc;
    11'b00110101100: data <= 32'hb8923ca7;
    11'b00110101101: data <= 32'h30ddbb55;
    11'b00110101110: data <= 32'h3983bca4;
    11'b00110101111: data <= 32'h3551b2f0;
    11'b00110110000: data <= 32'h324b28e0;
    11'b00110110001: data <= 32'h3d60b874;
    11'b00110110010: data <= 32'h411fb94c;
    11'b00110110011: data <= 32'h3f1527d2;
    11'b00110110100: data <= 32'hb9c73541;
    11'b00110110101: data <= 32'hc088b523;
    11'b00110110110: data <= 32'hbdd7bb78;
    11'b00110110111: data <= 32'h291fba6f;
    11'b00110111000: data <= 32'h3065b9ad;
    11'b00110111001: data <= 32'hba1ebd15;
    11'b00110111010: data <= 32'hbad7bd88;
    11'b00110111011: data <= 32'h2bf43188;
    11'b00110111100: data <= 32'h3726409e;
    11'b00110111101: data <= 32'hb5844147;
    11'b00110111110: data <= 32'hbc823aee;
    11'b00110111111: data <= 32'hbb7cb92f;
    11'b00111000000: data <= 32'hb60fb324;
    11'b00111000001: data <= 32'hb1463b1e;
    11'b00111000010: data <= 32'h3515397a;
    11'b00111000011: data <= 32'h3e9eb806;
    11'b00111000100: data <= 32'h415db9db;
    11'b00111000101: data <= 32'h3f41364b;
    11'b00111000110: data <= 32'hb4c33cbd;
    11'b00111000111: data <= 32'hbd003838;
    11'b00111001000: data <= 32'hb3bcb951;
    11'b00111001001: data <= 32'h3a62bce6;
    11'b00111001010: data <= 32'h3168bda9;
    11'b00111001011: data <= 32'hbc3cbf33;
    11'b00111001100: data <= 32'hbac0becc;
    11'b00111001101: data <= 32'h3890b4d6;
    11'b00111001110: data <= 32'h3c103d93;
    11'b00111001111: data <= 32'hb5133e1e;
    11'b00111010000: data <= 32'hbf3e31bb;
    11'b00111010001: data <= 32'hbfbeb85b;
    11'b00111010010: data <= 32'hbcaf3609;
    11'b00111010011: data <= 32'hb8d23d41;
    11'b00111010100: data <= 32'hac4438a4;
    11'b00111010101: data <= 32'h3c00ba7e;
    11'b00111010110: data <= 32'h3f78b8e4;
    11'b00111010111: data <= 32'h3d703cd4;
    11'b00111011000: data <= 32'h23fb40a9;
    11'b00111011001: data <= 32'hb5a83da5;
    11'b00111011010: data <= 32'h38acb48d;
    11'b00111011011: data <= 32'h3c43bc57;
    11'b00111011100: data <= 32'h2a64bc8f;
    11'b00111011101: data <= 32'hbb85bd88;
    11'b00111011110: data <= 32'hae45be3d;
    11'b00111011111: data <= 32'h3eb3bab8;
    11'b00111100000: data <= 32'h3f5e347f;
    11'b00111100001: data <= 32'haff7370b;
    11'b00111100010: data <= 32'hc00eb543;
    11'b00111100011: data <= 32'hc036b7f7;
    11'b00111100100: data <= 32'hbca3368c;
    11'b00111100101: data <= 32'hb9ef3aad;
    11'b00111100110: data <= 32'hba0bb4ac;
    11'b00111100111: data <= 32'hb25cbdd8;
    11'b00111101000: data <= 32'h399cb897;
    11'b00111101001: data <= 32'h3a6e3f2b;
    11'b00111101010: data <= 32'h306b41e0;
    11'b00111101011: data <= 32'hab023efe;
    11'b00111101100: data <= 32'h37f62326;
    11'b00111101101: data <= 32'h3872b670;
    11'b00111101110: data <= 32'hb5b2a654;
    11'b00111101111: data <= 32'hb9aab517;
    11'b00111110000: data <= 32'h39ffbc87;
    11'b00111110001: data <= 32'h4137bcb4;
    11'b00111110010: data <= 32'h40d4b5b5;
    11'b00111110011: data <= 32'h31f32eae;
    11'b00111110100: data <= 32'hbe29b26e;
    11'b00111110101: data <= 32'hbd0db53a;
    11'b00111110110: data <= 32'hb5782cb3;
    11'b00111110111: data <= 32'hb85cae77;
    11'b00111111000: data <= 32'hbd7abd6d;
    11'b00111111001: data <= 32'hbcbec03c;
    11'b00111111010: data <= 32'h9d36ba24;
    11'b00111111011: data <= 32'h391e3e96;
    11'b00111111100: data <= 32'h31ae4109;
    11'b00111111101: data <= 32'hb5d03d1d;
    11'b00111111110: data <= 32'hb5732c0e;
    11'b00111111111: data <= 32'hb6dc370d;
    11'b01000000000: data <= 32'hbb6a3cef;
    11'b01000000001: data <= 32'hb98b3931;
    11'b01000000010: data <= 32'h3c00ba97;
    11'b01000000011: data <= 32'h4158bd01;
    11'b01000000100: data <= 32'h40a8b391;
    11'b01000000101: data <= 32'h36e63983;
    11'b01000000110: data <= 32'hb8dc385d;
    11'b01000000111: data <= 32'h2e0f2816;
    11'b01000001000: data <= 32'h39d5b24a;
    11'b01000001001: data <= 32'hb3c8b9b5;
    11'b01000001010: data <= 32'hbe90bf5d;
    11'b01000001011: data <= 32'hbda1c0b4;
    11'b01000001100: data <= 32'h32cbbc73;
    11'b01000001101: data <= 32'h3c533a60;
    11'b01000001110: data <= 32'h34c13d20;
    11'b01000001111: data <= 32'hbae434ae;
    11'b01000010000: data <= 32'hbcdcaf0a;
    11'b01000010001: data <= 32'hbcbb3bfa;
    11'b01000010010: data <= 32'hbd533f86;
    11'b01000010011: data <= 32'hbc013ad4;
    11'b01000010100: data <= 32'h363cbbcd;
    11'b01000010101: data <= 32'h3efbbcd9;
    11'b01000010110: data <= 32'h3e6535ec;
    11'b01000010111: data <= 32'h378a3eb7;
    11'b01000011000: data <= 32'h33663d93;
    11'b01000011001: data <= 32'h3c8b36c8;
    11'b01000011010: data <= 32'h3d49acf2;
    11'b01000011011: data <= 32'hb193b74f;
    11'b01000011100: data <= 32'hbe59bd52;
    11'b01000011101: data <= 32'hbb10bfe2;
    11'b01000011110: data <= 32'h3c88bd92;
    11'b01000011111: data <= 32'h3f76b401;
    11'b01000100000: data <= 32'h384ba369;
    11'b01000100001: data <= 32'hbc2eb86f;
    11'b01000100010: data <= 32'hbd83b484;
    11'b01000100011: data <= 32'hbc643c4c;
    11'b01000100100: data <= 32'hbd183e87;
    11'b01000100101: data <= 32'hbdda3225;
    11'b01000100110: data <= 32'hb9f1be48;
    11'b01000100111: data <= 32'h361fbcfb;
    11'b01000101000: data <= 32'h39913b01;
    11'b01000101001: data <= 32'h358d4080;
    11'b01000101010: data <= 32'h386d3eb4;
    11'b01000101011: data <= 32'h3d26389d;
    11'b01000101100: data <= 32'h3c3536b9;
    11'b01000101101: data <= 32'hb80b38c9;
    11'b01000101110: data <= 32'hbdc2ad52;
    11'b01000101111: data <= 32'hb0d6bccc;
    11'b01000110000: data <= 32'h4003bdd9;
    11'b01000110001: data <= 32'h40cdbb1f;
    11'b01000110010: data <= 32'h3a06b8c1;
    11'b01000110011: data <= 32'hb992b999;
    11'b01000110100: data <= 32'hb8a8b2d9;
    11'b01000110101: data <= 32'haf793a9c;
    11'b01000110110: data <= 32'hba013abe;
    11'b01000110111: data <= 32'hbf36ba52;
    11'b01000111000: data <= 32'hbedcc068;
    11'b01000111001: data <= 32'hb891bd93;
    11'b01000111010: data <= 32'h333b3a90;
    11'b01000111011: data <= 32'h33f33f78;
    11'b01000111100: data <= 32'h353f3c43;
    11'b01000111101: data <= 32'h38fc3540;
    11'b01000111110: data <= 32'h31ae3bfa;
    11'b01000111111: data <= 32'hbc3e3f53;
    11'b01001000000: data <= 32'hbdaf3c86;
    11'b01001000001: data <= 32'h30a1b878;
    11'b01001000010: data <= 32'h402fbd72;
    11'b01001000011: data <= 32'h4066baba;
    11'b01001000100: data <= 32'h39e8b2a8;
    11'b01001000101: data <= 32'ha127ae1e;
    11'b01001000110: data <= 32'h39f8300a;
    11'b01001000111: data <= 32'h3ccb38b6;
    11'b01001001000: data <= 32'hae3a334f;
    11'b01001001001: data <= 32'hbf77bd24;
    11'b01001001010: data <= 32'hbff8c0b5;
    11'b01001001011: data <= 32'hb894be18;
    11'b01001001100: data <= 32'h37cc3219;
    11'b01001001101: data <= 32'h35583946;
    11'b01001001110: data <= 32'haf3bb107;
    11'b01001001111: data <= 32'hb2d5b28f;
    11'b01001010000: data <= 32'hb8983d49;
    11'b01001010001: data <= 32'hbda5410a;
    11'b01001010010: data <= 32'hbe423e4a;
    11'b01001010011: data <= 32'hb476b7d2;
    11'b01001010100: data <= 32'h3cc9bd0e;
    11'b01001010101: data <= 32'h3cffb4e0;
    11'b01001010110: data <= 32'h36be39a7;
    11'b01001010111: data <= 32'h38aa39da;
    11'b01001011000: data <= 32'h3f4737d8;
    11'b01001011001: data <= 32'h401738c5;
    11'b01001011010: data <= 32'h33723558;
    11'b01001011011: data <= 32'hbee2ba72;
    11'b01001011100: data <= 32'hbe2bbf1a;
    11'b01001011101: data <= 32'h33a9bdd9;
    11'b01001011110: data <= 32'h3ce7b8d9;
    11'b01001011111: data <= 32'h387eb94d;
    11'b01001100000: data <= 32'hb5c7bd18;
    11'b01001100001: data <= 32'hb7d1b968;
    11'b01001100010: data <= 32'hb82e3d18;
    11'b01001100011: data <= 32'hbcc340b1;
    11'b01001100100: data <= 32'hbedb3c34;
    11'b01001100101: data <= 32'hbca9bc09;
    11'b01001100110: data <= 32'hb1f0bd27;
    11'b01001100111: data <= 32'h2c3c333d;
    11'b01001101000: data <= 32'ha8633d6a;
    11'b01001101001: data <= 32'h39fd3c30;
    11'b01001101010: data <= 32'h40163821;
    11'b01001101011: data <= 32'h3fcb3a92;
    11'b01001101100: data <= 32'h22a53ca1;
    11'b01001101101: data <= 32'hbe3c373e;
    11'b01001101110: data <= 32'hba83b9ca;
    11'b01001101111: data <= 32'h3c9cbcb5;
    11'b01001110000: data <= 32'h3f2bbc3f;
    11'b01001110001: data <= 32'h397fbd43;
    11'b01001110010: data <= 32'hb39dbe81;
    11'b01001110011: data <= 32'h2e28ba18;
    11'b01001110100: data <= 32'h37603bfb;
    11'b01001110101: data <= 32'hb65f3e55;
    11'b01001110110: data <= 32'hbec22c00;
    11'b01001110111: data <= 32'hbfbabea9;
    11'b01001111000: data <= 32'hbcd8bd82;
    11'b01001111001: data <= 32'hb928359d;
    11'b01001111010: data <= 32'hb55d3c9f;
    11'b01001111011: data <= 32'h378e3717;
    11'b01001111100: data <= 32'h3db32567;
    11'b01001111101: data <= 32'h3c683c29;
    11'b01001111110: data <= 32'hb86a4058;
    11'b01001111111: data <= 32'hbe063ef1;
    11'b01010000000: data <= 32'hb61931fe;
    11'b01010000001: data <= 32'h3d9bba9c;
    11'b01010000010: data <= 32'h3e6ebb77;
    11'b01010000011: data <= 32'h3749bbe8;
    11'b01010000100: data <= 32'h2ef1bc5c;
    11'b01010000101: data <= 32'h3cd1b6f7;
    11'b01010000110: data <= 32'h3f5d39ef;
    11'b01010000111: data <= 32'h385d3af6;
    11'b01010001000: data <= 32'hbdd8b892;
    11'b01010001001: data <= 32'hc033bf61;
    11'b01010001010: data <= 32'hbd22bd4d;
    11'b01010001011: data <= 32'hb7ee2847;
    11'b01010001100: data <= 32'hb4c23140;
    11'b01010001101: data <= 32'h24eebab6;
    11'b01010001110: data <= 32'h3833ba81;
    11'b01010001111: data <= 32'h33933c2a;
    11'b01010010000: data <= 32'hbb8e4174;
    11'b01010010001: data <= 32'hbe074084;
    11'b01010010010: data <= 32'hb83336a0;
    11'b01010010011: data <= 32'h39b7b916;
    11'b01010010100: data <= 32'h38dab610;
    11'b01010010101: data <= 32'hb135a95c;
    11'b01010010110: data <= 32'h35c1b1c1;
    11'b01010010111: data <= 32'h403fa5ef;
    11'b01010011000: data <= 32'h418e3928;
    11'b01010011001: data <= 32'h3c4e39dc;
    11'b01010011010: data <= 32'hbcb3b4b4;
    11'b01010011011: data <= 32'hbe77bcec;
    11'b01010011100: data <= 32'hb774bbcb;
    11'b01010011101: data <= 32'h34a7b69e;
    11'b01010011110: data <= 32'ha6c6bbee;
    11'b01010011111: data <= 32'hb4d0c01c;
    11'b01010100000: data <= 32'h29babe1a;
    11'b01010100001: data <= 32'h2e0b3a72;
    11'b01010100010: data <= 32'hb9af40ff;
    11'b01010100011: data <= 32'hbd903f04;
    11'b01010100100: data <= 32'hbc42af42;
    11'b01010100101: data <= 32'hb7e0b980;
    11'b01010100110: data <= 32'hb9783272;
    11'b01010100111: data <= 32'hbb293a31;
    11'b01010101000: data <= 32'h34b23512;
    11'b01010101001: data <= 32'h408e22fc;
    11'b01010101010: data <= 32'h4172391a;
    11'b01010101011: data <= 32'h3b263ce3;
    11'b01010101100: data <= 32'hbc0e3a40;
    11'b01010101101: data <= 32'hbacfacb8;
    11'b01010101110: data <= 32'h38abb62e;
    11'b01010101111: data <= 32'h3c17b8ca;
    11'b01010110000: data <= 32'h3029be3b;
    11'b01010110001: data <= 32'hb5f3c0f3;
    11'b01010110010: data <= 32'h3514becb;
    11'b01010110011: data <= 32'h3b1d37e8;
    11'b01010110100: data <= 32'h31ae3ed0;
    11'b01010110101: data <= 32'hbc353946;
    11'b01010110110: data <= 32'hbe1fbb53;
    11'b01010110111: data <= 32'hbdaaba92;
    11'b01010111000: data <= 32'hbdf337bf;
    11'b01010111001: data <= 32'hbd593ae6;
    11'b01010111010: data <= 32'habb5adfc;
    11'b01010111011: data <= 32'h3e7fb879;
    11'b01010111100: data <= 32'h3f34385c;
    11'b01010111101: data <= 32'h32ad3fab;
    11'b01010111110: data <= 32'hbc0c3fcd;
    11'b01010111111: data <= 32'hb4a93b9e;
    11'b01011000000: data <= 32'h3c5f3111;
    11'b01011000001: data <= 32'h3c23b58b;
    11'b01011000010: data <= 32'hb0fcbcc5;
    11'b01011000011: data <= 32'hb522bf97;
    11'b01011000100: data <= 32'h3c65bd25;
    11'b01011000101: data <= 32'h40493494;
    11'b01011000110: data <= 32'h3d013b1d;
    11'b01011000111: data <= 32'hb8a9b2c0;
    11'b01011001000: data <= 32'hbe1dbd2d;
    11'b01011001001: data <= 32'hbdc6b9ee;
    11'b01011001010: data <= 32'hbd553705;
    11'b01011001011: data <= 32'hbd09323d;
    11'b01011001100: data <= 32'hb7b0bcf5;
    11'b01011001101: data <= 32'h3927be1d;
    11'b01011001110: data <= 32'h39cb3458;
    11'b01011001111: data <= 32'hb6214085;
    11'b01011010000: data <= 32'hbc0c40d6;
    11'b01011010001: data <= 32'hb2183cd9;
    11'b01011010010: data <= 32'h39cb35d2;
    11'b01011010011: data <= 32'h31c03278;
    11'b01011010100: data <= 32'hbb41b1bc;
    11'b01011010101: data <= 32'hb5deba71;
    11'b01011010110: data <= 32'h3f1bb973;
    11'b01011010111: data <= 32'h420a32cd;
    11'b01011011000: data <= 32'h3f66384b;
    11'b01011011001: data <= 32'hb32cb3d3;
    11'b01011011010: data <= 32'hbc0fbabb;
    11'b01011011011: data <= 32'hb88bb44d;
    11'b01011011100: data <= 32'hb66034c9;
    11'b01011011101: data <= 32'hba81b991;
    11'b01011011110: data <= 32'hba15c0c8;
    11'b01011011111: data <= 32'ha55dc0af;
    11'b01011100000: data <= 32'h3480adef;
    11'b01011100001: data <= 32'hb53e3fdb;
    11'b01011100010: data <= 32'hba5c3f72;
    11'b01011100011: data <= 32'hb6c43895;
    11'b01011100100: data <= 32'hb26d314f;
    11'b01011100101: data <= 32'hbc2839e6;
    11'b01011100110: data <= 32'hbf133a5a;
    11'b01011100111: data <= 32'hb8e7a560;
    11'b01011101000: data <= 32'h3f4bb72e;
    11'b01011101001: data <= 32'h41d4304d;
    11'b01011101010: data <= 32'h3e6339d6;
    11'b01011101011: data <= 32'hb15e3849;
    11'b01011101100: data <= 32'hb4963382;
    11'b01011101101: data <= 32'h38f1377f;
    11'b01011101110: data <= 32'h38d3356a;
    11'b01011101111: data <= 32'hb72ebc7b;
    11'b01011110000: data <= 32'hbaf8c189;
    11'b01011110001: data <= 32'ha6c8c0fa;
    11'b01011110010: data <= 32'h3a2db58d;
    11'b01011110011: data <= 32'h37653cc1;
    11'b01011110100: data <= 32'hb4c9392b;
    11'b01011110101: data <= 32'hb908b7a7;
    11'b01011110110: data <= 32'hbb9db1b9;
    11'b01011110111: data <= 32'hbf3d3c21;
    11'b01011111000: data <= 32'hc0773c8e;
    11'b01011111001: data <= 32'hbbb4afd4;
    11'b01011111010: data <= 32'h3cabbb36;
    11'b01011111011: data <= 32'h3f8eaef2;
    11'b01011111100: data <= 32'h39833c92;
    11'b01011111101: data <= 32'hb5f13e03;
    11'b01011111110: data <= 32'h34443ced;
    11'b01011111111: data <= 32'h3d733c54;
    11'b01100000000: data <= 32'h3b6b3927;
    11'b01100000001: data <= 32'hb8b9b9cf;
    11'b01100000010: data <= 32'hbba0c035;
    11'b01100000011: data <= 32'h3769bf8e;
    11'b01100000100: data <= 32'h3f34b5db;
    11'b01100000101: data <= 32'h3e063646;
    11'b01100000110: data <= 32'h3476b710;
    11'b01100000111: data <= 32'hb823bcae;
    11'b01100001000: data <= 32'hbb5fb444;
    11'b01100001001: data <= 32'hbe593c63;
    11'b01100001010: data <= 32'hc0053a1d;
    11'b01100001011: data <= 32'hbce4bc18;
    11'b01100001100: data <= 32'h32acbf56;
    11'b01100001101: data <= 32'h38e5b827;
    11'b01100001110: data <= 32'hb2e13d4e;
    11'b01100001111: data <= 32'hb87d3f8b;
    11'b01100010000: data <= 32'h373d3dc5;
    11'b01100010001: data <= 32'h3d213cc8;
    11'b01100010010: data <= 32'h35593c4b;
    11'b01100010011: data <= 32'hbd2b3450;
    11'b01100010100: data <= 32'hbc9cbaa2;
    11'b01100010101: data <= 32'h3b88bbd6;
    11'b01100010110: data <= 32'h4121b370;
    11'b01100010111: data <= 32'h4025a540;
    11'b01100011000: data <= 32'h38ccba11;
    11'b01100011001: data <= 32'hac9dbbfc;
    11'b01100011010: data <= 32'haaa6305b;
    11'b01100011011: data <= 32'hb7de3c77;
    11'b01100011100: data <= 32'hbd1e2e87;
    11'b01100011101: data <= 32'hbd26c014;
    11'b01100011110: data <= 32'hb7e8c143;
    11'b01100011111: data <= 32'haeedbb2f;
    11'b01100100000: data <= 32'hb75f3c2e;
    11'b01100100001: data <= 32'hb70e3d45;
    11'b01100100010: data <= 32'h35fd3957;
    11'b01100100011: data <= 32'h38de39f3;
    11'b01100100100: data <= 32'hb9d33d9a;
    11'b01100100101: data <= 32'hc04c3d0e;
    11'b01100100110: data <= 32'hbdd6331c;
    11'b01100100111: data <= 32'h3b9fb6d8;
    11'b01100101000: data <= 32'h40ddb1d6;
    11'b01100101001: data <= 32'h3ed727ef;
    11'b01100101010: data <= 32'h3717b3da;
    11'b01100101011: data <= 32'h3779ae87;
    11'b01100101100: data <= 32'h3c953afa;
    11'b01100101101: data <= 32'h3a1f3d06;
    11'b01100101110: data <= 32'hb8acb3af;
    11'b01100101111: data <= 32'hbcf5c0bf;
    11'b01100110000: data <= 32'hb8f8c164;
    11'b01100110001: data <= 32'h2e98bbe7;
    11'b01100110010: data <= 32'h2fcc36d5;
    11'b01100110011: data <= 32'h2a092dec;
    11'b01100110100: data <= 32'h34c3b8ff;
    11'b01100110101: data <= 32'ha4af2c35;
    11'b01100110110: data <= 32'hbdc33e0c;
    11'b01100110111: data <= 32'hc11f3ed6;
    11'b01100111000: data <= 32'hbecb3689;
    11'b01100111001: data <= 32'h36a9b924;
    11'b01100111010: data <= 32'h3d92b663;
    11'b01100111011: data <= 32'h38a234c1;
    11'b01100111100: data <= 32'had79387c;
    11'b01100111101: data <= 32'h3a963a93;
    11'b01100111110: data <= 32'h3fe53ddb;
    11'b01100111111: data <= 32'h3d873e07;
    11'b01101000000: data <= 32'hb7542cd1;
    11'b01101000001: data <= 32'hbd12bec6;
    11'b01101000010: data <= 32'hb48abf96;
    11'b01101000011: data <= 32'h3b83b99b;
    11'b01101000100: data <= 32'h3c4ab16a;
    11'b01101000101: data <= 32'h3902bc43;
    11'b01101000110: data <= 32'h368cbe73;
    11'b01101000111: data <= 32'ha5e9b517;
    11'b01101001000: data <= 32'hbccd3df8;
    11'b01101001001: data <= 32'hc0583dee;
    11'b01101001010: data <= 32'hbebcb467;
    11'b01101001011: data <= 32'hb596bdd5;
    11'b01101001100: data <= 32'h2ae9ba94;
    11'b01101001101: data <= 32'hb8fc36f4;
    11'b01101001110: data <= 32'hb8c43b79;
    11'b01101001111: data <= 32'h3b293c0d;
    11'b01101010000: data <= 32'h40113dcb;
    11'b01101010001: data <= 32'h3c1e3ed1;
    11'b01101010010: data <= 32'hbc0e3b26;
    11'b01101010011: data <= 32'hbdebb5d6;
    11'b01101010100: data <= 32'h2f2eb98b;
    11'b01101010101: data <= 32'h3e9db353;
    11'b01101010110: data <= 32'h3e77b710;
    11'b01101010111: data <= 32'h3addbe10;
    11'b01101011000: data <= 32'h3965bed1;
    11'b01101011001: data <= 32'h398eadf9;
    11'b01101011010: data <= 32'hab9f3e0f;
    11'b01101011011: data <= 32'hbca33b6b;
    11'b01101011100: data <= 32'hbd9cbcd3;
    11'b01101011101: data <= 32'hbb1fc073;
    11'b01101011110: data <= 32'hba55bc99;
    11'b01101011111: data <= 32'hbc9f3472;
    11'b01101100000: data <= 32'hb98637cb;
    11'b01101100001: data <= 32'h3a6a3261;
    11'b01101100010: data <= 32'h3def39ea;
    11'b01101100011: data <= 32'h2d5e3ec5;
    11'b01101100100: data <= 32'hbf513eda;
    11'b01101100101: data <= 32'hbf0f3a70;
    11'b01101100110: data <= 32'h32483152;
    11'b01101100111: data <= 32'h3e6f2cd9;
    11'b01101101000: data <= 32'h3ce2b59a;
    11'b01101101001: data <= 32'h37a1bc8d;
    11'b01101101010: data <= 32'h3b31bba8;
    11'b01101101011: data <= 32'h3edc38af;
    11'b01101101100: data <= 32'h3d3b3e9e;
    11'b01101101101: data <= 32'hb08d3877;
    11'b01101101110: data <= 32'hbc40be62;
    11'b01101101111: data <= 32'hbb97c088;
    11'b01101110000: data <= 32'hb9c9bc36;
    11'b01101110001: data <= 32'hba0eabb0;
    11'b01101110010: data <= 32'hb48db88d;
    11'b01101110011: data <= 32'h39eabcc7;
    11'b01101110100: data <= 32'h3af7b43f;
    11'b01101110101: data <= 32'hb93b3df0;
    11'b01101110110: data <= 32'hc075401f;
    11'b01101110111: data <= 32'hbf703c8d;
    11'b01101111000: data <= 32'hae753182;
    11'b01101111001: data <= 32'h39caa62a;
    11'b01101111010: data <= 32'h9a22ae5f;
    11'b01101111011: data <= 32'hb5fcb617;
    11'b01101111100: data <= 32'h3b5ba8dc;
    11'b01101111101: data <= 32'h40d93cb0;
    11'b01101111110: data <= 32'h40253f38;
    11'b01101111111: data <= 32'h33b03970;
    11'b01110000000: data <= 32'hbb76bc37;
    11'b01110000001: data <= 32'hb8efbd8a;
    11'b01110000010: data <= 32'h2893b752;
    11'b01110000011: data <= 32'h30f7b513;
    11'b01110000100: data <= 32'h34a3be62;
    11'b01110000101: data <= 32'h3a52c0ab;
    11'b01110000110: data <= 32'h39bfbb80;
    11'b01110000111: data <= 32'hb84a3d0e;
    11'b01110001000: data <= 32'hbf193f4a;
    11'b01110001001: data <= 32'hbe3f386c;
    11'b01110001010: data <= 32'hb849b88b;
    11'b01110001011: data <= 32'hb7a1b6ee;
    11'b01110001100: data <= 32'hbd702c3f;
    11'b01110001101: data <= 32'hbccd2e0c;
    11'b01110001110: data <= 32'h39fe341d;
    11'b01110001111: data <= 32'h40e73c73;
    11'b01110010000: data <= 32'h3f593f06;
    11'b01110010001: data <= 32'hb26c3cbf;
    11'b01110010010: data <= 32'hbc703050;
    11'b01110010011: data <= 32'hb2cba71b;
    11'b01110010100: data <= 32'h3a7b359f;
    11'b01110010101: data <= 32'h3a41b500;
    11'b01110010110: data <= 32'h3800bffa;
    11'b01110010111: data <= 32'h3ad2c11f;
    11'b01110011000: data <= 32'h3c9dbaf5;
    11'b01110011001: data <= 32'h37713ce2;
    11'b01110011010: data <= 32'hb8ed3d12;
    11'b01110011011: data <= 32'hbb79b66f;
    11'b01110011100: data <= 32'hba2fbd93;
    11'b01110011101: data <= 32'hbd05ba0a;
    11'b01110011110: data <= 32'hc0172c44;
    11'b01110011111: data <= 32'hbdfcaece;
    11'b01110100000: data <= 32'h3871b6b8;
    11'b01110100001: data <= 32'h3f9c3465;
    11'b01110100010: data <= 32'h3b323d9b;
    11'b01110100011: data <= 32'hbc323ebe;
    11'b01110100100: data <= 32'hbd993ce4;
    11'b01110100101: data <= 32'ha25b3c02;
    11'b01110100110: data <= 32'h3bc83b3a;
    11'b01110100111: data <= 32'h3825ad1f;
    11'b01110101000: data <= 32'h224ebe74;
    11'b01110101001: data <= 32'h3a08bf67;
    11'b01110101010: data <= 32'h3f66b20a;
    11'b01110101011: data <= 32'h3ef63d77;
    11'b01110101100: data <= 32'h38ad3a8a;
    11'b01110101101: data <= 32'hb4dcbbb4;
    11'b01110101110: data <= 32'hb92ebe3e;
    11'b01110101111: data <= 32'hbcb4b89e;
    11'b01110110000: data <= 32'hbede25b6;
    11'b01110110001: data <= 32'hbc82bac8;
    11'b01110110010: data <= 32'h37d8bedc;
    11'b01110110011: data <= 32'h3cf0bb5a;
    11'b01110110100: data <= 32'h25eb3af6;
    11'b01110110101: data <= 32'hbe443f3d;
    11'b01110110110: data <= 32'hbdc23e25;
    11'b01110110111: data <= 32'haaaf3c72;
    11'b01110111000: data <= 32'h362d3b1b;
    11'b01110111001: data <= 32'hb8d1322e;
    11'b01110111010: data <= 32'hbc19ba93;
    11'b01110111011: data <= 32'h36e7ba9d;
    11'b01110111100: data <= 32'h409b380f;
    11'b01110111101: data <= 32'h40f33df4;
    11'b01110111110: data <= 32'h3c6839c2;
    11'b01110111111: data <= 32'ha8aab996;
    11'b01111000000: data <= 32'hb42fba4e;
    11'b01111000001: data <= 32'hb657322f;
    11'b01111000010: data <= 32'hb9e12f52;
    11'b01111000011: data <= 32'hb758be63;
    11'b01111000100: data <= 32'h3847c1a2;
    11'b01111000101: data <= 32'h3b39bf05;
    11'b01111000110: data <= 32'haf5a3755;
    11'b01111000111: data <= 32'hbceb3dea;
    11'b01111001000: data <= 32'hbbe23b7f;
    11'b01111001001: data <= 32'hb095356e;
    11'b01111001010: data <= 32'hb8363694;
    11'b01111001011: data <= 32'hbfaa35a3;
    11'b01111001100: data <= 32'hc014b286;
    11'b01111001101: data <= 32'h2594b4cc;
    11'b01111001110: data <= 32'h4066389a;
    11'b01111001111: data <= 32'h40743d3e;
    11'b01111010000: data <= 32'h39573b30;
    11'b01111010001: data <= 32'hb3cf324e;
    11'b01111010010: data <= 32'h305b382d;
    11'b01111010011: data <= 32'h37d43cd6;
    11'b01111010100: data <= 32'h2e433666;
    11'b01111010101: data <= 32'haf4cbf52;
    11'b01111010110: data <= 32'h3804c211;
    11'b01111010111: data <= 32'h3c24beef;
    11'b01111011000: data <= 32'h38c1366c;
    11'b01111011001: data <= 32'hb0123b58;
    11'b01111011010: data <= 32'hb085aebd;
    11'b01111011011: data <= 32'hac47b94e;
    11'b01111011100: data <= 32'hbc6faa06;
    11'b01111011101: data <= 32'hc13136a5;
    11'b01111011110: data <= 32'hc0d9b04f;
    11'b01111011111: data <= 32'hb393b984;
    11'b01111100000: data <= 32'h3e7eb22c;
    11'b01111100001: data <= 32'h3ce239f4;
    11'b01111100010: data <= 32'hb53a3c40;
    11'b01111100011: data <= 32'hb94f3c43;
    11'b01111100100: data <= 32'h35f53e35;
    11'b01111100101: data <= 32'h3b1b3f94;
    11'b01111100110: data <= 32'h2f303a02;
    11'b01111100111: data <= 32'hb81cbd96;
    11'b01111101000: data <= 32'h329ec08a;
    11'b01111101001: data <= 32'h3d8fbb87;
    11'b01111101010: data <= 32'h3e84394a;
    11'b01111101011: data <= 32'h3c4c372f;
    11'b01111101100: data <= 32'h394cbafa;
    11'b01111101101: data <= 32'h336ebc63;
    11'b01111101110: data <= 32'hbb992653;
    11'b01111101111: data <= 32'hc0773855;
    11'b01111110000: data <= 32'hbff0b850;
    11'b01111110001: data <= 32'hb2d7beec;
    11'b01111110010: data <= 32'h3b91bd8a;
    11'b01111110011: data <= 32'h314d208a;
    11'b01111110100: data <= 32'hbc653bb5;
    11'b01111110101: data <= 32'hba9d3d13;
    11'b01111110110: data <= 32'h37933e93;
    11'b01111110111: data <= 32'h38fd3f6d;
    11'b01111111000: data <= 32'hb9f83bc9;
    11'b01111111001: data <= 32'hbe29b8c2;
    11'b01111111010: data <= 32'hb566bc5e;
    11'b01111111011: data <= 32'h3e509d7b;
    11'b01111111100: data <= 32'h40743b5b;
    11'b01111111101: data <= 32'h3e5e33af;
    11'b01111111110: data <= 32'h3baebb4a;
    11'b01111111111: data <= 32'h38eab8bc;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    