
module memory_rom_53(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3d7dba3e;
    11'b00000000001: data <= 32'h3a37b82d;
    11'b00000000010: data <= 32'hba3d36c1;
    11'b00000000011: data <= 32'hbf76304b;
    11'b00000000100: data <= 32'hbc28bd7c;
    11'b00000000101: data <= 32'h39b0c076;
    11'b00000000110: data <= 32'h3c38be3d;
    11'b00000000111: data <= 32'hb561b6bf;
    11'b00000001000: data <= 32'hbd57324b;
    11'b00000001001: data <= 32'hb90739ac;
    11'b00000001010: data <= 32'h352a3df4;
    11'b00000001011: data <= 32'hb5333e81;
    11'b00000001100: data <= 32'hbf6236e9;
    11'b00000001101: data <= 32'hbfffbaf2;
    11'b00000001110: data <= 32'hb583b877;
    11'b00000001111: data <= 32'h3d323b37;
    11'b00000010000: data <= 32'h3e7a3d8c;
    11'b00000010001: data <= 32'h3d17351c;
    11'b00000010010: data <= 32'h3c9db6bf;
    11'b00000010011: data <= 32'h3ace37fd;
    11'b00000010100: data <= 32'haf493e85;
    11'b00000010101: data <= 32'hba883ab9;
    11'b00000010110: data <= 32'hb218bda6;
    11'b00000010111: data <= 32'h3bc7c155;
    11'b00000011000: data <= 32'h3ba1bf98;
    11'b00000011001: data <= 32'hb201b88b;
    11'b00000011010: data <= 32'hb8d3ae25;
    11'b00000011011: data <= 32'h3577aabd;
    11'b00000011100: data <= 32'h3aa2363c;
    11'b00000011101: data <= 32'hb92139cc;
    11'b00000011110: data <= 32'hc15a30fe;
    11'b00000011111: data <= 32'hc180b91a;
    11'b00000100000: data <= 32'hba26b638;
    11'b00000100001: data <= 32'h3b7038a9;
    11'b00000100010: data <= 32'h3b6b3a1e;
    11'b00000100011: data <= 32'h34bf296b;
    11'b00000100100: data <= 32'h36072e30;
    11'b00000100101: data <= 32'h39cf3e69;
    11'b00000100110: data <= 32'h35b9415a;
    11'b00000100111: data <= 32'hb4873dac;
    11'b00000101000: data <= 32'had71bc82;
    11'b00000101001: data <= 32'h39a1c079;
    11'b00000101010: data <= 32'h3af4bcde;
    11'b00000101011: data <= 32'h3686a939;
    11'b00000101100: data <= 32'h389eb28c;
    11'b00000101101: data <= 32'h3df7ba73;
    11'b00000101110: data <= 32'h3dabb7d3;
    11'b00000101111: data <= 32'hb88a3458;
    11'b00000110000: data <= 32'hc14d31a4;
    11'b00000110001: data <= 32'hc0ffb90d;
    11'b00000110010: data <= 32'hb876bb4e;
    11'b00000110011: data <= 32'h38d7b79d;
    11'b00000110100: data <= 32'ha8efb480;
    11'b00000110101: data <= 32'hbaa8b699;
    11'b00000110110: data <= 32'hb4bd34d2;
    11'b00000110111: data <= 32'h3945400b;
    11'b00000111000: data <= 32'h374541cb;
    11'b00000111001: data <= 32'hb8a33e1b;
    11'b00000111010: data <= 32'hbaf4b967;
    11'b00000111011: data <= 32'hadeabce2;
    11'b00000111100: data <= 32'h392ca340;
    11'b00000111101: data <= 32'h3b323992;
    11'b00000111110: data <= 32'h3d85b26e;
    11'b00000111111: data <= 32'h4036bc99;
    11'b00001000000: data <= 32'h3f14b874;
    11'b00001000001: data <= 32'haef73986;
    11'b00001000010: data <= 32'hbf1e396b;
    11'b00001000011: data <= 32'hbdc1b928;
    11'b00001000100: data <= 32'h2cf6be8a;
    11'b00001000101: data <= 32'h3719be22;
    11'b00001000110: data <= 32'hb9a6bc83;
    11'b00001000111: data <= 32'hbd54bada;
    11'b00001001000: data <= 32'hb44ba6da;
    11'b00001001001: data <= 32'h3b473dd4;
    11'b00001001010: data <= 32'h34f34054;
    11'b00001001011: data <= 32'hbd963c8d;
    11'b00001001100: data <= 32'hc00ab4d4;
    11'b00001001101: data <= 32'hbbe2b422;
    11'b00001001110: data <= 32'h34953aff;
    11'b00001001111: data <= 32'h3ab23c0b;
    11'b00001010000: data <= 32'h3ce2b4c7;
    11'b00001010001: data <= 32'h3f2ebc27;
    11'b00001010010: data <= 32'h3ec73116;
    11'b00001010011: data <= 32'h37733f07;
    11'b00001010100: data <= 32'hb90c3dde;
    11'b00001010101: data <= 32'hb506b7f4;
    11'b00001010110: data <= 32'h38cebfb9;
    11'b00001010111: data <= 32'h3608bf43;
    11'b00001011000: data <= 32'hba4bbce3;
    11'b00001011001: data <= 32'hbb4ebc35;
    11'b00001011010: data <= 32'h3858b9c1;
    11'b00001011011: data <= 32'h3e02345e;
    11'b00001011100: data <= 32'h32d33c06;
    11'b00001011101: data <= 32'hc01938c4;
    11'b00001011110: data <= 32'hc16bb035;
    11'b00001011111: data <= 32'hbd972fbb;
    11'b00001100000: data <= 32'ha9a93afd;
    11'b00001100001: data <= 32'h31d5388c;
    11'b00001100010: data <= 32'h3164b93c;
    11'b00001100011: data <= 32'h3a4cba14;
    11'b00001100100: data <= 32'h3d3e3c38;
    11'b00001100101: data <= 32'h3adc4179;
    11'b00001100110: data <= 32'h2ddf4024;
    11'b00001100111: data <= 32'h2f4db22e;
    11'b00001101000: data <= 32'h384abe00;
    11'b00001101001: data <= 32'h3363bc42;
    11'b00001101010: data <= 32'hb712b7f5;
    11'b00001101011: data <= 32'h2873bb60;
    11'b00001101100: data <= 32'h3e7abd88;
    11'b00001101101: data <= 32'h404cba33;
    11'b00001101110: data <= 32'h35c73355;
    11'b00001101111: data <= 32'hbff23629;
    11'b00001110000: data <= 32'hc0caadb1;
    11'b00001110001: data <= 32'hbc1cb0d0;
    11'b00001110010: data <= 32'hb13d2c85;
    11'b00001110011: data <= 32'hb994b64c;
    11'b00001110100: data <= 32'hbc73bcc5;
    11'b00001110101: data <= 32'hb292b96d;
    11'b00001110110: data <= 32'h3bea3d9c;
    11'b00001110111: data <= 32'h3bb041cd;
    11'b00001111000: data <= 32'h296d4021;
    11'b00001111001: data <= 32'hb6482e3c;
    11'b00001111010: data <= 32'hb108b875;
    11'b00001111011: data <= 32'hadba346f;
    11'b00001111100: data <= 32'haf593865;
    11'b00001111101: data <= 32'h39deb934;
    11'b00001111110: data <= 32'h4061bed3;
    11'b00001111111: data <= 32'h40ddbc52;
    11'b00010000000: data <= 32'h39aa35a0;
    11'b00010000001: data <= 32'hbcad3a0e;
    11'b00010000010: data <= 32'hbcd59b7e;
    11'b00010000011: data <= 32'hae6db967;
    11'b00010000100: data <= 32'haaedbad1;
    11'b00010000101: data <= 32'hbd4cbcd0;
    11'b00010000110: data <= 32'hbf5cbe79;
    11'b00010000111: data <= 32'hb7dcbb98;
    11'b00010001000: data <= 32'h3c523af3;
    11'b00010001001: data <= 32'h3b38401e;
    11'b00010001010: data <= 32'hb8733da2;
    11'b00010001011: data <= 32'hbd8432a4;
    11'b00010001100: data <= 32'hbc0f35a2;
    11'b00010001101: data <= 32'hb79a3d89;
    11'b00010001110: data <= 32'hb1a03cc5;
    11'b00010001111: data <= 32'h38a7b874;
    11'b00010010000: data <= 32'h3f25bea6;
    11'b00010010001: data <= 32'h4041b8c2;
    11'b00010010010: data <= 32'h3c273ce6;
    11'b00010010011: data <= 32'had0d3e06;
    11'b00010010100: data <= 32'h300c3286;
    11'b00010010101: data <= 32'h3a1abb5d;
    11'b00010010110: data <= 32'h2e63bc77;
    11'b00010010111: data <= 32'hbdcdbce8;
    11'b00010011000: data <= 32'hbea2be85;
    11'b00010011001: data <= 32'h2e6bbdb7;
    11'b00010011010: data <= 32'h3e77b421;
    11'b00010011011: data <= 32'h3b1b399c;
    11'b00010011100: data <= 32'hbc75382b;
    11'b00010011101: data <= 32'hc00c303a;
    11'b00010011110: data <= 32'hbd833a0d;
    11'b00010011111: data <= 32'hb9673e81;
    11'b00010100000: data <= 32'hb94a3bfe;
    11'b00010100001: data <= 32'hb6b7baad;
    11'b00010100010: data <= 32'h38c5bde8;
    11'b00010100011: data <= 32'h3d9e3176;
    11'b00010100100: data <= 32'h3cab4045;
    11'b00010100101: data <= 32'h39334027;
    11'b00010100110: data <= 32'h3a7036e0;
    11'b00010100111: data <= 32'h3bd5b8e2;
    11'b00010101000: data <= 32'h2bb8b67a;
    11'b00010101001: data <= 32'hbcccb574;
    11'b00010101010: data <= 32'hbaf5bcb8;
    11'b00010101011: data <= 32'h3c55bf4e;
    11'b00010101100: data <= 32'h407cbd30;
    11'b00010101101: data <= 32'h3c05b546;
    11'b00010101110: data <= 32'hbc7e96cf;
    11'b00010101111: data <= 32'hbef12848;
    11'b00010110000: data <= 32'hbaf83895;
    11'b00010110001: data <= 32'hb80e3c09;
    11'b00010110010: data <= 32'hbd223101;
    11'b00010110011: data <= 32'hbebabd6f;
    11'b00010110100: data <= 32'hb930bd9f;
    11'b00010110101: data <= 32'h39f5385d;
    11'b00010110110: data <= 32'h3c5f40a0;
    11'b00010110111: data <= 32'h39683fd7;
    11'b00010111000: data <= 32'h380e3794;
    11'b00010111001: data <= 32'h37022e32;
    11'b00010111010: data <= 32'hb3b63b50;
    11'b00010111011: data <= 32'hbb543b9f;
    11'b00010111100: data <= 32'hb1ebb86e;
    11'b00010111101: data <= 32'h3ea0bfc2;
    11'b00010111110: data <= 32'h40e5bea6;
    11'b00010111111: data <= 32'h3c9cb6fe;
    11'b00011000000: data <= 32'hb81731bd;
    11'b00011000001: data <= 32'hb8922d51;
    11'b00011000010: data <= 32'h34b02f55;
    11'b00011000011: data <= 32'ha8d83070;
    11'b00011000100: data <= 32'hbeb7b924;
    11'b00011000101: data <= 32'hc0e9bef0;
    11'b00011000110: data <= 32'hbcbbbe1c;
    11'b00011000111: data <= 32'h38d431e0;
    11'b00011001000: data <= 32'h3bc63df9;
    11'b00011001001: data <= 32'h31013c57;
    11'b00011001010: data <= 32'hb63e3367;
    11'b00011001011: data <= 32'hb6423a1c;
    11'b00011001100: data <= 32'hb8d3401d;
    11'b00011001101: data <= 32'hbb093f70;
    11'b00011001110: data <= 32'hb270b207;
    11'b00011001111: data <= 32'h3d1cbf33;
    11'b00011010000: data <= 32'h3fccbd09;
    11'b00011010001: data <= 32'h3c993505;
    11'b00011010010: data <= 32'h355d3afd;
    11'b00011010011: data <= 32'h3a5a3482;
    11'b00011010100: data <= 32'h3dbbb1cb;
    11'b00011010101: data <= 32'h36c6b324;
    11'b00011010110: data <= 32'hbeb5b98e;
    11'b00011010111: data <= 32'hc0b5be5a;
    11'b00011011000: data <= 32'hb9f6bed2;
    11'b00011011001: data <= 32'h3c36b9a7;
    11'b00011011010: data <= 32'h3b9c2f19;
    11'b00011011011: data <= 32'hb6a0ad97;
    11'b00011011100: data <= 32'hbc62b1cb;
    11'b00011011101: data <= 32'hba413c0a;
    11'b00011011110: data <= 32'hb97640c2;
    11'b00011011111: data <= 32'hbc6b3f68;
    11'b00011100000: data <= 32'hbbd9b578;
    11'b00011100001: data <= 32'h2c78be65;
    11'b00011100010: data <= 32'h3b89b812;
    11'b00011100011: data <= 32'h3b603cff;
    11'b00011100100: data <= 32'h3b0b3de0;
    11'b00011100101: data <= 32'h3e3536c8;
    11'b00011100110: data <= 32'h3f7aad59;
    11'b00011100111: data <= 32'h3868349b;
    11'b00011101000: data <= 32'hbd933265;
    11'b00011101001: data <= 32'hbe69baf1;
    11'b00011101010: data <= 32'h3358bef4;
    11'b00011101011: data <= 32'h3ec7be2b;
    11'b00011101100: data <= 32'h3c0fbbfd;
    11'b00011101101: data <= 32'hb8b5bae9;
    11'b00011101110: data <= 32'hbbdab7e6;
    11'b00011101111: data <= 32'hb4723a2c;
    11'b00011110000: data <= 32'hb4503f43;
    11'b00011110001: data <= 32'hbd7d3c36;
    11'b00011110010: data <= 32'hc00fbaec;
    11'b00011110011: data <= 32'hbd01bdfd;
    11'b00011110100: data <= 32'h1408a1ca;
    11'b00011110101: data <= 32'h38b23e4f;
    11'b00011110110: data <= 32'h3a983d77;
    11'b00011110111: data <= 32'h3d4a3419;
    11'b00011111000: data <= 32'h3da534a8;
    11'b00011111001: data <= 32'h34623d92;
    11'b00011111010: data <= 32'hbc603e42;
    11'b00011111011: data <= 32'hbaa82b79;
    11'b00011111100: data <= 32'h3b6cbe35;
    11'b00011111101: data <= 32'h3fb4bf30;
    11'b00011111110: data <= 32'h3be7bcbf;
    11'b00011111111: data <= 32'hb477ba7c;
    11'b00100000000: data <= 32'ha6d8b807;
    11'b00100000001: data <= 32'h3b9b34d2;
    11'b00100000010: data <= 32'h380d3b27;
    11'b00100000011: data <= 32'hbdc130ed;
    11'b00100000100: data <= 32'hc156bd1e;
    11'b00100000101: data <= 32'hbf81bdef;
    11'b00100000110: data <= 32'hb504aeb5;
    11'b00100000111: data <= 32'h35c63ba9;
    11'b00100001000: data <= 32'h349536ff;
    11'b00100001001: data <= 32'h3677b4a2;
    11'b00100001010: data <= 32'h381938e8;
    11'b00100001011: data <= 32'hb02d40c4;
    11'b00100001100: data <= 32'hbbab4125;
    11'b00100001101: data <= 32'hb8ef3920;
    11'b00100001110: data <= 32'h39efbd08;
    11'b00100001111: data <= 32'h3d8fbd71;
    11'b00100010000: data <= 32'h3991b712;
    11'b00100010001: data <= 32'h3305ad4c;
    11'b00100010010: data <= 32'h3cb3b44b;
    11'b00100010011: data <= 32'h4066abd7;
    11'b00100010100: data <= 32'h3ce53568;
    11'b00100010101: data <= 32'hbcf1ad3c;
    11'b00100010110: data <= 32'hc107bc77;
    11'b00100010111: data <= 32'hbde0bd98;
    11'b00100011000: data <= 32'h3013b939;
    11'b00100011001: data <= 32'h35bcb410;
    11'b00100011010: data <= 32'hb544bacb;
    11'b00100011011: data <= 32'hb75abbeb;
    11'b00100011100: data <= 32'haa7638ef;
    11'b00100011101: data <= 32'hb3024145;
    11'b00100011110: data <= 32'hbba5413c;
    11'b00100011111: data <= 32'hbc463857;
    11'b00100100000: data <= 32'hb49dbc2f;
    11'b00100100001: data <= 32'h3452b89b;
    11'b00100100010: data <= 32'h310938f1;
    11'b00100100011: data <= 32'h37c83958;
    11'b00100100100: data <= 32'h3f63ae31;
    11'b00100100101: data <= 32'h416eb0e4;
    11'b00100100110: data <= 32'h3dd4385a;
    11'b00100100111: data <= 32'hbb3c3908;
    11'b00100101000: data <= 32'hbeebb4be;
    11'b00100101001: data <= 32'hb669bc72;
    11'b00100101010: data <= 32'h3b38bcbc;
    11'b00100101011: data <= 32'h3770bd0f;
    11'b00100101100: data <= 32'hb93ebeec;
    11'b00100101101: data <= 32'hb8fcbdd8;
    11'b00100101110: data <= 32'h343f349b;
    11'b00100101111: data <= 32'h34634012;
    11'b00100110000: data <= 32'hbb473f07;
    11'b00100110001: data <= 32'hbf2fad8b;
    11'b00100110010: data <= 32'hbdffbbec;
    11'b00100110011: data <= 32'hba602980;
    11'b00100110100: data <= 32'hb6353cc9;
    11'b00100110101: data <= 32'h34b83a0d;
    11'b00100110110: data <= 32'h3e50b51c;
    11'b00100110111: data <= 32'h4075acb2;
    11'b00100111000: data <= 32'h3c713d4a;
    11'b00100111001: data <= 32'hb9273f7c;
    11'b00100111010: data <= 32'hbae63a28;
    11'b00100111011: data <= 32'h3830b95b;
    11'b00100111100: data <= 32'h3d4dbd09;
    11'b00100111101: data <= 32'h368cbda2;
    11'b00100111110: data <= 32'hb8ecbebe;
    11'b00100111111: data <= 32'h20b6bdcc;
    11'b00101000000: data <= 32'h3d72b11b;
    11'b00101000001: data <= 32'h3cc63c24;
    11'b00101000010: data <= 32'hb9813940;
    11'b00101000011: data <= 32'hc06eb987;
    11'b00101000100: data <= 32'hc025bbca;
    11'b00101000101: data <= 32'hbca33210;
    11'b00101000110: data <= 32'hb92d3b22;
    11'b00101000111: data <= 32'hb3f3a756;
    11'b00101001000: data <= 32'h38c4bc03;
    11'b00101001001: data <= 32'h3ca1ab47;
    11'b00101001010: data <= 32'h38304021;
    11'b00101001011: data <= 32'hb83c41a4;
    11'b00101001100: data <= 32'hb6fb3dbe;
    11'b00101001101: data <= 32'h3925b48d;
    11'b00101001110: data <= 32'h3b94ba3d;
    11'b00101001111: data <= 32'h9eafb8de;
    11'b00101010000: data <= 32'hb6deba92;
    11'b00101010001: data <= 32'h3b88bc33;
    11'b00101010010: data <= 32'h4118b7c7;
    11'b00101010011: data <= 32'h400d34c6;
    11'b00101010100: data <= 32'hb5673005;
    11'b00101010101: data <= 32'hbfecb9a1;
    11'b00101010110: data <= 32'hbe76ba4d;
    11'b00101010111: data <= 32'hb8f8aa59;
    11'b00101011000: data <= 32'hb825a89c;
    11'b00101011001: data <= 32'hba99bcfc;
    11'b00101011010: data <= 32'hb6c1bf61;
    11'b00101011011: data <= 32'h3504b402;
    11'b00101011100: data <= 32'h33c84064;
    11'b00101011101: data <= 32'hb74641a5;
    11'b00101011110: data <= 32'hb8bb3d22;
    11'b00101011111: data <= 32'hade6b124;
    11'b00101100000: data <= 32'hadfea694;
    11'b00101100001: data <= 32'hb9a138ac;
    11'b00101100010: data <= 32'hb6683222;
    11'b00101100011: data <= 32'h3dd8b967;
    11'b00101100100: data <= 32'h420cb8f2;
    11'b00101100101: data <= 32'h40803341;
    11'b00101100110: data <= 32'ha9be3843;
    11'b00101100111: data <= 32'hbcd4255b;
    11'b00101101000: data <= 32'hb6e6b564;
    11'b00101101001: data <= 32'h364ab4f8;
    11'b00101101010: data <= 32'hb29fbaed;
    11'b00101101011: data <= 32'hbca8c032;
    11'b00101101100: data <= 32'hbabbc0b5;
    11'b00101101101: data <= 32'h3521b8c3;
    11'b00101101110: data <= 32'h38f13e57;
    11'b00101101111: data <= 32'hb40b3f71;
    11'b00101110000: data <= 32'hbc1d3719;
    11'b00101110001: data <= 32'hbc62b4cf;
    11'b00101110010: data <= 32'hbc8c38b6;
    11'b00101110011: data <= 32'hbd553d96;
    11'b00101110100: data <= 32'hb95138ba;
    11'b00101110101: data <= 32'h3c9eba09;
    11'b00101110110: data <= 32'h40e8b966;
    11'b00101110111: data <= 32'h3eec39a7;
    11'b00101111000: data <= 32'h29183e2f;
    11'b00101111001: data <= 32'hb5a53c3f;
    11'b00101111010: data <= 32'h39aa334f;
    11'b00101111011: data <= 32'h3c81b421;
    11'b00101111100: data <= 32'hae1abb8c;
    11'b00101111101: data <= 32'hbcf1bff6;
    11'b00101111110: data <= 32'hb80cc06d;
    11'b00101111111: data <= 32'h3cabbb30;
    11'b00110000000: data <= 32'h3e0438cc;
    11'b00110000001: data <= 32'h2f9b387f;
    11'b00110000010: data <= 32'hbd16b77c;
    11'b00110000011: data <= 32'hbe4eb78c;
    11'b00110000100: data <= 32'hbdd33a91;
    11'b00110000101: data <= 32'hbe113d88;
    11'b00110000110: data <= 32'hbc6c2c98;
    11'b00110000111: data <= 32'h31cdbd8e;
    11'b00110001000: data <= 32'h3cd1ba93;
    11'b00110001001: data <= 32'h3ac63cf1;
    11'b00110001010: data <= 32'haa1f40c0;
    11'b00110001011: data <= 32'h304e3ed1;
    11'b00110001100: data <= 32'h3c7338bf;
    11'b00110001101: data <= 32'h3c20316d;
    11'b00110001110: data <= 32'hb70eb089;
    11'b00110001111: data <= 32'hbcdcbbc2;
    11'b00110010000: data <= 32'h31f6be28;
    11'b00110010001: data <= 32'h406cbc12;
    11'b00110010010: data <= 32'h40a7b1b6;
    11'b00110010011: data <= 32'h3803b3e2;
    11'b00110010100: data <= 32'hbc23ba43;
    11'b00110010101: data <= 32'hbc68b61e;
    11'b00110010110: data <= 32'hba4e39ec;
    11'b00110010111: data <= 32'hbc9539b7;
    11'b00110011000: data <= 32'hbdeebbde;
    11'b00110011001: data <= 32'hbae6c076;
    11'b00110011010: data <= 32'h2decbc5f;
    11'b00110011011: data <= 32'h33e63d41;
    11'b00110011100: data <= 32'hae7240af;
    11'b00110011101: data <= 32'h2fe83dcb;
    11'b00110011110: data <= 32'h39353829;
    11'b00110011111: data <= 32'h31a539fa;
    11'b00110100000: data <= 32'hbc8f3c45;
    11'b00110100001: data <= 32'hbd3334c7;
    11'b00110100010: data <= 32'h38dbbaad;
    11'b00110100011: data <= 32'h4147bbf0;
    11'b00110100100: data <= 32'h40f4b600;
    11'b00110100101: data <= 32'h392eaffa;
    11'b00110100110: data <= 32'hb676b454;
    11'b00110100111: data <= 32'h2e4d2bf2;
    11'b00110101000: data <= 32'h376f38f5;
    11'b00110101001: data <= 32'hb80b25d9;
    11'b00110101010: data <= 32'hbe91bf15;
    11'b00110101011: data <= 32'hbd8ac165;
    11'b00110101100: data <= 32'hb232bd62;
    11'b00110101101: data <= 32'h360e3a72;
    11'b00110101110: data <= 32'h2cd93d72;
    11'b00110101111: data <= 32'hb1083642;
    11'b00110110000: data <= 32'hb1bd2bf5;
    11'b00110110001: data <= 32'hba4d3cad;
    11'b00110110010: data <= 32'hbf053fdd;
    11'b00110110011: data <= 32'hbe1b3bf7;
    11'b00110110100: data <= 32'h35c9b91e;
    11'b00110110101: data <= 32'h4018bbf6;
    11'b00110110110: data <= 32'h3f0fab0a;
    11'b00110110111: data <= 32'h36ff397b;
    11'b00110111000: data <= 32'h341f3960;
    11'b00110111001: data <= 32'h3d3f3914;
    11'b00110111010: data <= 32'h3dfe3981;
    11'b00110111011: data <= 32'hadf2acb6;
    11'b00110111100: data <= 32'hbe83be8f;
    11'b00110111101: data <= 32'hbcd1c0cb;
    11'b00110111110: data <= 32'h36c9bd8c;
    11'b00110111111: data <= 32'h3c901a04;
    11'b00111000000: data <= 32'h377298ca;
    11'b00111000001: data <= 32'hb56eba90;
    11'b00111000010: data <= 32'hb916b6e8;
    11'b00111000011: data <= 32'hbc563d25;
    11'b00111000100: data <= 32'hbf474032;
    11'b00111000101: data <= 32'hbf0239d3;
    11'b00111000110: data <= 32'hb726bc7c;
    11'b00111000111: data <= 32'h39e7bca1;
    11'b00111001000: data <= 32'h38b1360b;
    11'b00111001001: data <= 32'h22713dce;
    11'b00111001010: data <= 32'h38d83d26;
    11'b00111001011: data <= 32'h3f6a3b5f;
    11'b00111001100: data <= 32'h3eb43b9f;
    11'b00111001101: data <= 32'hb40938b7;
    11'b00111001110: data <= 32'hbe71b88c;
    11'b00111001111: data <= 32'hb90cbdc5;
    11'b00111010000: data <= 32'h3d7abcaa;
    11'b00111010001: data <= 32'h3fb7b8f0;
    11'b00111010010: data <= 32'h3a73bb88;
    11'b00111010011: data <= 32'hb2b0bdb8;
    11'b00111010100: data <= 32'hb44bb885;
    11'b00111010101: data <= 32'hb5f83cc2;
    11'b00111010110: data <= 32'hbcc83e41;
    11'b00111010111: data <= 32'hbf32b24e;
    11'b00111011000: data <= 32'hbd49bfaa;
    11'b00111011001: data <= 32'hb7f8bdaa;
    11'b00111011010: data <= 32'hb53d3817;
    11'b00111011011: data <= 32'hb4d23df7;
    11'b00111011100: data <= 32'h386f3bfd;
    11'b00111011101: data <= 32'h3e25390c;
    11'b00111011110: data <= 32'h3bdc3ce7;
    11'b00111011111: data <= 32'hbb183e84;
    11'b00111100000: data <= 32'hbed03a86;
    11'b00111100001: data <= 32'hb266b693;
    11'b00111100010: data <= 32'h3f59bac0;
    11'b00111100011: data <= 32'h401cb9f8;
    11'b00111100100: data <= 32'h3a35bbc4;
    11'b00111100101: data <= 32'h30f1bc74;
    11'b00111100110: data <= 32'h3a2bb2bd;
    11'b00111100111: data <= 32'h3be43c5a;
    11'b00111101000: data <= 32'hb32d3b33;
    11'b00111101001: data <= 32'hbe8abbf7;
    11'b00111101010: data <= 32'hbf00c0bc;
    11'b00111101011: data <= 32'hbb84be24;
    11'b00111101100: data <= 32'hb6dc3342;
    11'b00111101101: data <= 32'hb3ff393e;
    11'b00111101110: data <= 32'h34aab0ff;
    11'b00111101111: data <= 32'h3a22b0c7;
    11'b00111110000: data <= 32'h28b33d40;
    11'b00111110001: data <= 32'hbdf940d3;
    11'b00111110010: data <= 32'hbf5b3eae;
    11'b00111110011: data <= 32'hb4492aab;
    11'b00111110100: data <= 32'h3d7eb970;
    11'b00111110101: data <= 32'h3d09b6ee;
    11'b00111110110: data <= 32'h342fb3fc;
    11'b00111110111: data <= 32'h37b2b31e;
    11'b00111111000: data <= 32'h3f6e35aa;
    11'b00111111001: data <= 32'h405b3c6b;
    11'b00111111010: data <= 32'h37cf395f;
    11'b00111111011: data <= 32'hbda4bbce;
    11'b00111111100: data <= 32'hbe3bc000;
    11'b00111111101: data <= 32'hb6ebbd34;
    11'b00111111110: data <= 32'h33d7b40d;
    11'b00111111111: data <= 32'h2fb7b89d;
    11'b01000000000: data <= 32'h2dabbe1c;
    11'b01000000001: data <= 32'h3323bbbf;
    11'b01000000010: data <= 32'hb5a13cb8;
    11'b01000000011: data <= 32'hbe0d4106;
    11'b01000000100: data <= 32'hbf4e3e20;
    11'b01000000101: data <= 32'hba34b4cc;
    11'b01000000110: data <= 32'h324dba68;
    11'b01000000111: data <= 32'hacf913c4;
    11'b01000001000: data <= 32'hb80b3880;
    11'b01000001001: data <= 32'h3861376f;
    11'b01000001010: data <= 32'h40b238f3;
    11'b01000001011: data <= 32'h41013cb4;
    11'b01000001100: data <= 32'h38023c42;
    11'b01000001101: data <= 32'hbd47a881;
    11'b01000001110: data <= 32'hbbecbb2e;
    11'b01000001111: data <= 32'h382eb9d8;
    11'b01000010000: data <= 32'h3c53b88c;
    11'b01000010001: data <= 32'h374ebdce;
    11'b01000010010: data <= 32'h2c9cc09a;
    11'b01000010011: data <= 32'h35b6bd46;
    11'b01000010100: data <= 32'h335d3bc8;
    11'b01000010101: data <= 32'hba103fee;
    11'b01000010110: data <= 32'hbe203905;
    11'b01000010111: data <= 32'hbd54bc75;
    11'b01000011000: data <= 32'hbbb4bc40;
    11'b01000011001: data <= 32'hbcb133b1;
    11'b01000011010: data <= 32'hbc523a61;
    11'b01000011011: data <= 32'h358534cc;
    11'b01000011100: data <= 32'h400f3310;
    11'b01000011101: data <= 32'h3f713c84;
    11'b01000011110: data <= 32'hafbb3f24;
    11'b01000011111: data <= 32'hbda83d0d;
    11'b01000100000: data <= 32'hb7ca353d;
    11'b01000100001: data <= 32'h3c98aedb;
    11'b01000100010: data <= 32'h3d4cb80a;
    11'b01000100011: data <= 32'h358dbde4;
    11'b01000100100: data <= 32'h30bec023;
    11'b01000100101: data <= 32'h3c5abc10;
    11'b01000100110: data <= 32'h3dfc3ae4;
    11'b01000100111: data <= 32'h368f3d16;
    11'b01000101000: data <= 32'hbc23b4b8;
    11'b01000101001: data <= 32'hbe1fbeb3;
    11'b01000101010: data <= 32'hbd8dbc84;
    11'b01000101011: data <= 32'hbd90328a;
    11'b01000101100: data <= 32'hbc843403;
    11'b01000101101: data <= 32'h2aa8ba0c;
    11'b01000101110: data <= 32'h3cedba01;
    11'b01000101111: data <= 32'h3a963aed;
    11'b01000110000: data <= 32'hba9d409e;
    11'b01000110001: data <= 32'hbe18402f;
    11'b01000110010: data <= 32'hb5873b85;
    11'b01000110011: data <= 32'h3b9d32bd;
    11'b01000110100: data <= 32'h390db02f;
    11'b01000110101: data <= 32'hb586b9e2;
    11'b01000110110: data <= 32'h2fdebc7b;
    11'b01000110111: data <= 32'h3f94b5e7;
    11'b01000111000: data <= 32'h41503af8;
    11'b01000111001: data <= 32'h3d333afb;
    11'b01000111010: data <= 32'hb8d3b827;
    11'b01000111011: data <= 32'hbcf5bdae;
    11'b01000111100: data <= 32'hbaf9b9e9;
    11'b01000111101: data <= 32'hb9982c46;
    11'b01000111110: data <= 32'hb9a1b98e;
    11'b01000111111: data <= 32'hb0b2c02e;
    11'b01001000000: data <= 32'h386dbf14;
    11'b01001000001: data <= 32'h32d837a9;
    11'b01001000010: data <= 32'hbbbd408a;
    11'b01001000011: data <= 32'hbd873fca;
    11'b01001000100: data <= 32'hb83d38e2;
    11'b01001000101: data <= 32'h2c1a2cb0;
    11'b01001000110: data <= 32'hb94d34d0;
    11'b01001000111: data <= 32'hbd5031c9;
    11'b01001001000: data <= 32'haea4b3a5;
    11'b01001001001: data <= 32'h406d2624;
    11'b01001001010: data <= 32'h41f43ac8;
    11'b01001001011: data <= 32'h3d823bc0;
    11'b01001001100: data <= 32'hb7b5304c;
    11'b01001001101: data <= 32'hb947b5e1;
    11'b01001001110: data <= 32'h31372afb;
    11'b01001001111: data <= 32'h34d42cb2;
    11'b01001010000: data <= 32'hb39fbd79;
    11'b01001010001: data <= 32'hb332c1ba;
    11'b01001010010: data <= 32'h36c7c074;
    11'b01001010011: data <= 32'h381e320b;
    11'b01001010100: data <= 32'hb4703ed2;
    11'b01001010101: data <= 32'hbaf53bdc;
    11'b01001010110: data <= 32'hb9f9b561;
    11'b01001010111: data <= 32'hbafdb4f3;
    11'b01001011000: data <= 32'hbf0d389b;
    11'b01001011001: data <= 32'hc01a3929;
    11'b01001011010: data <= 32'hb715b037;
    11'b01001011011: data <= 32'h3f57b4a2;
    11'b01001011100: data <= 32'h409438d1;
    11'b01001011101: data <= 32'h39453d61;
    11'b01001011110: data <= 32'hb96d3cc5;
    11'b01001011111: data <= 32'hb0613aec;
    11'b01001100000: data <= 32'h3be53aec;
    11'b01001100001: data <= 32'h3a713537;
    11'b01001100010: data <= 32'hb3d3bd35;
    11'b01001100011: data <= 32'hb51cc134;
    11'b01001100100: data <= 32'h3a8bbf7b;
    11'b01001100101: data <= 32'h3e1d30d4;
    11'b01001100110: data <= 32'h3b283bda;
    11'b01001100111: data <= 32'hb10aaf28;
    11'b01001101000: data <= 32'hb9a9bc92;
    11'b01001101001: data <= 32'hbcbbb7ef;
    11'b01001101010: data <= 32'hbfe3396e;
    11'b01001101011: data <= 32'hc03136b3;
    11'b01001101100: data <= 32'hb99bbb6b;
    11'b01001101101: data <= 32'h3c16bd05;
    11'b01001101110: data <= 32'h3c6a2edf;
    11'b01001101111: data <= 32'hb46b3e5e;
    11'b01001110000: data <= 32'hbb593f86;
    11'b01001110001: data <= 32'h2f453df1;
    11'b01001110010: data <= 32'h3c5c3ced;
    11'b01001110011: data <= 32'h360c39b6;
    11'b01001110100: data <= 32'hbb52b852;
    11'b01001110101: data <= 32'hb8a1be21;
    11'b01001110110: data <= 32'h3d4abc11;
    11'b01001110111: data <= 32'h410c34c1;
    11'b01001111000: data <= 32'h3f3b3800;
    11'b01001111001: data <= 32'h3605b8ee;
    11'b01001111010: data <= 32'hb594bca2;
    11'b01001111011: data <= 32'hb905b0b3;
    11'b01001111100: data <= 32'hbcbc3a22;
    11'b01001111101: data <= 32'hbdfdb2bb;
    11'b01001111110: data <= 32'hba25c028;
    11'b01001111111: data <= 32'h3485c09d;
    11'b01010000000: data <= 32'h3381b6db;
    11'b01010000001: data <= 32'hb98a3dbb;
    11'b01010000010: data <= 32'hbabf3eb5;
    11'b01010000011: data <= 32'h30643c5a;
    11'b01010000100: data <= 32'h38313bb9;
    11'b01010000101: data <= 32'hb9c13c21;
    11'b01010000110: data <= 32'hbfbf36bc;
    11'b01010000111: data <= 32'hbbf0b697;
    11'b01010001000: data <= 32'h3de3b585;
    11'b01010001001: data <= 32'h418935dd;
    11'b01010001010: data <= 32'h3f603696;
    11'b01010001011: data <= 32'h36b8b48f;
    11'b01010001100: data <= 32'h30ceb518;
    11'b01010001101: data <= 32'h37203977;
    11'b01010001110: data <= 32'h281a3be6;
    11'b01010001111: data <= 32'hba10b967;
    11'b01010010000: data <= 32'hb9d7c185;
    11'b01010010001: data <= 32'h9ca9c181;
    11'b01010010010: data <= 32'h32ecb992;
    11'b01010010011: data <= 32'hb37c3b42;
    11'b01010010100: data <= 32'hb4e63963;
    11'b01010010101: data <= 32'h30d3aa1c;
    11'b01010010110: data <= 32'hb17f352f;
    11'b01010010111: data <= 32'hbedb3cb5;
    11'b01010011000: data <= 32'hc15a3c0f;
    11'b01010011001: data <= 32'hbd751f46;
    11'b01010011010: data <= 32'h3c59b685;
    11'b01010011011: data <= 32'h40122f8c;
    11'b01010011100: data <= 32'h3bb8386c;
    11'b01010011101: data <= 32'ha0cc380c;
    11'b01010011110: data <= 32'h38513a5b;
    11'b01010011111: data <= 32'h3d823e24;
    11'b01010100000: data <= 32'h3ab23d50;
    11'b01010100001: data <= 32'hb7ebb875;
    11'b01010100010: data <= 32'hba64c0e6;
    11'b01010100011: data <= 32'h3134c088;
    11'b01010100100: data <= 32'h3b8bb84b;
    11'b01010100101: data <= 32'h3a6834e8;
    11'b01010100110: data <= 32'h376db81d;
    11'b01010100111: data <= 32'h353cbc93;
    11'b01010101000: data <= 32'hb62eb0a7;
    11'b01010101001: data <= 32'hbf7b3ce6;
    11'b01010101010: data <= 32'hc1423c00;
    11'b01010101011: data <= 32'hbde2b7d0;
    11'b01010101100: data <= 32'h360fbcdb;
    11'b01010101101: data <= 32'h3a23b709;
    11'b01010101110: data <= 32'hb3e638fd;
    11'b01010101111: data <= 32'hb8523c3b;
    11'b01010110000: data <= 32'h39ac3d70;
    11'b01010110001: data <= 32'h3eb23f68;
    11'b01010110010: data <= 32'h39c03e78;
    11'b01010110011: data <= 32'hbbdc300c;
    11'b01010110100: data <= 32'hbc74bd37;
    11'b01010110101: data <= 32'h3772bc9e;
    11'b01010110110: data <= 32'h3f11ae70;
    11'b01010110111: data <= 32'h3e9bacc2;
    11'b01010111000: data <= 32'h3be8bcc8;
    11'b01010111001: data <= 32'h392ebde7;
    11'b01010111010: data <= 32'h30059dfc;
    11'b01010111011: data <= 32'hbc0f3d67;
    11'b01010111100: data <= 32'hbf3238b2;
    11'b01010111101: data <= 32'hbd0abdc0;
    11'b01010111110: data <= 32'hb3eec064;
    11'b01010111111: data <= 32'hb43dbc00;
    11'b01011000000: data <= 32'hbbe5371d;
    11'b01011000001: data <= 32'hb99d3ae0;
    11'b01011000010: data <= 32'h39ff3b37;
    11'b01011000011: data <= 32'h3d503d90;
    11'b01011000100: data <= 32'hb0d43ebd;
    11'b01011000101: data <= 32'hbfaf3bc7;
    11'b01011000110: data <= 32'hbe4fa86f;
    11'b01011000111: data <= 32'h3859b0f4;
    11'b01011001000: data <= 32'h3fe83375;
    11'b01011001001: data <= 32'h3e8cb0e5;
    11'b01011001010: data <= 32'h3b0cbc56;
    11'b01011001011: data <= 32'h3b79bb19;
    11'b01011001100: data <= 32'h3c5d39ca;
    11'b01011001101: data <= 32'h35613e8c;
    11'b01011001110: data <= 32'hb9df338a;
    11'b01011001111: data <= 32'hbb7bc01a;
    11'b01011010000: data <= 32'hb7f8c130;
    11'b01011010001: data <= 32'hb800bca7;
    11'b01011010010: data <= 32'hba6e2d43;
    11'b01011010011: data <= 32'hb4a3ab0a;
    11'b01011010100: data <= 32'h3aaab5b3;
    11'b01011010101: data <= 32'h3a3d36fb;
    11'b01011010110: data <= 32'hbc313e1f;
    11'b01011010111: data <= 32'hc13e3e05;
    11'b01011011000: data <= 32'hbf8f38c4;
    11'b01011011001: data <= 32'h344f2d53;
    11'b01011011010: data <= 32'h3d3e3088;
    11'b01011011011: data <= 32'h392eace0;
    11'b01011011100: data <= 32'h3128b77b;
    11'b01011011101: data <= 32'h3c1d2e59;
    11'b01011011110: data <= 32'h3fc83e2a;
    11'b01011011111: data <= 32'h3d613fd9;
    11'b01011100000: data <= 32'hb0c234ba;
    11'b01011100001: data <= 32'hba7bbf21;
    11'b01011100010: data <= 32'hb610c007;
    11'b01011100011: data <= 32'h283cb9f4;
    11'b01011100100: data <= 32'h2cb4b3a4;
    11'b01011100101: data <= 32'h3716bca2;
    11'b01011100110: data <= 32'h3c1fbe98;
    11'b01011100111: data <= 32'h3877b5f2;
    11'b01011101000: data <= 32'hbce43d66;
    11'b01011101001: data <= 32'hc0ff3e10;
    11'b01011101010: data <= 32'hbf1b34e7;
    11'b01011101011: data <= 32'hb1ffb843;
    11'b01011101100: data <= 32'h3002b5d6;
    11'b01011101101: data <= 32'hba07aae3;
    11'b01011101110: data <= 32'hb9bd29a6;
    11'b01011101111: data <= 32'h3b853946;
    11'b01011110000: data <= 32'h407d3f37;
    11'b01011110001: data <= 32'h3dc44028;
    11'b01011110010: data <= 32'hb6973a1a;
    11'b01011110011: data <= 32'hbc33b9b7;
    11'b01011110100: data <= 32'hb071b9ca;
    11'b01011110101: data <= 32'h3a35293d;
    11'b01011110110: data <= 32'h3b28b57b;
    11'b01011110111: data <= 32'h3b78bf4b;
    11'b01011111000: data <= 32'h3cecc068;
    11'b01011111001: data <= 32'h3b2bb7d8;
    11'b01011111010: data <= 32'hb6fe3d7a;
    11'b01011111011: data <= 32'hbe053cab;
    11'b01011111100: data <= 32'hbce8b83c;
    11'b01011111101: data <= 32'hb836bdd4;
    11'b01011111110: data <= 32'hbb04bb3e;
    11'b01011111111: data <= 32'hbee4b135;
    11'b01100000000: data <= 32'hbcafa6f6;
    11'b01100000001: data <= 32'h3ab63431;
    11'b01100000010: data <= 32'h3fd53ccf;
    11'b01100000011: data <= 32'h39b13f52;
    11'b01100000100: data <= 32'hbd0e3d4a;
    11'b01100000101: data <= 32'hbdfd381f;
    11'b01100000110: data <= 32'ha83d381a;
    11'b01100000111: data <= 32'h3c433996;
    11'b01100001000: data <= 32'h3b6bb3cd;
    11'b01100001001: data <= 32'h39b6bf0c;
    11'b01100001010: data <= 32'h3cf4bf1d;
    11'b01100001011: data <= 32'h3e5c2fbe;
    11'b01100001100: data <= 32'h3af13e89;
    11'b01100001101: data <= 32'hb27f3a91;
    11'b01100001110: data <= 32'hb86bbcb9;
    11'b01100001111: data <= 32'hb884bf91;
    11'b01100010000: data <= 32'hbc9abbe1;
    11'b01100010001: data <= 32'hbeeab4ab;
    11'b01100010010: data <= 32'hbb51b98f;
    11'b01100010011: data <= 32'h3b1abb93;
    11'b01100010100: data <= 32'h3dbf24b0;
    11'b01100010101: data <= 32'hb1f13d3f;
    11'b01100010110: data <= 32'hbff23e75;
    11'b01100010111: data <= 32'hbf043cb0;
    11'b01100011000: data <= 32'hafd53bb7;
    11'b01100011001: data <= 32'h38ea3a72;
    11'b01100011010: data <= 32'ha1c2aeed;
    11'b01100011011: data <= 32'hb30dbcc0;
    11'b01100011100: data <= 32'h3bc1ba9c;
    11'b01100011101: data <= 32'h405e3b8d;
    11'b01100011110: data <= 32'h3f913fb5;
    11'b01100011111: data <= 32'h38f139f1;
    11'b01100100000: data <= 32'hb1d3bc5e;
    11'b01100100001: data <= 32'hb5acbd72;
    11'b01100100010: data <= 32'hb959b5fa;
    11'b01100100011: data <= 32'hbb5fb439;
    11'b01100100100: data <= 32'hb259be21;
    11'b01100100101: data <= 32'h3c48c07e;
    11'b01100100110: data <= 32'h3c7cbc2b;
    11'b01100100111: data <= 32'hb80d3abe;
    11'b01100101000: data <= 32'hbfa93dfd;
    11'b01100101001: data <= 32'hbde83b7d;
    11'b01100101010: data <= 32'hb4173745;
    11'b01100101011: data <= 32'hb4f3358f;
    11'b01100101100: data <= 32'hbda7ad04;
    11'b01100101101: data <= 32'hbd73b8f7;
    11'b01100101110: data <= 32'h3876b0e4;
    11'b01100101111: data <= 32'h40a43d0b;
    11'b01100110000: data <= 32'h40143fa8;
    11'b01100110001: data <= 32'h37f43b5d;
    11'b01100110010: data <= 32'hb553b460;
    11'b01100110011: data <= 32'hae77acb9;
    11'b01100110100: data <= 32'h2e3b396d;
    11'b01100110101: data <= 32'ha562a523;
    11'b01100110110: data <= 32'h3591c003;
    11'b01100110111: data <= 32'h3cb5c1b3;
    11'b01100111000: data <= 32'h3cd7bd5a;
    11'b01100111001: data <= 32'h29a639d2;
    11'b01100111010: data <= 32'hbb763c78;
    11'b01100111011: data <= 32'hb9532e6c;
    11'b01100111100: data <= 32'hb37db81b;
    11'b01100111101: data <= 32'hbc67b3c0;
    11'b01100111110: data <= 32'hc0deb014;
    11'b01100111111: data <= 32'hc00eb7cd;
    11'b01101000000: data <= 32'h3460b558;
    11'b01101000001: data <= 32'h3fe93977;
    11'b01101000010: data <= 32'h3d4e3daf;
    11'b01101000011: data <= 32'hb5ca3c79;
    11'b01101000100: data <= 32'hba8239d9;
    11'b01101000101: data <= 32'h29173cdb;
    11'b01101000110: data <= 32'h38633e52;
    11'b01101000111: data <= 32'h329634f3;
    11'b01101001000: data <= 32'h3153bf71;
    11'b01101001001: data <= 32'h3bc2c0e9;
    11'b01101001010: data <= 32'h3e38ba12;
    11'b01101001011: data <= 32'h3c773c01;
    11'b01101001100: data <= 32'h36b839fe;
    11'b01101001101: data <= 32'h347bb964;
    11'b01101001110: data <= 32'h19d9bc78;
    11'b01101001111: data <= 32'hbd0db5f9;
    11'b01101010000: data <= 32'hc0f7acf9;
    11'b01101010001: data <= 32'hbf61baa4;
    11'b01101010010: data <= 32'h34c2bd3c;
    11'b01101010011: data <= 32'h3dc0b85b;
    11'b01101010100: data <= 32'h356538ee;
    11'b01101010101: data <= 32'hbceb3c65;
    11'b01101010110: data <= 32'hbc883d01;
    11'b01101010111: data <= 32'h2de33ee5;
    11'b01101011000: data <= 32'h36403f3c;
    11'b01101011001: data <= 32'hb8063817;
    11'b01101011010: data <= 32'hba66bd0d;
    11'b01101011011: data <= 32'h3696bdc1;
    11'b01101011100: data <= 32'h3f4031e0;
    11'b01101011101: data <= 32'h3fed3d71;
    11'b01101011110: data <= 32'h3d3f3882;
    11'b01101011111: data <= 32'h3a90bac3;
    11'b01101100000: data <= 32'h3541ba7c;
    11'b01101100001: data <= 32'hb9f7340f;
    11'b01101100010: data <= 32'hbe8e334b;
    11'b01101100011: data <= 32'hbc2abd47;
    11'b01101100100: data <= 32'h385cc0dd;
    11'b01101100101: data <= 32'h3c2dbebe;
    11'b01101100110: data <= 32'hb2c6ac60;
    11'b01101100111: data <= 32'hbd7f3a83;
    11'b01101101000: data <= 32'hbade3bb3;
    11'b01101101001: data <= 32'h32e43cd0;
    11'b01101101010: data <= 32'hb1ff3d36;
    11'b01101101011: data <= 32'hbee037d7;
    11'b01101101100: data <= 32'hc00eb920;
    11'b01101101101: data <= 32'hb407b88c;
    11'b01101101110: data <= 32'h3eee39af;
    11'b01101101111: data <= 32'h401c3d7e;
    11'b01101110000: data <= 32'h3cd4381b;
    11'b01101110001: data <= 32'h395bb5ce;
    11'b01101110010: data <= 32'h38743488;
    11'b01101110011: data <= 32'h2bdd3d91;
    11'b01101110100: data <= 32'hb89339ff;
    11'b01101110101: data <= 32'hb4bbbe26;
    11'b01101110110: data <= 32'h3998c1e3;
    11'b01101110111: data <= 32'h3b80c00b;
    11'b01101111000: data <= 32'h24a3b394;
    11'b01101111001: data <= 32'hb8bd36bc;
    11'b01101111010: data <= 32'h28212dc6;
    11'b01101111011: data <= 32'h383d2e7c;
    11'b01101111100: data <= 32'hb9893840;
    11'b01101111101: data <= 32'hc1433600;
    11'b01101111110: data <= 32'hc184b58c;
    11'b01101111111: data <= 32'hb926b728;
    11'b01110000000: data <= 32'h3d533577;
    11'b01110000001: data <= 32'h3d363a89;
    11'b01110000010: data <= 32'h33d436a5;
    11'b01110000011: data <= 32'h2867355b;
    11'b01110000100: data <= 32'h38ff3dd0;
    11'b01110000101: data <= 32'h392140c3;
    11'b01110000110: data <= 32'hac243cf4;
    11'b01110000111: data <= 32'hb424bd27;
    11'b01110001000: data <= 32'h373fc101;
    11'b01110001001: data <= 32'h3bf6bd7c;
    11'b01110001010: data <= 32'h3a2a30fa;
    11'b01110001011: data <= 32'h390b2fb2;
    11'b01110001100: data <= 32'h3c57ba4d;
    11'b01110001101: data <= 32'h3bcbba14;
    11'b01110001110: data <= 32'hb9a831a0;
    11'b01110001111: data <= 32'hc14136f5;
    11'b01110010000: data <= 32'hc113b6c8;
    11'b01110010001: data <= 32'hb85abc63;
    11'b01110010010: data <= 32'h3abdb9f1;
    11'b01110010011: data <= 32'h3343aec1;
    11'b01110010100: data <= 32'hbada30ba;
    11'b01110010101: data <= 32'hb8143954;
    11'b01110010110: data <= 32'h39453f9e;
    11'b01110010111: data <= 32'h39c44139;
    11'b01110011000: data <= 32'hb7343dab;
    11'b01110011001: data <= 32'hbc43b9b9;
    11'b01110011010: data <= 32'hb30abda4;
    11'b01110011011: data <= 32'h3bd2b30a;
    11'b01110011100: data <= 32'h3da539e0;
    11'b01110011101: data <= 32'h3dd6a66d;
    11'b01110011110: data <= 32'h3eaabcad;
    11'b01110011111: data <= 32'h3d55ba29;
    11'b01110100000: data <= 32'hb1cf3903;
    11'b01110100001: data <= 32'hbedd3abb;
    11'b01110100010: data <= 32'hbe37b901;
    11'b01110100011: data <= 32'hadd3bfdf;
    11'b01110100100: data <= 32'h3806bf41;
    11'b01110100101: data <= 32'hb80ebaef;
    11'b01110100110: data <= 32'hbd3eb35c;
    11'b01110100111: data <= 32'hb6dd354c;
    11'b01110101000: data <= 32'h3ae63d4c;
    11'b01110101001: data <= 32'h36e63fd7;
    11'b01110101010: data <= 32'hbd933cdb;
    11'b01110101011: data <= 32'hc06db0ed;
    11'b01110101100: data <= 32'hbbe8b605;
    11'b01110101101: data <= 32'h39ff38e0;
    11'b01110101110: data <= 32'h3d983bab;
    11'b01110101111: data <= 32'h3d35b029;
    11'b01110110000: data <= 32'h3da8bbbb;
    11'b01110110001: data <= 32'h3dac28dc;
    11'b01110110010: data <= 32'h388c3eb2;
    11'b01110110011: data <= 32'hb80c3df2;
    11'b01110110100: data <= 32'hb821b932;
    11'b01110110101: data <= 32'h34a8c0b5;
    11'b01110110110: data <= 32'h35edc035;
    11'b01110110111: data <= 32'hb85bbbd9;
    11'b01110111000: data <= 32'hba9db83c;
    11'b01110111001: data <= 32'h35afb7fd;
    11'b01110111010: data <= 32'h3d3b2e2c;
    11'b01110111011: data <= 32'h30f33b51;
    11'b01110111100: data <= 32'hc04c3ae5;
    11'b01110111101: data <= 32'hc1ce3072;
    11'b01110111110: data <= 32'hbd7d99a4;
    11'b01110111111: data <= 32'h362f3866;
    11'b01111000000: data <= 32'h394e383d;
    11'b01111000001: data <= 32'h3355b5b5;
    11'b01111000010: data <= 32'h383db82b;
    11'b01111000011: data <= 32'h3d013c19;
    11'b01111000100: data <= 32'h3c804140;
    11'b01111000101: data <= 32'h33924006;
    11'b01111000110: data <= 32'hb11cb619;
    11'b01111000111: data <= 32'h3262bf9b;
    11'b01111001000: data <= 32'h34ffbd6d;
    11'b01111001001: data <= 32'habc0b5fc;
    11'b01111001010: data <= 32'h320cb8e5;
    11'b01111001011: data <= 32'h3d7dbd5d;
    11'b01111001100: data <= 32'h3f51bbdb;
    11'b01111001101: data <= 32'h32ce3374;
    11'b01111001110: data <= 32'hc03639e7;
    11'b01111001111: data <= 32'hc13530f8;
    11'b01111010000: data <= 32'hbc67b608;
    11'b01111010001: data <= 32'h2d8bb4da;
    11'b01111010010: data <= 32'hb601b5a1;
    11'b01111010011: data <= 32'hbc4ab9de;
    11'b01111010100: data <= 32'hb572b4fd;
    11'b01111010101: data <= 32'h3c4e3da5;
    11'b01111010110: data <= 32'h3d164197;
    11'b01111010111: data <= 32'h300c4021;
    11'b01111011000: data <= 32'hb9b02942;
    11'b01111011001: data <= 32'hb6adbaba;
    11'b01111011010: data <= 32'h314aa4f7;
    11'b01111011011: data <= 32'h36a33832;
    11'b01111011100: data <= 32'h3b6cb83d;
    11'b01111011101: data <= 32'h3fa8bf0e;
    11'b01111011110: data <= 32'h403bbd0d;
    11'b01111011111: data <= 32'h3911367b;
    11'b01111100000: data <= 32'hbcdc3c42;
    11'b01111100001: data <= 32'hbdcc2db6;
    11'b01111100010: data <= 32'hb577bc31;
    11'b01111100011: data <= 32'ha4b3bd09;
    11'b01111100100: data <= 32'hbc86bc5d;
    11'b01111100101: data <= 32'hbf2dbc5f;
    11'b01111100110: data <= 32'hb87ab8be;
    11'b01111100111: data <= 32'h3cae3ab6;
    11'b01111101000: data <= 32'h3c723ffd;
    11'b01111101001: data <= 32'hb8be3e54;
    11'b01111101010: data <= 32'hbedf35f0;
    11'b01111101011: data <= 32'hbcb23274;
    11'b01111101100: data <= 32'hae083c4a;
    11'b01111101101: data <= 32'h36773c46;
    11'b01111101110: data <= 32'h3a1ab7ec;
    11'b01111101111: data <= 32'h3e2bbeb7;
    11'b01111110000: data <= 32'h3fd5b992;
    11'b01111110001: data <= 32'h3caa3d24;
    11'b01111110010: data <= 32'h9cd23ecb;
    11'b01111110011: data <= 32'hb0f6305b;
    11'b01111110100: data <= 32'h360bbd8c;
    11'b01111110101: data <= 32'h24dbbe19;
    11'b01111110110: data <= 32'hbd15bc76;
    11'b01111110111: data <= 32'hbe42bccb;
    11'b01111111000: data <= 32'h27bfbcef;
    11'b01111111001: data <= 32'h3e63b62b;
    11'b01111111010: data <= 32'h3b7839a5;
    11'b01111111011: data <= 32'hbd093b11;
    11'b01111111100: data <= 32'hc0bb3779;
    11'b01111111101: data <= 32'hbdfe3948;
    11'b01111111110: data <= 32'hb5143d20;
    11'b01111111111: data <= 32'hb1bc3aec;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    