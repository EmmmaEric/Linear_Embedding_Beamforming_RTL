
module memory_rom_13(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hb8a33de9;
    11'b00000000001: data <= 32'hb4583a58;
    11'b00000000010: data <= 32'h36bcbb36;
    11'b00000000011: data <= 32'h3dc8bcc7;
    11'b00000000100: data <= 32'h3e8838b5;
    11'b00000000101: data <= 32'h39e74080;
    11'b00000000110: data <= 32'h2f643f27;
    11'b00000000111: data <= 32'h388e253c;
    11'b00000001000: data <= 32'h3b5fbbf8;
    11'b00000001001: data <= 32'ha6f9bb76;
    11'b00000001010: data <= 32'hbcd0bc03;
    11'b00000001011: data <= 32'hb921be0c;
    11'b00000001100: data <= 32'h3d40bdbc;
    11'b00000001101: data <= 32'h402cb780;
    11'b00000001110: data <= 32'h377233e6;
    11'b00000001111: data <= 32'hbeb62b47;
    11'b00000010000: data <= 32'hc031adb0;
    11'b00000010001: data <= 32'hbc8e38a6;
    11'b00000010010: data <= 32'hb9403c1e;
    11'b00000010011: data <= 32'hbc012692;
    11'b00000010100: data <= 32'hbaedbdaa;
    11'b00000010101: data <= 32'h32a8bc47;
    11'b00000010110: data <= 32'h3c253c9d;
    11'b00000010111: data <= 32'h3aa54179;
    11'b00000011000: data <= 32'h36573fec;
    11'b00000011001: data <= 32'h381a33d5;
    11'b00000011010: data <= 32'h3817b474;
    11'b00000011011: data <= 32'hb4d53487;
    11'b00000011100: data <= 32'hbb1f30ce;
    11'b00000011101: data <= 32'h31c0bc2f;
    11'b00000011110: data <= 32'h403ebf10;
    11'b00000011111: data <= 32'h4107bc72;
    11'b00000100000: data <= 32'h3996af98;
    11'b00000100001: data <= 32'hbca52e78;
    11'b00000100010: data <= 32'hbc99a8c1;
    11'b00000100011: data <= 32'hb308314f;
    11'b00000100100: data <= 32'hb6a82fdf;
    11'b00000100101: data <= 32'hbe80bb44;
    11'b00000100110: data <= 32'hbf88bfb0;
    11'b00000100111: data <= 32'hb84abcbf;
    11'b00000101000: data <= 32'h3a733bce;
    11'b00000101001: data <= 32'h3a31406d;
    11'b00000101010: data <= 32'h241d3d9f;
    11'b00000101011: data <= 32'hb4d033d3;
    11'b00000101100: data <= 32'hb57838a2;
    11'b00000101101: data <= 32'hb9b53e5b;
    11'b00000101110: data <= 32'hba583cad;
    11'b00000101111: data <= 32'h3644b975;
    11'b00000110000: data <= 32'h4023bf16;
    11'b00000110001: data <= 32'h40a2bb81;
    11'b00000110010: data <= 32'h3b26371d;
    11'b00000110011: data <= 32'hb2b839d1;
    11'b00000110100: data <= 32'h3436312d;
    11'b00000110101: data <= 32'h3b4cb23a;
    11'b00000110110: data <= 32'habadb730;
    11'b00000110111: data <= 32'hbf64bd0a;
    11'b00000111000: data <= 32'hc026c010;
    11'b00000111001: data <= 32'hb585bded;
    11'b00000111010: data <= 32'h3c922e51;
    11'b00000111011: data <= 32'h39fa3b4d;
    11'b00000111100: data <= 32'hb89a35b1;
    11'b00000111101: data <= 32'hbc912549;
    11'b00000111110: data <= 32'hbba43c66;
    11'b00000111111: data <= 32'hbbca4073;
    11'b00001000000: data <= 32'hbc2c3da3;
    11'b00001000001: data <= 32'hb421b9e7;
    11'b00001000010: data <= 32'h3c41be6d;
    11'b00001000011: data <= 32'h3e15b3ec;
    11'b00001000100: data <= 32'h3b243d9f;
    11'b00001000101: data <= 32'h38d53dbf;
    11'b00001000110: data <= 32'h3d343656;
    11'b00001000111: data <= 32'h3e2eb0b6;
    11'b00001001000: data <= 32'h2e62b0c6;
    11'b00001001001: data <= 32'hbebcb932;
    11'b00001001010: data <= 32'hbdefbe47;
    11'b00001001011: data <= 32'h3859beea;
    11'b00001001100: data <= 32'h3f2dbb87;
    11'b00001001101: data <= 32'h3aa0b63b;
    11'b00001001110: data <= 32'hbabdb838;
    11'b00001001111: data <= 32'hbd0fb378;
    11'b00001010000: data <= 32'hba0a3c4e;
    11'b00001010001: data <= 32'hba873fae;
    11'b00001010010: data <= 32'hbde13a4d;
    11'b00001010011: data <= 32'hbd9cbccf;
    11'b00001010100: data <= 32'hb525bdf3;
    11'b00001010101: data <= 32'h38ad3572;
    11'b00001010110: data <= 32'h39a13fc4;
    11'b00001010111: data <= 32'h3ab73e63;
    11'b00001011000: data <= 32'h3d9c36df;
    11'b00001011001: data <= 32'h3d4534d9;
    11'b00001011010: data <= 32'hae6b3b6f;
    11'b00001011011: data <= 32'hbd8d3923;
    11'b00001011100: data <= 32'hb96aba14;
    11'b00001011101: data <= 32'h3d81bf01;
    11'b00001011110: data <= 32'h4069be10;
    11'b00001011111: data <= 32'h3b53bb65;
    11'b00001100000: data <= 32'hb86ab9aa;
    11'b00001100001: data <= 32'hb71bb4a7;
    11'b00001100010: data <= 32'h34a23975;
    11'b00001100011: data <= 32'hb39b3c3e;
    11'b00001100100: data <= 32'hbf15b094;
    11'b00001100101: data <= 32'hc0abbece;
    11'b00001100110: data <= 32'hbcfabe02;
    11'b00001100111: data <= 32'h2dac358c;
    11'b00001101000: data <= 32'h37f13e21;
    11'b00001101001: data <= 32'h37953b4c;
    11'b00001101010: data <= 32'h39542f13;
    11'b00001101011: data <= 32'h37fc3ab3;
    11'b00001101100: data <= 32'hb8104046;
    11'b00001101101: data <= 32'hbce93f62;
    11'b00001101110: data <= 32'hb527ae04;
    11'b00001101111: data <= 32'h3db6be41;
    11'b00001110000: data <= 32'h3fadbd60;
    11'b00001110001: data <= 32'h3a92b774;
    11'b00001110010: data <= 32'h2d8fb0ec;
    11'b00001110011: data <= 32'h3af0ae9e;
    11'b00001110100: data <= 32'h3e7034a4;
    11'b00001110101: data <= 32'h372b362f;
    11'b00001110110: data <= 32'hbf0bb8b5;
    11'b00001110111: data <= 32'hc106beff;
    11'b00001111000: data <= 32'hbcbabe2d;
    11'b00001111001: data <= 32'h34f4b398;
    11'b00001111010: data <= 32'h36ff355c;
    11'b00001111011: data <= 32'hb012b52e;
    11'b00001111100: data <= 32'hb39ab763;
    11'b00001111101: data <= 32'hb22f3c60;
    11'b00001111110: data <= 32'hb9e0417d;
    11'b00001111111: data <= 32'hbd14407a;
    11'b00010000000: data <= 32'hb9a3226d;
    11'b00010000001: data <= 32'h3839bd57;
    11'b00010000010: data <= 32'h3b91b93c;
    11'b00010000011: data <= 32'h376c382d;
    11'b00010000100: data <= 32'h38ec38ea;
    11'b00010000101: data <= 32'h3f782f9c;
    11'b00010000110: data <= 32'h40d63199;
    11'b00010000111: data <= 32'h3a893732;
    11'b00010001000: data <= 32'hbdfead8e;
    11'b00010001001: data <= 32'hbfb1bc85;
    11'b00010001010: data <= 32'hb4d1bdc4;
    11'b00010001011: data <= 32'h3bf2bbd5;
    11'b00010001100: data <= 32'h3825bb60;
    11'b00010001101: data <= 32'hb81fbd9f;
    11'b00010001110: data <= 32'hb882bbc6;
    11'b00010001111: data <= 32'haead3b78;
    11'b00010010000: data <= 32'hb72340e3;
    11'b00010010001: data <= 32'hbd773ea1;
    11'b00010010010: data <= 32'hbe30b73b;
    11'b00010010011: data <= 32'hba70bcde;
    11'b00010010100: data <= 32'hb2902570;
    11'b00010010101: data <= 32'ha5f33ce9;
    11'b00010010110: data <= 32'h39693b16;
    11'b00010010111: data <= 32'h3fe22acf;
    11'b00010011000: data <= 32'h40893539;
    11'b00010011001: data <= 32'h39433cef;
    11'b00010011010: data <= 32'hbcc63c93;
    11'b00010011011: data <= 32'hbc37ae4f;
    11'b00010011100: data <= 32'h395ebc88;
    11'b00010011101: data <= 32'h3e0cbd61;
    11'b00010011110: data <= 32'h384bbdd5;
    11'b00010011111: data <= 32'hb7c8becf;
    11'b00010100000: data <= 32'ha61dbc79;
    11'b00010100001: data <= 32'h3af63817;
    11'b00010100010: data <= 32'h35933e2c;
    11'b00010100011: data <= 32'hbd4538f2;
    11'b00010100100: data <= 32'hc07cbc35;
    11'b00010100101: data <= 32'hbee8bcc2;
    11'b00010100110: data <= 32'hbad93406;
    11'b00010100111: data <= 32'hb5fa3c53;
    11'b00010101000: data <= 32'h34173481;
    11'b00010101001: data <= 32'h3cd6b779;
    11'b00010101010: data <= 32'h3d813810;
    11'b00010101011: data <= 32'h31324060;
    11'b00010101100: data <= 32'hbc0d40b0;
    11'b00010101101: data <= 32'hb8163a0d;
    11'b00010101110: data <= 32'h3bbfb9fb;
    11'b00010101111: data <= 32'h3d46bc56;
    11'b00010110000: data <= 32'h343abbe5;
    11'b00010110001: data <= 32'hb227bc76;
    11'b00010110010: data <= 32'h3c18baf2;
    11'b00010110011: data <= 32'h405e2f2f;
    11'b00010110100: data <= 32'h3cff39b4;
    11'b00010110101: data <= 32'hbc3eab1c;
    11'b00010110110: data <= 32'hc098bcd3;
    11'b00010110111: data <= 32'hbea6bc55;
    11'b00010111000: data <= 32'hb92d9cbf;
    11'b00010111001: data <= 32'hb68630e1;
    11'b00010111010: data <= 32'hb59fbb8c;
    11'b00010111011: data <= 32'h31c5bd16;
    11'b00010111100: data <= 32'h379e37a8;
    11'b00010111101: data <= 32'hb1db4148;
    11'b00010111110: data <= 32'hbb83417c;
    11'b00010111111: data <= 32'hb8b53b60;
    11'b00011000000: data <= 32'h3569b7f4;
    11'b00011000001: data <= 32'h35ddb60e;
    11'b00011000010: data <= 32'hb5562e61;
    11'b00011000011: data <= 32'h25afb151;
    11'b00011000100: data <= 32'h3f63b82b;
    11'b00011000101: data <= 32'h4205ad74;
    11'b00011000110: data <= 32'h3ee637fd;
    11'b00011000111: data <= 32'hb9c931a6;
    11'b00011001000: data <= 32'hbeb1b900;
    11'b00011001001: data <= 32'hb9a2b9f4;
    11'b00011001010: data <= 32'h31eab6a1;
    11'b00011001011: data <= 32'hb2a7bb45;
    11'b00011001100: data <= 32'hba5bc01b;
    11'b00011001101: data <= 32'hb64abfbc;
    11'b00011001110: data <= 32'h34c3321e;
    11'b00011001111: data <= 32'h29c74091;
    11'b00011010000: data <= 32'hba8a4036;
    11'b00011010001: data <= 32'hbc5e3590;
    11'b00011010010: data <= 32'hba43b7ae;
    11'b00011010011: data <= 32'hba8d355c;
    11'b00011010100: data <= 32'hbc0e3c19;
    11'b00011010101: data <= 32'hae1035de;
    11'b00011010110: data <= 32'h3f7cb805;
    11'b00011010111: data <= 32'h41a6b000;
    11'b00011011000: data <= 32'h3e003b95;
    11'b00011011001: data <= 32'hb7e13cb9;
    11'b00011011010: data <= 32'hba303708;
    11'b00011011011: data <= 32'h3760b2bf;
    11'b00011011100: data <= 32'h3ba5b873;
    11'b00011011101: data <= 32'had71bd61;
    11'b00011011110: data <= 32'hbb68c0ae;
    11'b00011011111: data <= 32'hb1a5c021;
    11'b00011100000: data <= 32'h3c22b236;
    11'b00011100001: data <= 32'h3ae63d67;
    11'b00011100010: data <= 32'hb8343b2e;
    11'b00011100011: data <= 32'hbe19b7d9;
    11'b00011100100: data <= 32'hbe57b891;
    11'b00011100101: data <= 32'hbdf23992;
    11'b00011100110: data <= 32'hbda03cbe;
    11'b00011100111: data <= 32'hb8302225;
    11'b00011101000: data <= 32'h3c4cbc1d;
    11'b00011101001: data <= 32'h3f28b214;
    11'b00011101010: data <= 32'h3a4e3e73;
    11'b00011101011: data <= 32'hb6fd407c;
    11'b00011101100: data <= 32'haffb3d55;
    11'b00011101101: data <= 32'h3c343460;
    11'b00011101110: data <= 32'h3c16b395;
    11'b00011101111: data <= 32'hb571baa5;
    11'b00011110000: data <= 32'hbaf6be90;
    11'b00011110001: data <= 32'h3888be87;
    11'b00011110010: data <= 32'h4062b78d;
    11'b00011110011: data <= 32'h3f4436fa;
    11'b00011110100: data <= 32'hafb8aad8;
    11'b00011110101: data <= 32'hbde1bb51;
    11'b00011110110: data <= 32'hbdddb810;
    11'b00011110111: data <= 32'hbccb394d;
    11'b00011111000: data <= 32'hbd34388e;
    11'b00011111001: data <= 32'hbc1abc2b;
    11'b00011111010: data <= 32'ha648bf93;
    11'b00011111011: data <= 32'h390ab683;
    11'b00011111100: data <= 32'h314c3fa5;
    11'b00011111101: data <= 32'hb6f34126;
    11'b00011111110: data <= 32'h0d4a3dd1;
    11'b00011111111: data <= 32'h39e736ff;
    11'b00100000000: data <= 32'h341d3649;
    11'b00100000001: data <= 32'hbbfa350f;
    11'b00100000010: data <= 32'hbaf8b742;
    11'b00100000011: data <= 32'h3cc9bc08;
    11'b00100000100: data <= 32'h41e1b897;
    11'b00100000101: data <= 32'h4090297d;
    11'b00100000110: data <= 32'h3204b085;
    11'b00100000111: data <= 32'hbb14b856;
    11'b00100001000: data <= 32'hb737afc0;
    11'b00100001001: data <= 32'hb0fa37c8;
    11'b00100001010: data <= 32'hbab2b44c;
    11'b00100001011: data <= 32'hbd6dc022;
    11'b00100001100: data <= 32'hba08c127;
    11'b00100001101: data <= 32'h3037b9c7;
    11'b00100001110: data <= 32'h311d3e33;
    11'b00100001111: data <= 32'hb4923f87;
    11'b00100010000: data <= 32'hb4373999;
    11'b00100010001: data <= 32'hb04932e6;
    11'b00100010010: data <= 32'hbaa93bec;
    11'b00100010011: data <= 32'hbee93d82;
    11'b00100010100: data <= 32'hbc483650;
    11'b00100010101: data <= 32'h3cb5b9dc;
    11'b00100010110: data <= 32'h4167b8e5;
    11'b00100010111: data <= 32'h3fa63413;
    11'b00100011000: data <= 32'h32ec38bc;
    11'b00100011001: data <= 32'hadf33694;
    11'b00100011010: data <= 32'h3aaf37bc;
    11'b00100011011: data <= 32'h3b62379b;
    11'b00100011100: data <= 32'hb704b8fb;
    11'b00100011101: data <= 32'hbdd3c09b;
    11'b00100011110: data <= 32'hba1ac137;
    11'b00100011111: data <= 32'h389fbb99;
    11'b00100100000: data <= 32'h3ac039ab;
    11'b00100100001: data <= 32'h2d6d387f;
    11'b00100100010: data <= 32'hb834b6f1;
    11'b00100100011: data <= 32'hba89b124;
    11'b00100100100: data <= 32'hbdd03d2d;
    11'b00100100101: data <= 32'hc0213f00;
    11'b00100100110: data <= 32'hbd933580;
    11'b00100100111: data <= 32'h372bbc63;
    11'b00100101000: data <= 32'h3e43b9ff;
    11'b00100101001: data <= 32'h3b6339c6;
    11'b00100101010: data <= 32'ha30d3e00;
    11'b00100101011: data <= 32'h37ae3d08;
    11'b00100101100: data <= 32'h3e7f3ba7;
    11'b00100101101: data <= 32'h3d3939fa;
    11'b00100101110: data <= 32'hb807b0b9;
    11'b00100101111: data <= 32'hbdd4be10;
    11'b00100110000: data <= 32'hb37bbfb1;
    11'b00100110001: data <= 32'h3e36bb9f;
    11'b00100110010: data <= 32'h3efcafa3;
    11'b00100110011: data <= 32'h3823b89f;
    11'b00100110100: data <= 32'hb760bcc0;
    11'b00100110101: data <= 32'hb9a6b515;
    11'b00100110110: data <= 32'hbc5e3d2f;
    11'b00100110111: data <= 32'hbefd3d6b;
    11'b00100111000: data <= 32'hbe94b802;
    11'b00100111001: data <= 32'hb87bbf99;
    11'b00100111010: data <= 32'h3345bc16;
    11'b00100111011: data <= 32'ha8d33bad;
    11'b00100111100: data <= 32'hb42b3f3d;
    11'b00100111101: data <= 32'h38f03d49;
    11'b00100111110: data <= 32'h3e273ba6;
    11'b00100111111: data <= 32'h3a373ca7;
    11'b00101000000: data <= 32'hbc523b4f;
    11'b00101000001: data <= 32'hbe1fb136;
    11'b00101000010: data <= 32'h34b3bbaf;
    11'b00101000011: data <= 32'h407fba40;
    11'b00101000100: data <= 32'h4055b802;
    11'b00101000101: data <= 32'h39b0bb28;
    11'b00101000110: data <= 32'ha94ebc51;
    11'b00101000111: data <= 32'h338aa881;
    11'b00101001000: data <= 32'h2e793ccb;
    11'b00101001001: data <= 32'hbba3393b;
    11'b00101001010: data <= 32'hbec2bdc7;
    11'b00101001011: data <= 32'hbd06c11a;
    11'b00101001100: data <= 32'hb801bd15;
    11'b00101001101: data <= 32'hb56639b4;
    11'b00101001110: data <= 32'hb3f43caf;
    11'b00101001111: data <= 32'h36dd36f2;
    11'b00101010000: data <= 32'h3aa436da;
    11'b00101010001: data <= 32'hb2953de7;
    11'b00101010010: data <= 32'hbf263fb4;
    11'b00101010011: data <= 32'hbed43b4f;
    11'b00101010100: data <= 32'h3571b5cf;
    11'b00101010101: data <= 32'h4018b929;
    11'b00101010110: data <= 32'h3ebeb5a3;
    11'b00101010111: data <= 32'h3776b593;
    11'b00101011000: data <= 32'h37acb434;
    11'b00101011001: data <= 32'h3dde385c;
    11'b00101011010: data <= 32'h3d9d3cd1;
    11'b00101011011: data <= 32'hb2d8347c;
    11'b00101011100: data <= 32'hbe50becf;
    11'b00101011101: data <= 32'hbd3ec0fc;
    11'b00101011110: data <= 32'hb42bbd11;
    11'b00101011111: data <= 32'h31942f82;
    11'b00101100000: data <= 32'h2d89adea;
    11'b00101100001: data <= 32'h32cdbb56;
    11'b00101100010: data <= 32'h317cb4d8;
    11'b00101100011: data <= 32'hbaa43e28;
    11'b00101100100: data <= 32'hc02040a6;
    11'b00101100101: data <= 32'hbf643c55;
    11'b00101100110: data <= 32'hb1a7b824;
    11'b00101100111: data <= 32'h3bb5b9cc;
    11'b00101101000: data <= 32'h37d02aa0;
    11'b00101101001: data <= 32'hafb937ee;
    11'b00101101010: data <= 32'h3a58388b;
    11'b00101101011: data <= 32'h40883bdb;
    11'b00101101100: data <= 32'h400a3d60;
    11'b00101101101: data <= 32'ha7de38a6;
    11'b00101101110: data <= 32'hbdf6bbb6;
    11'b00101101111: data <= 32'hbaccbe79;
    11'b00101110000: data <= 32'h38edbb5f;
    11'b00101110001: data <= 32'h3c25b712;
    11'b00101110010: data <= 32'h3802bcee;
    11'b00101110011: data <= 32'h3245bfac;
    11'b00101110100: data <= 32'h30c8b9f6;
    11'b00101110101: data <= 32'hb8213dac;
    11'b00101110110: data <= 32'hbe533ffc;
    11'b00101110111: data <= 32'hbf1835e1;
    11'b00101111000: data <= 32'hbb55bd02;
    11'b00101111001: data <= 32'hb5e4bbe4;
    11'b00101111010: data <= 32'hb9d7353d;
    11'b00101111011: data <= 32'hb97f3b2a;
    11'b00101111100: data <= 32'h3a2d3965;
    11'b00101111101: data <= 32'h407b3ace;
    11'b00101111110: data <= 32'h3e983de2;
    11'b00101111111: data <= 32'hb80b3d8a;
    11'b00110000000: data <= 32'hbe333602;
    11'b00110000001: data <= 32'hb515b64e;
    11'b00110000010: data <= 32'h3d74b670;
    11'b00110000011: data <= 32'h3dfab910;
    11'b00110000100: data <= 32'h38c9be6c;
    11'b00110000101: data <= 32'h35efbffc;
    11'b00110000110: data <= 32'h3ad7b8d4;
    11'b00110000111: data <= 32'h39423d2c;
    11'b00110001000: data <= 32'hb8433d41;
    11'b00110001001: data <= 32'hbdd0b8bd;
    11'b00110001010: data <= 32'hbd95bfb9;
    11'b00110001011: data <= 32'hbc96bcae;
    11'b00110001100: data <= 32'hbcfd3471;
    11'b00110001101: data <= 32'hbae43778;
    11'b00110001110: data <= 32'h3849b1fd;
    11'b00110001111: data <= 32'h3e482d59;
    11'b00110010000: data <= 32'h39793dab;
    11'b00110010001: data <= 32'hbce84052;
    11'b00110010010: data <= 32'hbec03dfc;
    11'b00110010011: data <= 32'hafb63732;
    11'b00110010100: data <= 32'h3d5da81f;
    11'b00110010101: data <= 32'h3c2db686;
    11'b00110010110: data <= 32'h3073bc70;
    11'b00110010111: data <= 32'h3851bcf0;
    11'b00110011000: data <= 32'h3f5fa731;
    11'b00110011001: data <= 32'h3ffe3d1e;
    11'b00110011010: data <= 32'h37a03aa8;
    11'b00110011011: data <= 32'hbc40bc01;
    11'b00110011100: data <= 32'hbd5bbfa5;
    11'b00110011101: data <= 32'hbbb7bbdc;
    11'b00110011110: data <= 32'hbaa32086;
    11'b00110011111: data <= 32'hb87cb875;
    11'b00110100000: data <= 32'h34f2be4a;
    11'b00110100001: data <= 32'h3ab8bb70;
    11'b00110100010: data <= 32'hac1f3ca9;
    11'b00110100011: data <= 32'hbe3240d6;
    11'b00110100100: data <= 32'hbeb83eeb;
    11'b00110100101: data <= 32'hb57a36e3;
    11'b00110100110: data <= 32'h37d3a8b4;
    11'b00110100111: data <= 32'hb1ca20ae;
    11'b00110101000: data <= 32'hb9e0b342;
    11'b00110101001: data <= 32'h3819b4f1;
    11'b00110101010: data <= 32'h40f33765;
    11'b00110101011: data <= 32'h415e3d3c;
    11'b00110101100: data <= 32'h3ab13aff;
    11'b00110101101: data <= 32'hbad2b7bf;
    11'b00110101110: data <= 32'hbad0bc13;
    11'b00110101111: data <= 32'hacdfb5b4;
    11'b00110110000: data <= 32'h2df3b247;
    11'b00110110001: data <= 32'hae0fbe0d;
    11'b00110110010: data <= 32'h32fac14b;
    11'b00110110011: data <= 32'h38cdbe5a;
    11'b00110110100: data <= 32'h292d3af9;
    11'b00110110101: data <= 32'hbc444015;
    11'b00110110110: data <= 32'hbd5e3c17;
    11'b00110110111: data <= 32'hb9cfb537;
    11'b00110111000: data <= 32'hb92bb565;
    11'b00110111001: data <= 32'hbdea3552;
    11'b00110111010: data <= 32'hbe36359d;
    11'b00110111011: data <= 32'h345ca02a;
    11'b00110111100: data <= 32'h40c13596;
    11'b00110111101: data <= 32'h40ae3cce;
    11'b00110111110: data <= 32'h36163d54;
    11'b00110111111: data <= 32'hbb6a3934;
    11'b00111000000: data <= 32'hb49a3498;
    11'b00111000001: data <= 32'h3a80371b;
    11'b00111000010: data <= 32'h39d0b002;
    11'b00111000011: data <= 32'h2931bf2b;
    11'b00111000100: data <= 32'h323dc18b;
    11'b00111000101: data <= 32'h3bd6be0b;
    11'b00111000110: data <= 32'h3c0539d5;
    11'b00111000111: data <= 32'h2b543d54;
    11'b00111001000: data <= 32'hb9c8aa08;
    11'b00111001001: data <= 32'hbb41bca4;
    11'b00111001010: data <= 32'hbd3eb896;
    11'b00111001011: data <= 32'hc0213714;
    11'b00111001100: data <= 32'hbf5d3312;
    11'b00111001101: data <= 32'ha5bbb946;
    11'b00111001110: data <= 32'h3eb6b7ac;
    11'b00111001111: data <= 32'h3d2c3ac1;
    11'b00111010000: data <= 32'hb78f3f24;
    11'b00111010001: data <= 32'hbc803e90;
    11'b00111010010: data <= 32'h28813ce0;
    11'b00111010011: data <= 32'h3c3d3bd9;
    11'b00111010100: data <= 32'h37c83290;
    11'b00111010101: data <= 32'hb760bd09;
    11'b00111010110: data <= 32'h2c8dbfd5;
    11'b00111010111: data <= 32'h3e87baac;
    11'b00111011000: data <= 32'h40663a32;
    11'b00111011001: data <= 32'h3cae3a06;
    11'b00111011010: data <= 32'haf74b994;
    11'b00111011011: data <= 32'hb992bd65;
    11'b00111011100: data <= 32'hbc54b5dd;
    11'b00111011101: data <= 32'hbe823721;
    11'b00111011110: data <= 32'hbdebb778;
    11'b00111011111: data <= 32'hb268bf8d;
    11'b00111100000: data <= 32'h3afcbe6a;
    11'b00111100001: data <= 32'h354a3561;
    11'b00111100010: data <= 32'hbc013f5d;
    11'b00111100011: data <= 32'hbc7e3f41;
    11'b00111100100: data <= 32'h2b6d3cda;
    11'b00111100101: data <= 32'h384b3bb9;
    11'b00111100110: data <= 32'hb89438c6;
    11'b00111100111: data <= 32'hbdc9b515;
    11'b00111101000: data <= 32'hb3a9bac6;
    11'b00111101001: data <= 32'h400db08d;
    11'b00111101010: data <= 32'h41a03aae;
    11'b00111101011: data <= 32'h3e4d38a6;
    11'b00111101100: data <= 32'h3073b7fb;
    11'b00111101101: data <= 32'hb260b911;
    11'b00111101110: data <= 32'hb09435d7;
    11'b00111101111: data <= 32'hb864384f;
    11'b00111110000: data <= 32'hba9bbc9e;
    11'b00111110001: data <= 32'hb3b6c1c2;
    11'b00111110010: data <= 32'h3738c0ad;
    11'b00111110011: data <= 32'h3023ab7b;
    11'b00111110100: data <= 32'hb9aa3da6;
    11'b00111110101: data <= 32'hb9913c3b;
    11'b00111110110: data <= 32'ha60b355b;
    11'b00111110111: data <= 32'hb4f43803;
    11'b00111111000: data <= 32'hbf1e3ae1;
    11'b00111111001: data <= 32'hc0bc3697;
    11'b00111111010: data <= 32'hb913b415;
    11'b00111111011: data <= 32'h3f55aa96;
    11'b00111111100: data <= 32'h40d6394e;
    11'b00111111101: data <= 32'h3c2239f3;
    11'b00111111110: data <= 32'hac023556;
    11'b00111111111: data <= 32'h34ed3895;
    11'b01000000000: data <= 32'h3afb3d29;
    11'b01000000001: data <= 32'h35b63a81;
    11'b01000000010: data <= 32'hb799bd32;
    11'b01000000011: data <= 32'hb4c2c1e9;
    11'b01000000100: data <= 32'h386bc06d;
    11'b01000000101: data <= 32'h3a42af92;
    11'b01000000110: data <= 32'h34d639f6;
    11'b01000000111: data <= 32'h2bceafbe;
    11'b01000001000: data <= 32'h2903ba01;
    11'b01000001001: data <= 32'hba6f29b7;
    11'b01000001010: data <= 32'hc0a33bca;
    11'b01000001011: data <= 32'hc14e384a;
    11'b01000001100: data <= 32'hbb2fb8ba;
    11'b01000001101: data <= 32'h3c9bb9fc;
    11'b01000001110: data <= 32'h3d1a316d;
    11'b01000001111: data <= 32'ha9f03b66;
    11'b01000010000: data <= 32'hb7a93c7b;
    11'b01000010001: data <= 32'h38e43dd7;
    11'b01000010010: data <= 32'h3d663f79;
    11'b01000010011: data <= 32'h36e93cad;
    11'b01000010100: data <= 32'hba96ba0d;
    11'b01000010101: data <= 32'hb85bc01d;
    11'b01000010110: data <= 32'h3b57bd5c;
    11'b01000010111: data <= 32'h3efd303f;
    11'b01000011000: data <= 32'h3d793267;
    11'b01000011001: data <= 32'h3a00bbd4;
    11'b01000011010: data <= 32'h3558bd03;
    11'b01000011011: data <= 32'hb8432ce2;
    11'b01000011100: data <= 32'hbf3d3c50;
    11'b01000011101: data <= 32'hc0433070;
    11'b01000011110: data <= 32'hbb27be45;
    11'b01000011111: data <= 32'h3632bf47;
    11'b01000100000: data <= 32'h2ff2b741;
    11'b01000100001: data <= 32'hbb173abb;
    11'b01000100010: data <= 32'hb9633cdf;
    11'b01000100011: data <= 32'h39af3d96;
    11'b01000100100: data <= 32'h3c723ef4;
    11'b01000100101: data <= 32'hb5bf3da8;
    11'b01000100110: data <= 32'hbefa30b0;
    11'b01000100111: data <= 32'hbbedba31;
    11'b01000101000: data <= 32'h3c80b57f;
    11'b01000101001: data <= 32'h40803687;
    11'b01000101010: data <= 32'h3eeca576;
    11'b01000101011: data <= 32'h3b8abc3b;
    11'b01000101100: data <= 32'h39ddba8f;
    11'b01000101101: data <= 32'h360d39d0;
    11'b01000101110: data <= 32'hb8a23d44;
    11'b01000101111: data <= 32'hbcbfb544;
    11'b01000110000: data <= 32'hb9a9c0d8;
    11'b01000110001: data <= 32'hab99c10b;
    11'b01000110010: data <= 32'hb584bab2;
    11'b01000110011: data <= 32'hbb23374c;
    11'b01000110100: data <= 32'hb597378b;
    11'b01000110101: data <= 32'h3a2d3630;
    11'b01000110110: data <= 32'h38133c0a;
    11'b01000110111: data <= 32'hbd9e3dcd;
    11'b01000111000: data <= 32'hc1493b0a;
    11'b01000111001: data <= 32'hbdb02cb7;
    11'b01000111010: data <= 32'h3b602c08;
    11'b01000111011: data <= 32'h3f6035e6;
    11'b01000111100: data <= 32'h3c4f206b;
    11'b01000111101: data <= 32'h3819b7ca;
    11'b01000111110: data <= 32'h3c1c3276;
    11'b01000111111: data <= 32'h3d8a3e8a;
    11'b01001000000: data <= 32'h388d3eac;
    11'b01001000001: data <= 32'hb810b692;
    11'b01001000010: data <= 32'hb8cdc0ed;
    11'b01001000011: data <= 32'hac91c09e;
    11'b01001000100: data <= 32'h287db9b1;
    11'b01001000101: data <= 32'hadcba6d5;
    11'b01001000110: data <= 32'h3633b98f;
    11'b01001000111: data <= 32'h3b92bb6a;
    11'b01001001000: data <= 32'h2ff8330d;
    11'b01001001001: data <= 32'hbf8e3d7e;
    11'b01001001010: data <= 32'hc1ba3c60;
    11'b01001001011: data <= 32'hbe342472;
    11'b01001001100: data <= 32'h3634b65c;
    11'b01001001101: data <= 32'h39aeadda;
    11'b01001001110: data <= 32'hb2e02b21;
    11'b01001001111: data <= 32'hb37330cb;
    11'b01001010000: data <= 32'h3c7b3c0f;
    11'b01001010001: data <= 32'h3fb7405a;
    11'b01001010010: data <= 32'h3b673fc6;
    11'b01001010011: data <= 32'hb8bb26d3;
    11'b01001010100: data <= 32'hba52be44;
    11'b01001010101: data <= 32'h30d3bcf7;
    11'b01001010110: data <= 32'h3a86b0ab;
    11'b01001010111: data <= 32'h3b0cb5a6;
    11'b01001011000: data <= 32'h3c3fbe69;
    11'b01001011001: data <= 32'h3cddbed8;
    11'b01001011010: data <= 32'h3564a90d;
    11'b01001011011: data <= 32'hbd803d8f;
    11'b01001011100: data <= 32'hc0593ab1;
    11'b01001011101: data <= 32'hbd07b9fb;
    11'b01001011110: data <= 32'hb120bd66;
    11'b01001011111: data <= 32'hb7afb9b6;
    11'b01001100000: data <= 32'hbd59aacc;
    11'b01001100001: data <= 32'hb9f13422;
    11'b01001100010: data <= 32'h3c673b86;
    11'b01001100011: data <= 32'h3f493fa3;
    11'b01001100100: data <= 32'h35e23fbf;
    11'b01001100101: data <= 32'hbd7839d0;
    11'b01001100110: data <= 32'hbcf5b40b;
    11'b01001100111: data <= 32'h34ac2884;
    11'b01001101000: data <= 32'h3d23376f;
    11'b01001101001: data <= 32'h3ce4b6cf;
    11'b01001101010: data <= 32'h3c9dbf34;
    11'b01001101011: data <= 32'h3da4be1e;
    11'b01001101100: data <= 32'h3c4636fa;
    11'b01001101101: data <= 32'hafaf3e7f;
    11'b01001101110: data <= 32'hbbaa376c;
    11'b01001101111: data <= 32'hb9c9be1b;
    11'b01001110000: data <= 32'hb6ecc00b;
    11'b01001110001: data <= 32'hbc3abc21;
    11'b01001110010: data <= 32'hbe74b49f;
    11'b01001110011: data <= 32'hb905b575;
    11'b01001110100: data <= 32'h3c92adbd;
    11'b01001110101: data <= 32'h3d553b6b;
    11'b01001110110: data <= 32'hb88d3e81;
    11'b01001110111: data <= 32'hc0723d11;
    11'b01001111000: data <= 32'hbe8b3988;
    11'b01001111001: data <= 32'h31de39d9;
    11'b01001111010: data <= 32'h3be5395f;
    11'b01001111011: data <= 32'h386bb5a6;
    11'b01001111100: data <= 32'h37f4bd6b;
    11'b01001111101: data <= 32'h3d80b930;
    11'b01001111110: data <= 32'h3f7f3d25;
    11'b01001111111: data <= 32'h3c753fdd;
    11'b01010000000: data <= 32'h26713567;
    11'b01010000001: data <= 32'hb54fbe8f;
    11'b01010000010: data <= 32'hb5f6bf2d;
    11'b01010000011: data <= 32'hba77b9b7;
    11'b01010000100: data <= 32'hbbe0b78a;
    11'b01010000101: data <= 32'h27a7bd3e;
    11'b01010000110: data <= 32'h3d4abdec;
    11'b01010000111: data <= 32'h3b94b196;
    11'b01010001000: data <= 32'hbc5c3ced;
    11'b01010001001: data <= 32'hc0de3d83;
    11'b01010001010: data <= 32'hbe703a24;
    11'b01010001011: data <= 32'hadbe37a1;
    11'b01010001100: data <= 32'h288f3524;
    11'b01010001101: data <= 32'hba7cb511;
    11'b01010001110: data <= 32'hb879ba0a;
    11'b01010001111: data <= 32'h3c84316a;
    11'b01010010000: data <= 32'h40933f48;
    11'b01010010001: data <= 32'h3e684041;
    11'b01010010010: data <= 32'h31c83879;
    11'b01010010011: data <= 32'hb5f5bb40;
    11'b01010010100: data <= 32'hb0f0b94d;
    11'b01010010101: data <= 32'hae1530e5;
    11'b01010010110: data <= 32'ha965b734;
    11'b01010010111: data <= 32'h3998c022;
    11'b01010011000: data <= 32'h3e12c0c9;
    11'b01010011001: data <= 32'h3beeb9a1;
    11'b01010011010: data <= 32'hb9c03c39;
    11'b01010011011: data <= 32'hbec33c6d;
    11'b01010011100: data <= 32'hbc212de9;
    11'b01010011101: data <= 32'hb4b2b694;
    11'b01010011110: data <= 32'hbbf2b4a3;
    11'b01010011111: data <= 32'hc01fb633;
    11'b01010100000: data <= 32'hbd76b837;
    11'b01010100001: data <= 32'h3aff32e0;
    11'b01010100010: data <= 32'h40493e11;
    11'b01010100011: data <= 32'h3c993f77;
    11'b01010100100: data <= 32'hb7e43b70;
    11'b01010100101: data <= 32'hba5833bb;
    11'b01010100110: data <= 32'h0d6539ed;
    11'b01010100111: data <= 32'h37283c54;
    11'b01010101000: data <= 32'h3654b401;
    11'b01010101001: data <= 32'h3a2ec068;
    11'b01010101010: data <= 32'h3e00c0a9;
    11'b01010101011: data <= 32'h3dadb5e8;
    11'b01010101100: data <= 32'h35f13cf0;
    11'b01010101101: data <= 32'hb5a139dd;
    11'b01010101110: data <= 32'hb14eb9c3;
    11'b01010101111: data <= 32'hb431bc9c;
    11'b01010110000: data <= 32'hbdf3b8d6;
    11'b01010110001: data <= 32'hc0f0b747;
    11'b01010110010: data <= 32'hbdbabadf;
    11'b01010110011: data <= 32'h3a9db93e;
    11'b01010110100: data <= 32'h3e9e36c6;
    11'b01010110101: data <= 32'h32ca3ce1;
    11'b01010110110: data <= 32'hbd903c93;
    11'b01010110111: data <= 32'hbcc93c58;
    11'b01010111000: data <= 32'h24363e55;
    11'b01010111001: data <= 32'h36063e0e;
    11'b01010111010: data <= 32'hafe7aa13;
    11'b01010111011: data <= 32'h256fbf04;
    11'b01010111100: data <= 32'h3c8fbde8;
    11'b01010111101: data <= 32'h3f8e37e4;
    11'b01010111110: data <= 32'h3df83e58;
    11'b01010111111: data <= 32'h3a503827;
    11'b01011000000: data <= 32'h37e6bc14;
    11'b01011000001: data <= 32'ha71bbc43;
    11'b01011000010: data <= 32'hbce6b2d8;
    11'b01011000011: data <= 32'hbf95b569;
    11'b01011000100: data <= 32'hba60bdfc;
    11'b01011000101: data <= 32'h3c0abfb1;
    11'b01011000110: data <= 32'h3cd8babe;
    11'b01011000111: data <= 32'hb753382a;
    11'b01011001000: data <= 32'hbeec3c24;
    11'b01011001001: data <= 32'hbc7b3c89;
    11'b01011001010: data <= 32'h20663da6;
    11'b01011001011: data <= 32'hb41e3cea;
    11'b01011001100: data <= 32'hbd6e11d5;
    11'b01011001101: data <= 32'hbccbbc79;
    11'b01011001110: data <= 32'h3882b85e;
    11'b01011001111: data <= 32'h40163c95;
    11'b01011010000: data <= 32'h3fbe3ee2;
    11'b01011010001: data <= 32'h3c3a381b;
    11'b01011010010: data <= 32'h388ab8a6;
    11'b01011010011: data <= 32'h335fac2a;
    11'b01011010100: data <= 32'hb7d83a7d;
    11'b01011010101: data <= 32'hbafe2693;
    11'b01011010110: data <= 32'ha61ebfdf;
    11'b01011010111: data <= 32'h3ccfc18f;
    11'b01011011000: data <= 32'h3c45be0b;
    11'b01011011001: data <= 32'hb5b531b4;
    11'b01011011010: data <= 32'hbc7c397f;
    11'b01011011011: data <= 32'hb6653719;
    11'b01011011100: data <= 32'h30b537b2;
    11'b01011011101: data <= 32'hbbe1384c;
    11'b01011011110: data <= 32'hc115ad41;
    11'b01011011111: data <= 32'hc055b9f1;
    11'b01011100000: data <= 32'h2ddeb419;
    11'b01011100001: data <= 32'h3f1f3bda;
    11'b01011100010: data <= 32'h3ddf3d5b;
    11'b01011100011: data <= 32'h3602386c;
    11'b01011100100: data <= 32'h2e563423;
    11'b01011100101: data <= 32'h35e53d11;
    11'b01011100110: data <= 32'h31473faf;
    11'b01011100111: data <= 32'hb31337cd;
    11'b01011101000: data <= 32'h3233bfc7;
    11'b01011101001: data <= 32'h3c5ec165;
    11'b01011101010: data <= 32'h3cc0bcd1;
    11'b01011101011: data <= 32'h36cf35cf;
    11'b01011101100: data <= 32'h306d3523;
    11'b01011101101: data <= 32'h3949b743;
    11'b01011101110: data <= 32'h37a6b720;
    11'b01011101111: data <= 32'hbd222cdf;
    11'b01011110000: data <= 32'hc1dcadb9;
    11'b01011110001: data <= 32'hc099ba61;
    11'b01011110010: data <= 32'h18afba98;
    11'b01011110011: data <= 32'h3d1fa5f6;
    11'b01011110100: data <= 32'h376f37f2;
    11'b01011110101: data <= 32'hb969370d;
    11'b01011110110: data <= 32'hb7203b05;
    11'b01011110111: data <= 32'h36a6402d;
    11'b01011111000: data <= 32'h355e40ea;
    11'b01011111001: data <= 32'hb72e3a46;
    11'b01011111010: data <= 32'hb747bdd2;
    11'b01011111011: data <= 32'h385fbf2a;
    11'b01011111100: data <= 32'h3d44b307;
    11'b01011111101: data <= 32'h3d2f3abb;
    11'b01011111110: data <= 32'h3d082e36;
    11'b01011111111: data <= 32'h3ddcbbae;
    11'b01100000000: data <= 32'h3ae4b914;
    11'b01100000001: data <= 32'hbb9a3596;
    11'b01100000010: data <= 32'hc0a1321f;
    11'b01100000011: data <= 32'hbe4fbc61;
    11'b01100000100: data <= 32'h34a8bf4c;
    11'b01100000101: data <= 32'h3ab3bd0f;
    11'b01100000110: data <= 32'hb61db617;
    11'b01100000111: data <= 32'hbd1b3024;
    11'b01100001000: data <= 32'hb8033a93;
    11'b01100001001: data <= 32'h38593f8f;
    11'b01100001010: data <= 32'h274e4042;
    11'b01100001011: data <= 32'hbd9f3a14;
    11'b01100001100: data <= 32'hbe92ba96;
    11'b01100001101: data <= 32'hb361b9ab;
    11'b01100001110: data <= 32'h3ce3396c;
    11'b01100001111: data <= 32'h3e693c7c;
    11'b01100010000: data <= 32'h3e0ba365;
    11'b01100010001: data <= 32'h3e2cbaa2;
    11'b01100010010: data <= 32'h3c5c2d65;
    11'b01100010011: data <= 32'hb2d23d53;
    11'b01100010100: data <= 32'hbcaa3a20;
    11'b01100010101: data <= 32'hb8a3bd20;
    11'b01100010110: data <= 32'h3919c107;
    11'b01100010111: data <= 32'h38f2bfb5;
    11'b01100011000: data <= 32'hb888ba3a;
    11'b01100011001: data <= 32'hbb9cb3c6;
    11'b01100011010: data <= 32'h312d2f3d;
    11'b01100011011: data <= 32'h3b223ad4;
    11'b01100011100: data <= 32'hb6433cf5;
    11'b01100011101: data <= 32'hc0cc382d;
    11'b01100011110: data <= 32'hc13ab65c;
    11'b01100011111: data <= 32'hba73b0fe;
    11'b01100100000: data <= 32'h3b043a65;
    11'b01100100001: data <= 32'h3c603a89;
    11'b01100100010: data <= 32'h39f9b18a;
    11'b01100100011: data <= 32'h3b4eb4ef;
    11'b01100100100: data <= 32'h3c563cd5;
    11'b01100100101: data <= 32'h378b40e7;
    11'b01100100110: data <= 32'hb4613d7e;
    11'b01100100111: data <= 32'hacbcbc7e;
    11'b01100101000: data <= 32'h3907c0bb;
    11'b01100101001: data <= 32'h387abe3e;
    11'b01100101010: data <= 32'haed8b7a0;
    11'b01100101011: data <= 32'h2d72b7d9;
    11'b01100101100: data <= 32'h3cefba6d;
    11'b01100101101: data <= 32'h3d9cb49c;
    11'b01100101110: data <= 32'hb81137e3;
    11'b01100101111: data <= 32'hc1653632;
    11'b01100110000: data <= 32'hc16ab4cf;
    11'b01100110001: data <= 32'hbaa1b678;
    11'b01100110010: data <= 32'h37552872;
    11'b01100110011: data <= 32'h2ca2a7e7;
    11'b01100110100: data <= 32'hb7f5b7d8;
    11'b01100110101: data <= 32'h2e032da7;
    11'b01100110110: data <= 32'h3be13fae;
    11'b01100110111: data <= 32'h3a1c41f2;
    11'b01100111000: data <= 32'hb2173ea0;
    11'b01100111001: data <= 32'hb771b95d;
    11'b01100111010: data <= 32'h2dffbdbd;
    11'b01100111011: data <= 32'h378cb683;
    11'b01100111100: data <= 32'h38123420;
    11'b01100111101: data <= 32'h3c50b878;
    11'b01100111110: data <= 32'h4018bd9e;
    11'b01100111111: data <= 32'h3f50ba36;
    11'b01101000000: data <= 32'hb13d37e0;
    11'b01101000001: data <= 32'hc0193910;
    11'b01101000010: data <= 32'hbf5fb622;
    11'b01101000011: data <= 32'hb4fabc80;
    11'b01101000100: data <= 32'h316cbc3e;
    11'b01101000101: data <= 32'hbacdbb7e;
    11'b01101000110: data <= 32'hbd89bb2c;
    11'b01101000111: data <= 32'hb3fba72a;
    11'b01101001000: data <= 32'h3c333eb6;
    11'b01101001001: data <= 32'h3944410f;
    11'b01101001010: data <= 32'hbad33dc3;
    11'b01101001011: data <= 32'hbdf3b1be;
    11'b01101001100: data <= 32'hb9c5b49d;
    11'b01101001101: data <= 32'h338f3a1b;
    11'b01101001110: data <= 32'h39a73aae;
    11'b01101001111: data <= 32'h3d1bb8a1;
    11'b01101010000: data <= 32'h4018bdd4;
    11'b01101010001: data <= 32'h3fa7b5c3;
    11'b01101010010: data <= 32'h374d3d26;
    11'b01101010011: data <= 32'hbac23cfa;
    11'b01101010100: data <= 32'hb8b1b651;
    11'b01101010101: data <= 32'h3563bea6;
    11'b01101010110: data <= 32'h2c32bea2;
    11'b01101010111: data <= 32'hbccbbd2b;
    11'b01101011000: data <= 32'hbd76bcba;
    11'b01101011001: data <= 32'h3284b938;
    11'b01101011010: data <= 32'h3db238bb;
    11'b01101011011: data <= 32'h36ef3d9c;
    11'b01101011100: data <= 32'hbea23b3d;
    11'b01101011101: data <= 32'hc0c32f2c;
    11'b01101011110: data <= 32'hbd28368c;
    11'b01101011111: data <= 32'had2d3ccb;
    11'b01101100000: data <= 32'h33b83a21;
    11'b01101100001: data <= 32'h3772b9f5;
    11'b01101100010: data <= 32'h3cd4bc8f;
    11'b01101100011: data <= 32'h3e813861;
    11'b01101100100: data <= 32'h3bfa40a2;
    11'b01101100101: data <= 32'h31a33f7d;
    11'b01101100110: data <= 32'h3394b2a9;
    11'b01101100111: data <= 32'h38babe0f;
    11'b01101101000: data <= 32'h2635bcfb;
    11'b01101101001: data <= 32'hbb8eba89;
    11'b01101101010: data <= 32'hb88ebcb8;
    11'b01101101011: data <= 32'h3caebdb5;
    11'b01101101100: data <= 32'h3fe6b94f;
    11'b01101101101: data <= 32'h364f356d;
    11'b01101101110: data <= 32'hbfaa37b7;
    11'b01101101111: data <= 32'hc0dc3131;
    11'b01101110000: data <= 32'hbcb535ce;
    11'b01101110001: data <= 32'hb4b13992;
    11'b01101110010: data <= 32'hb938298c;
    11'b01101110011: data <= 32'hbb0bbc74;
    11'b01101110100: data <= 32'h2d02bae5;
    11'b01101110101: data <= 32'h3ce23cba;
    11'b01101110110: data <= 32'h3cda4197;
    11'b01101110111: data <= 32'h373f4020;
    11'b01101111000: data <= 32'h302f2da7;
    11'b01101111001: data <= 32'h32b3b980;
    11'b01101111010: data <= 32'haf5b0ed0;
    11'b01101111011: data <= 32'hb7ab32cc;
    11'b01101111100: data <= 32'h3503bb7b;
    11'b01101111101: data <= 32'h3fc4bfb7;
    11'b01101111110: data <= 32'h40b3bd56;
    11'b01101111111: data <= 32'h39172841;
    11'b01110000000: data <= 32'hbd603852;
    11'b01110000001: data <= 32'hbdec2f9a;
    11'b01110000010: data <= 32'hb633b1e6;
    11'b01110000011: data <= 32'hb46db41d;
    11'b01110000100: data <= 32'hbdd9ba8d;
    11'b01110000101: data <= 32'hbfc1be0a;
    11'b01110000110: data <= 32'hb8b1bb71;
    11'b01110000111: data <= 32'h3c3f3be8;
    11'b01110001000: data <= 32'h3c80408f;
    11'b01110001001: data <= 32'ha5aa3e6c;
    11'b01110001010: data <= 32'hb9bc34b0;
    11'b01110001011: data <= 32'hb86b3578;
    11'b01110001100: data <= 32'hb5fc3d57;
    11'b01110001101: data <= 32'hb4923c7e;
    11'b01110001110: data <= 32'h383fb999;
    11'b01110001111: data <= 32'h3f8abfe4;
    11'b01110010000: data <= 32'h4078bc73;
    11'b01110010001: data <= 32'h3bff38fa;
    11'b01110010010: data <= 32'hb40b3c50;
    11'b01110010011: data <= 32'hac4430d6;
    11'b01110010100: data <= 32'h38cfb95c;
    11'b01110010101: data <= 32'hae4cbac1;
    11'b01110010110: data <= 32'hbf1dbc89;
    11'b01110010111: data <= 32'hc03dbe92;
    11'b01110011000: data <= 32'hb5eebd5a;
    11'b01110011001: data <= 32'h3d581eca;
    11'b01110011010: data <= 32'h3b9c3c05;
    11'b01110011011: data <= 32'hb9e939d8;
    11'b01110011100: data <= 32'hbe48348b;
    11'b01110011101: data <= 32'hbc5e3be7;
    11'b01110011110: data <= 32'hb8b53fe4;
    11'b01110011111: data <= 32'hb8a83d4a;
    11'b01110100000: data <= 32'hb208b9de;
    11'b01110100001: data <= 32'h3b51bed1;
    11'b01110100010: data <= 32'h3e7db528;
    11'b01110100011: data <= 32'h3ced3e54;
    11'b01110100100: data <= 32'h399b3ebe;
    11'b01110100101: data <= 32'h3bb5347e;
    11'b01110100110: data <= 32'h3c9fb920;
    11'b01110100111: data <= 32'h2778b80c;
    11'b01110101000: data <= 32'hbe40b863;
    11'b01110101001: data <= 32'hbddbbd5e;
    11'b01110101010: data <= 32'h37f2bf3d;
    11'b01110101011: data <= 32'h3f76bcae;
    11'b01110101100: data <= 32'h3b25b446;
    11'b01110101101: data <= 32'hbc45a5ca;
    11'b01110101110: data <= 32'hbeb3300f;
    11'b01110101111: data <= 32'hbb263bba;
    11'b01110110000: data <= 32'hb8533e89;
    11'b01110110001: data <= 32'hbcc539de;
    11'b01110110010: data <= 32'hbdcebc48;
    11'b01110110011: data <= 32'hb6b7bdbd;
    11'b01110110100: data <= 32'h3aeb3574;
    11'b01110110101: data <= 32'h3cd14032;
    11'b01110110110: data <= 32'h3be23f40;
    11'b01110110111: data <= 32'h3c2a35cc;
    11'b01110111000: data <= 32'h3b93ac43;
    11'b01110111001: data <= 32'haba43943;
    11'b01110111010: data <= 32'hbc81396b;
    11'b01110111011: data <= 32'hb8b9b9e6;
    11'b01110111100: data <= 32'h3d28c014;
    11'b01110111101: data <= 32'h4066bf54;
    11'b01110111110: data <= 32'h3bbcba35;
    11'b01110111111: data <= 32'hb9b3b1c9;
    11'b01111000000: data <= 32'hba6f1ae0;
    11'b01111000001: data <= 32'h2d003752;
    11'b01111000010: data <= 32'hb16539cd;
    11'b01111000011: data <= 32'hbedeb025;
    11'b01111000100: data <= 32'hc0f9bdca;
    11'b01111000101: data <= 32'hbd37bd86;
    11'b01111000110: data <= 32'h3722353c;
    11'b01111000111: data <= 32'h3bff3ea2;
    11'b01111001000: data <= 32'h38683cc7;
    11'b01111001001: data <= 32'h345e334c;
    11'b01111001010: data <= 32'h32c73965;
    11'b01111001011: data <= 32'hb4f83fd9;
    11'b01111001100: data <= 32'hbad63f47;
    11'b01111001101: data <= 32'hb358b27b;
    11'b01111001110: data <= 32'h3d38bfb6;
    11'b01111001111: data <= 32'h3fcebe95;
    11'b01111010000: data <= 32'h3c13b4c9;
    11'b01111010001: data <= 32'h2e3a34ba;
    11'b01111010010: data <= 32'h389726fd;
    11'b01111010011: data <= 32'h3d3aac6e;
    11'b01111010100: data <= 32'h35732827;
    11'b01111010101: data <= 32'hbf5db820;
    11'b01111010110: data <= 32'hc164bdea;
    11'b01111010111: data <= 32'hbcecbe0e;
    11'b01111011000: data <= 32'h38ecb630;
    11'b01111011001: data <= 32'h3a6f36c8;
    11'b01111011010: data <= 32'hb1c32cf3;
    11'b01111011011: data <= 32'hb930b04d;
    11'b01111011100: data <= 32'hb6463c66;
    11'b01111011101: data <= 32'hb752413f;
    11'b01111011110: data <= 32'hbb5c4063;
    11'b01111011111: data <= 32'hb99cad7c;
    11'b01111100000: data <= 32'h361ebe75;
    11'b01111100001: data <= 32'h3c6cbadf;
    11'b01111100010: data <= 32'h3b17398b;
    11'b01111100011: data <= 32'h3a793b9f;
    11'b01111100100: data <= 32'h3e802f85;
    11'b01111100101: data <= 32'h4022b335;
    11'b01111100110: data <= 32'h395630bc;
    11'b01111100111: data <= 32'hbe3522b0;
    11'b01111101000: data <= 32'hc01cbbba;
    11'b01111101001: data <= 32'hb5dbbe80;
    11'b01111101010: data <= 32'h3cb3bd3c;
    11'b01111101011: data <= 32'h39ccbaee;
    11'b01111101100: data <= 32'hb936bb49;
    11'b01111101101: data <= 32'hbb97b84f;
    11'b01111101110: data <= 32'hb4283bc8;
    11'b01111101111: data <= 32'hb34a409d;
    11'b01111110000: data <= 32'hbcc03e93;
    11'b01111110001: data <= 32'hbed0b6cf;
    11'b01111110010: data <= 32'hbbb8bd54;
    11'b01111110011: data <= 32'h2dd8ad9d;
    11'b01111110100: data <= 32'h388b3d84;
    11'b01111110101: data <= 32'h3ba73c9e;
    11'b01111110110: data <= 32'h3ef22a90;
    11'b01111110111: data <= 32'h3fc2285e;
    11'b01111111000: data <= 32'h38e53c37;
    11'b01111111001: data <= 32'hbc673cf9;
    11'b01111111010: data <= 32'hbc6aae0f;
    11'b01111111011: data <= 32'h388cbe1f;
    11'b01111111100: data <= 32'h3e5cbf36;
    11'b01111111101: data <= 32'h397bbdaa;
    11'b01111111110: data <= 32'hb89fbcc8;
    11'b01111111111: data <= 32'hb53bb9f0;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    