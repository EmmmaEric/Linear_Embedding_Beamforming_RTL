
module memory_rom_25(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3cefbbf8;
    11'b00000000001: data <= 32'h392ab8a4;
    11'b00000000010: data <= 32'hba3b3887;
    11'b00000000011: data <= 32'hbf5c35b2;
    11'b00000000100: data <= 32'hbca8bd1f;
    11'b00000000101: data <= 32'h36f4c0a4;
    11'b00000000110: data <= 32'h3a4dbe8f;
    11'b00000000111: data <= 32'hb758b515;
    11'b00000001000: data <= 32'hbd2b368c;
    11'b00000001001: data <= 32'hb7573a88;
    11'b00000001010: data <= 32'h386c3dcf;
    11'b00000001011: data <= 32'hb0d93e8f;
    11'b00000001100: data <= 32'hbf493913;
    11'b00000001101: data <= 32'hc021b8cb;
    11'b00000001110: data <= 32'hb538b761;
    11'b00000001111: data <= 32'h3de13a03;
    11'b00000010000: data <= 32'h3f2a3c75;
    11'b00000010001: data <= 32'h3d242cc0;
    11'b00000010010: data <= 32'h3c4fb8a3;
    11'b00000010011: data <= 32'h3b283702;
    11'b00000010100: data <= 32'h2d2d3e9a;
    11'b00000010101: data <= 32'hb9993af0;
    11'b00000010110: data <= 32'hb5b2bde2;
    11'b00000010111: data <= 32'h38d4c195;
    11'b00000011000: data <= 32'h3919bfcd;
    11'b00000011001: data <= 32'hb4f5b7c2;
    11'b00000011010: data <= 32'hb8bb9f31;
    11'b00000011011: data <= 32'h3617ae68;
    11'b00000011100: data <= 32'h3adf34ae;
    11'b00000011101: data <= 32'hb9033a91;
    11'b00000011110: data <= 32'hc160381d;
    11'b00000011111: data <= 32'hc186b40b;
    11'b00000100000: data <= 32'hb9b2b3f8;
    11'b00000100001: data <= 32'h3c2e377f;
    11'b00000100010: data <= 32'h3bfc38d4;
    11'b00000100011: data <= 32'h347ca6dc;
    11'b00000100100: data <= 32'h36972d0e;
    11'b00000100101: data <= 32'h3bbc3e38;
    11'b00000100110: data <= 32'h39b74132;
    11'b00000100111: data <= 32'hae7e3d5e;
    11'b00000101000: data <= 32'hb373bcd0;
    11'b00000101001: data <= 32'h3659c09f;
    11'b00000101010: data <= 32'h396abd0d;
    11'b00000101011: data <= 32'h362eacd3;
    11'b00000101100: data <= 32'h388eb528;
    11'b00000101101: data <= 32'h3d8dbc1f;
    11'b00000101110: data <= 32'h3d23b932;
    11'b00000101111: data <= 32'hb9083635;
    11'b00000110000: data <= 32'hc14d3854;
    11'b00000110001: data <= 32'hc103b4c9;
    11'b00000110010: data <= 32'hb8c9ba99;
    11'b00000110011: data <= 32'h384cb851;
    11'b00000110100: data <= 32'hb020b454;
    11'b00000110101: data <= 32'hbb1db47b;
    11'b00000110110: data <= 32'hb2273659;
    11'b00000110111: data <= 32'h3bd93fe6;
    11'b00000111000: data <= 32'h3aaa4195;
    11'b00000111001: data <= 32'hb6713e01;
    11'b00000111010: data <= 32'hbb9eb8ec;
    11'b00000111011: data <= 32'hb32dbcb0;
    11'b00000111100: data <= 32'h3951aaac;
    11'b00000111101: data <= 32'h3c01385f;
    11'b00000111110: data <= 32'h3d71b76c;
    11'b00000111111: data <= 32'h3fbabdd5;
    11'b00001000000: data <= 32'h3e7cb9f7;
    11'b00001000001: data <= 32'hae3b39fe;
    11'b00001000010: data <= 32'hbecc3b2a;
    11'b00001000011: data <= 32'hbde0b7f9;
    11'b00001000100: data <= 32'haf1cbe9d;
    11'b00001000101: data <= 32'h320abe3c;
    11'b00001000110: data <= 32'hbb58bbee;
    11'b00001000111: data <= 32'hbdb5b915;
    11'b00001001000: data <= 32'hb22c2bba;
    11'b00001001001: data <= 32'h3c8f3d77;
    11'b00001001010: data <= 32'h38704031;
    11'b00001001011: data <= 32'hbd283d12;
    11'b00001001100: data <= 32'hc010a966;
    11'b00001001101: data <= 32'hbb8bad21;
    11'b00001001110: data <= 32'h37503ade;
    11'b00001001111: data <= 32'h3be13ab8;
    11'b00001010000: data <= 32'h3cb7b853;
    11'b00001010001: data <= 32'h3e92bd1e;
    11'b00001010010: data <= 32'h3eb69c4d;
    11'b00001010011: data <= 32'h39453ede;
    11'b00001010100: data <= 32'hb6fe3dee;
    11'b00001010101: data <= 32'hb5afb856;
    11'b00001010110: data <= 32'h3548c00d;
    11'b00001010111: data <= 32'h2c53bf45;
    11'b00001011000: data <= 32'hbbf8bc48;
    11'b00001011001: data <= 32'hbc13bb45;
    11'b00001011010: data <= 32'h3813ba29;
    11'b00001011011: data <= 32'h3e1b2e55;
    11'b00001011100: data <= 32'h342b3be2;
    11'b00001011101: data <= 32'hc00c3aea;
    11'b00001011110: data <= 32'hc15a33f7;
    11'b00001011111: data <= 32'hbd24358e;
    11'b00001100000: data <= 32'h2faf3b10;
    11'b00001100001: data <= 32'h340237db;
    11'b00001100010: data <= 32'h2cfbb9bd;
    11'b00001100011: data <= 32'h39acba9d;
    11'b00001100100: data <= 32'h3ddf3b9a;
    11'b00001100101: data <= 32'h3cdd413a;
    11'b00001100110: data <= 32'h35cc3fd1;
    11'b00001100111: data <= 32'h2dc0b4e0;
    11'b00001101000: data <= 32'h350dbe4c;
    11'b00001101001: data <= 32'h29d3bc2e;
    11'b00001101010: data <= 32'hb82db6c6;
    11'b00001101011: data <= 32'haa2cbba8;
    11'b00001101100: data <= 32'h3ddabe74;
    11'b00001101101: data <= 32'h3ff2bc1f;
    11'b00001101110: data <= 32'h3482330d;
    11'b00001101111: data <= 32'hbfec3956;
    11'b00001110000: data <= 32'hc0b233b5;
    11'b00001110001: data <= 32'hbbc71a2d;
    11'b00001110010: data <= 32'hb0d02dec;
    11'b00001110011: data <= 32'hba50b51f;
    11'b00001110100: data <= 32'hbd10bc23;
    11'b00001110101: data <= 32'hb36cb8a9;
    11'b00001110110: data <= 32'h3cea3d58;
    11'b00001110111: data <= 32'h3d62417f;
    11'b00001111000: data <= 32'h34b93fd6;
    11'b00001111001: data <= 32'hb6212d64;
    11'b00001111010: data <= 32'hb324b81c;
    11'b00001111011: data <= 32'haa18353e;
    11'b00001111100: data <= 32'ha6083841;
    11'b00001111101: data <= 32'h3974ba9d;
    11'b00001111110: data <= 32'h3fdcc00e;
    11'b00001111111: data <= 32'h406fbd6f;
    11'b00010000000: data <= 32'h394734ec;
    11'b00010000001: data <= 32'hbc613b49;
    11'b00010000010: data <= 32'hbca43012;
    11'b00010000011: data <= 32'hb138b964;
    11'b00010000100: data <= 32'hb2f8bab1;
    11'b00010000101: data <= 32'hbe2ebc0c;
    11'b00010000110: data <= 32'hc011bd57;
    11'b00010000111: data <= 32'hb842ba86;
    11'b00010001000: data <= 32'h3cfa3a37;
    11'b00010001001: data <= 32'h3c943faf;
    11'b00010001010: data <= 32'hb6a03db4;
    11'b00010001011: data <= 32'hbd5e360e;
    11'b00010001100: data <= 32'hbb583845;
    11'b00010001101: data <= 32'hb3eb3dde;
    11'b00010001110: data <= 32'h21aa3c98;
    11'b00010001111: data <= 32'h3840b9cd;
    11'b00010010000: data <= 32'h3e45bfa6;
    11'b00010010001: data <= 32'h4004ba82;
    11'b00010010010: data <= 32'h3c9b3c80;
    11'b00010010011: data <= 32'h2f703de1;
    11'b00010010100: data <= 32'h31b82f2e;
    11'b00010010101: data <= 32'h38f9bc32;
    11'b00010010110: data <= 32'hb019bc6e;
    11'b00010010111: data <= 32'hbeaebc08;
    11'b00010011000: data <= 32'hbf59bd8d;
    11'b00010011001: data <= 32'ha1edbda1;
    11'b00010011010: data <= 32'h3e5cb6fd;
    11'b00010011011: data <= 32'h3b3c38ba;
    11'b00010011100: data <= 32'hbc6d3952;
    11'b00010011101: data <= 32'hbfeb36e1;
    11'b00010011110: data <= 32'hbcd03bed;
    11'b00010011111: data <= 32'hb6a53ee0;
    11'b00010100000: data <= 32'hb82b3c11;
    11'b00010100001: data <= 32'hb823bab9;
    11'b00010100010: data <= 32'h36dabe1b;
    11'b00010100011: data <= 32'h3dc32c0b;
    11'b00010100100: data <= 32'h3dcb3ffa;
    11'b00010100101: data <= 32'h3b713fa0;
    11'b00010100110: data <= 32'h3aee336a;
    11'b00010100111: data <= 32'h3ae7ba0e;
    11'b00010101000: data <= 32'hab97b61d;
    11'b00010101001: data <= 32'hbd14b1ad;
    11'b00010101010: data <= 32'hbbcfbc60;
    11'b00010101011: data <= 32'h3b24bfec;
    11'b00010101100: data <= 32'h4010be45;
    11'b00010101101: data <= 32'h3ad8b6da;
    11'b00010101110: data <= 32'hbcba318c;
    11'b00010101111: data <= 32'hbec334bb;
    11'b00010110000: data <= 32'hb9dc39c2;
    11'b00010110001: data <= 32'hb5ed3c46;
    11'b00010110010: data <= 32'hbd2f3483;
    11'b00010110011: data <= 32'hbf6abc96;
    11'b00010110100: data <= 32'hba2ebd03;
    11'b00010110101: data <= 32'h3afe3837;
    11'b00010110110: data <= 32'h3da94053;
    11'b00010110111: data <= 32'h3b703f22;
    11'b00010111000: data <= 32'h3884357a;
    11'b00010111001: data <= 32'h36f82b1f;
    11'b00010111010: data <= 32'hb07c3bd4;
    11'b00010111011: data <= 32'hba363c27;
    11'b00010111100: data <= 32'hb29ab8e4;
    11'b00010111101: data <= 32'h3db2c066;
    11'b00010111110: data <= 32'h4056bfd0;
    11'b00010111111: data <= 32'h3bfdb854;
    11'b00011000000: data <= 32'hb82c3437;
    11'b00011000001: data <= 32'hb82830f7;
    11'b00011000010: data <= 32'h35492cc5;
    11'b00011000011: data <= 32'haccc3061;
    11'b00011000100: data <= 32'hbf54b6e9;
    11'b00011000101: data <= 32'hc158bd8c;
    11'b00011000110: data <= 32'hbd33bd31;
    11'b00011000111: data <= 32'h39853163;
    11'b00011001000: data <= 32'h3ca53d6d;
    11'b00011001001: data <= 32'h344d3c0b;
    11'b00011001010: data <= 32'hb5c63465;
    11'b00011001011: data <= 32'hb4463af4;
    11'b00011001100: data <= 32'hb4ea4053;
    11'b00011001101: data <= 32'hb8d23fa0;
    11'b00011001110: data <= 32'hb1e7b441;
    11'b00011001111: data <= 32'h3c38c000;
    11'b00011010000: data <= 32'h3efabddc;
    11'b00011010001: data <= 32'h3c903293;
    11'b00011010010: data <= 32'h37353a73;
    11'b00011010011: data <= 32'h3ae62ffe;
    11'b00011010100: data <= 32'h3d8db651;
    11'b00011010101: data <= 32'h34ccb46a;
    11'b00011010110: data <= 32'hbf5fb777;
    11'b00011010111: data <= 32'hc113bd0a;
    11'b00011011000: data <= 32'hbb18be44;
    11'b00011011001: data <= 32'h3be7ba76;
    11'b00011011010: data <= 32'h3b49a1de;
    11'b00011011011: data <= 32'hb7b1a8c0;
    11'b00011011100: data <= 32'hbc6e1daf;
    11'b00011011101: data <= 32'hb8c63cbc;
    11'b00011011110: data <= 32'hb55c40f7;
    11'b00011011111: data <= 32'hbac73fae;
    11'b00011100000: data <= 32'hbc03b4b6;
    11'b00011100001: data <= 32'haf37be65;
    11'b00011100010: data <= 32'h3b16b87b;
    11'b00011100011: data <= 32'h3c5d3c9d;
    11'b00011100100: data <= 32'h3c633d28;
    11'b00011100101: data <= 32'h3e80308b;
    11'b00011100110: data <= 32'h3f44b595;
    11'b00011100111: data <= 32'h3800337a;
    11'b00011101000: data <= 32'hbda73616;
    11'b00011101001: data <= 32'hbeb0b97a;
    11'b00011101010: data <= 32'h2c15bf20;
    11'b00011101011: data <= 32'h3de3bf01;
    11'b00011101100: data <= 32'h3a54bc72;
    11'b00011101101: data <= 32'hba16ba0f;
    11'b00011101110: data <= 32'hbc13b4f4;
    11'b00011101111: data <= 32'hb0023aeb;
    11'b00011110000: data <= 32'ha7ef3f67;
    11'b00011110001: data <= 32'hbd103cb3;
    11'b00011110010: data <= 32'hc047b90d;
    11'b00011110011: data <= 32'hbd96bd1e;
    11'b00011110100: data <= 32'h2b172c83;
    11'b00011110101: data <= 32'h3a9e3e05;
    11'b00011110110: data <= 32'h3c193cba;
    11'b00011110111: data <= 32'h3d732604;
    11'b00011111000: data <= 32'h3daf2fd2;
    11'b00011111001: data <= 32'h36943d8e;
    11'b00011111010: data <= 32'hbb203eb5;
    11'b00011111011: data <= 32'hba272d89;
    11'b00011111100: data <= 32'h3a18bee7;
    11'b00011111101: data <= 32'h3e91c015;
    11'b00011111110: data <= 32'h39eabd21;
    11'b00011111111: data <= 32'hb6b7b9fc;
    11'b00100000000: data <= 32'haac1b79f;
    11'b00100000001: data <= 32'h3c0d3249;
    11'b00100000010: data <= 32'h38883a8e;
    11'b00100000011: data <= 32'hbdfc3507;
    11'b00100000100: data <= 32'hc1aebb5e;
    11'b00100000101: data <= 32'hc000bcaa;
    11'b00100000110: data <= 32'hb42a1ca7;
    11'b00100000111: data <= 32'h38073b3a;
    11'b00100001000: data <= 32'h35683588;
    11'b00100001001: data <= 32'h35e6b592;
    11'b00100001010: data <= 32'h38c838e1;
    11'b00100001011: data <= 32'h31f140e1;
    11'b00100001100: data <= 32'hb8c34146;
    11'b00100001101: data <= 32'hb7bb38e7;
    11'b00100001110: data <= 32'h38cabda1;
    11'b00100001111: data <= 32'h3cb1be10;
    11'b00100010000: data <= 32'h38b3b7f8;
    11'b00100010001: data <= 32'h32edafa6;
    11'b00100010010: data <= 32'h3cbcb735;
    11'b00100010011: data <= 32'h405bb5d0;
    11'b00100010100: data <= 32'h3cab3188;
    11'b00100010101: data <= 32'hbd5c2cbb;
    11'b00100010110: data <= 32'hc14fba31;
    11'b00100010111: data <= 32'hbe4fbca6;
    11'b00100011000: data <= 32'h2d2bb914;
    11'b00100011001: data <= 32'h34b1b4f4;
    11'b00100011010: data <= 32'hb7adba8e;
    11'b00100011011: data <= 32'hb8a5bb0c;
    11'b00100011100: data <= 32'h2c4239b9;
    11'b00100011101: data <= 32'h30ce4165;
    11'b00100011110: data <= 32'hb8c74158;
    11'b00100011111: data <= 32'hbbc738b7;
    11'b00100100000: data <= 32'hb674bc15;
    11'b00100100001: data <= 32'h3247b871;
    11'b00100100010: data <= 32'h33dd38fa;
    11'b00100100011: data <= 32'h38ef3871;
    11'b00100100100: data <= 32'h3f7fb66e;
    11'b00100100101: data <= 32'h4152b833;
    11'b00100100110: data <= 32'h3db435da;
    11'b00100100111: data <= 32'hbb2139f2;
    11'b00100101000: data <= 32'hbef5add4;
    11'b00100101001: data <= 32'hb7bdbc47;
    11'b00100101010: data <= 32'h39eabd35;
    11'b00100101011: data <= 32'h3312bd4f;
    11'b00100101100: data <= 32'hbb7abe81;
    11'b00100101101: data <= 32'hba53bd3e;
    11'b00100101110: data <= 32'h35943562;
    11'b00100101111: data <= 32'h38554009;
    11'b00100110000: data <= 32'hb9ad3f43;
    11'b00100110001: data <= 32'hbf3f2e82;
    11'b00100110010: data <= 32'hbe61ba09;
    11'b00100110011: data <= 32'hb9fc3322;
    11'b00100110100: data <= 32'hb2073d06;
    11'b00100110101: data <= 32'h3715392f;
    11'b00100110110: data <= 32'h3e43b8a7;
    11'b00100110111: data <= 32'h4061b593;
    11'b00100111000: data <= 32'h3ce13cdb;
    11'b00100111001: data <= 32'hb6b43fbf;
    11'b00100111010: data <= 32'hb9b13a7f;
    11'b00100111011: data <= 32'h37a7ba5c;
    11'b00100111100: data <= 32'h3c79bdc9;
    11'b00100111101: data <= 32'h3058bdd1;
    11'b00100111110: data <= 32'hbaf2be56;
    11'b00100111111: data <= 32'hb05fbda1;
    11'b00101000000: data <= 32'h3d7bb4b5;
    11'b00101000001: data <= 32'h3d1d3b09;
    11'b00101000010: data <= 32'hb97939b0;
    11'b00101000011: data <= 32'hc0a8b670;
    11'b00101000100: data <= 32'hc04eb916;
    11'b00101000101: data <= 32'hbc4d368d;
    11'b00101000110: data <= 32'hb7f53bbc;
    11'b00101000111: data <= 32'hb365ab46;
    11'b00101001000: data <= 32'h37b6bc5d;
    11'b00101001001: data <= 32'h3c98b07a;
    11'b00101001010: data <= 32'h3a42401a;
    11'b00101001011: data <= 32'hb08741b3;
    11'b00101001100: data <= 32'hb24b3d92;
    11'b00101001101: data <= 32'h3908b6ed;
    11'b00101001110: data <= 32'h3a68bb3a;
    11'b00101001111: data <= 32'hb08ab8bc;
    11'b00101010000: data <= 32'hb831ba2b;
    11'b00101010001: data <= 32'h3aeabcbb;
    11'b00101010010: data <= 32'h40f9ba8d;
    11'b00101010011: data <= 32'h3fe2271d;
    11'b00101010100: data <= 32'hb6d53109;
    11'b00101010101: data <= 32'hc02eb6e2;
    11'b00101010110: data <= 32'hbea7b834;
    11'b00101010111: data <= 32'hb8b82c34;
    11'b00101011000: data <= 32'hb84d206e;
    11'b00101011001: data <= 32'hbc08bcad;
    11'b00101011010: data <= 32'hb934befc;
    11'b00101011011: data <= 32'h34f1b1f6;
    11'b00101011100: data <= 32'h38644071;
    11'b00101011101: data <= 32'hac3841a8;
    11'b00101011110: data <= 32'hb6503d13;
    11'b00101011111: data <= 32'hae6db1a0;
    11'b00101100000: data <= 32'haf3d25e3;
    11'b00101100001: data <= 32'hb9053988;
    11'b00101100010: data <= 32'hb51d326c;
    11'b00101100011: data <= 32'h3dc1bb5c;
    11'b00101100100: data <= 32'h41dabc1d;
    11'b00101100101: data <= 32'h405bab98;
    11'b00101100110: data <= 32'habb1384c;
    11'b00101100111: data <= 32'hbcc7317a;
    11'b00101101000: data <= 32'hb6c5b47c;
    11'b00101101001: data <= 32'h358eb5ed;
    11'b00101101010: data <= 32'hb637baee;
    11'b00101101011: data <= 32'hbdf1bfcb;
    11'b00101101100: data <= 32'hbc81c05a;
    11'b00101101101: data <= 32'h3499b848;
    11'b00101101110: data <= 32'h3aa93e2c;
    11'b00101101111: data <= 32'ha7963f5f;
    11'b00101110000: data <= 32'hbbd33839;
    11'b00101110001: data <= 32'hbc7db015;
    11'b00101110010: data <= 32'hbc283a72;
    11'b00101110011: data <= 32'hbc723e4f;
    11'b00101110100: data <= 32'hb82538de;
    11'b00101110101: data <= 32'h3c71bbb6;
    11'b00101110110: data <= 32'h40b2bbe1;
    11'b00101110111: data <= 32'h3f033824;
    11'b00101111000: data <= 32'h32b43e25;
    11'b00101111001: data <= 32'hb1833c3c;
    11'b00101111010: data <= 32'h3a3a2d8f;
    11'b00101111011: data <= 32'h3c33b6fe;
    11'b00101111100: data <= 32'hb4f4bb9e;
    11'b00101111101: data <= 32'hbe20bf4c;
    11'b00101111110: data <= 32'hba00c032;
    11'b00101111111: data <= 32'h3c5dbbeb;
    11'b00110000000: data <= 32'h3e3136a3;
    11'b00110000001: data <= 32'h2f993817;
    11'b00110000010: data <= 32'hbd79b4e1;
    11'b00110000011: data <= 32'hbe78b24f;
    11'b00110000100: data <= 32'hbd3f3c54;
    11'b00110000101: data <= 32'hbd333e47;
    11'b00110000110: data <= 32'hbc3730a7;
    11'b00110000111: data <= 32'h2874bdbe;
    11'b00110001000: data <= 32'h3c64bb56;
    11'b00110001001: data <= 32'h3beb3cc2;
    11'b00110001010: data <= 32'h347840bb;
    11'b00110001011: data <= 32'h369b3e6d;
    11'b00110001100: data <= 32'h3cda362a;
    11'b00110001101: data <= 32'h3c0023cb;
    11'b00110001110: data <= 32'hb83aade0;
    11'b00110001111: data <= 32'hbd56ba97;
    11'b00110010000: data <= 32'h2b21be42;
    11'b00110010001: data <= 32'h4034bd31;
    11'b00110010010: data <= 32'h4074b7d4;
    11'b00110010011: data <= 32'h35d9b53f;
    11'b00110010100: data <= 32'hbcb0b905;
    11'b00110010101: data <= 32'hbc7bb194;
    11'b00110010110: data <= 32'hb9543b13;
    11'b00110010111: data <= 32'hbc3e3aa6;
    11'b00110011000: data <= 32'hbe79babb;
    11'b00110011001: data <= 32'hbc8ac02e;
    11'b00110011010: data <= 32'ha6a4bc00;
    11'b00110011011: data <= 32'h36fd3d6b;
    11'b00110011100: data <= 32'h338840a7;
    11'b00110011101: data <= 32'h35a23d6b;
    11'b00110011110: data <= 32'h39cf3677;
    11'b00110011111: data <= 32'h339439f8;
    11'b00110100000: data <= 32'hbc143ce2;
    11'b00110100001: data <= 32'hbcd236ce;
    11'b00110100010: data <= 32'h38a8bbb5;
    11'b00110100011: data <= 32'h4107bd6c;
    11'b00110100100: data <= 32'h40adb999;
    11'b00110100101: data <= 32'h3857b2bc;
    11'b00110100110: data <= 32'hb719b2a7;
    11'b00110100111: data <= 32'h30a92c81;
    11'b00110101000: data <= 32'h384a386f;
    11'b00110101001: data <= 32'hb88a2970;
    11'b00110101010: data <= 32'hbfacbe56;
    11'b00110101011: data <= 32'hbee1c0eb;
    11'b00110101100: data <= 32'hb53bbcd8;
    11'b00110101101: data <= 32'h38053a7d;
    11'b00110101110: data <= 32'h340c3d43;
    11'b00110101111: data <= 32'haebe35dc;
    11'b00110110000: data <= 32'hb1942f42;
    11'b00110110001: data <= 32'hb9253d59;
    11'b00110110010: data <= 32'hbde74067;
    11'b00110110011: data <= 32'hbd483c81;
    11'b00110110100: data <= 32'h35a7ba05;
    11'b00110110101: data <= 32'h3fa9bd10;
    11'b00110110110: data <= 32'h3ec4b420;
    11'b00110110111: data <= 32'h37da390f;
    11'b00110111000: data <= 32'h362438ec;
    11'b00110111001: data <= 32'h3dbd36f5;
    11'b00110111010: data <= 32'h3e2d374f;
    11'b00110111011: data <= 32'hb265aec5;
    11'b00110111100: data <= 32'hbf8dbdc6;
    11'b00110111101: data <= 32'hbdebc063;
    11'b00110111110: data <= 32'h34a3bd7f;
    11'b00110111111: data <= 32'h3c83b018;
    11'b00111000000: data <= 32'h3697ae3c;
    11'b00111000001: data <= 32'hb7b1ba3b;
    11'b00111000010: data <= 32'hb98eb460;
    11'b00111000011: data <= 32'hbb3b3e0a;
    11'b00111000100: data <= 32'hbe1240a8;
    11'b00111000101: data <= 32'hbe6a3b09;
    11'b00111000110: data <= 32'hb85cbc6a;
    11'b00111000111: data <= 32'h38b9bcd6;
    11'b00111001000: data <= 32'h38ed35cf;
    11'b00111001001: data <= 32'h33203dcd;
    11'b00111001010: data <= 32'h3ab73c9e;
    11'b00111001011: data <= 32'h40023909;
    11'b00111001100: data <= 32'h3ef539a5;
    11'b00111001101: data <= 32'hb42f38c5;
    11'b00111001110: data <= 32'hbec5b617;
    11'b00111001111: data <= 32'hba02bd70;
    11'b00111010000: data <= 32'h3d06bd56;
    11'b00111010001: data <= 32'h3f2ebb10;
    11'b00111010010: data <= 32'h38c1bc48;
    11'b00111010011: data <= 32'hb6fabd83;
    11'b00111010100: data <= 32'hb54cb72c;
    11'b00111010101: data <= 32'hb2ab3d30;
    11'b00111010110: data <= 32'hbc003ec1;
    11'b00111010111: data <= 32'hbf4da7a3;
    11'b00111011000: data <= 32'hbe37bef4;
    11'b00111011001: data <= 32'hb953bd0a;
    11'b00111011010: data <= 32'hb3c2390e;
    11'b00111011011: data <= 32'habe43e13;
    11'b00111011100: data <= 32'h39f13aee;
    11'b00111011101: data <= 32'h3e85367a;
    11'b00111011110: data <= 32'h3c5b3c73;
    11'b00111011111: data <= 32'hb9bc3ef9;
    11'b00111100000: data <= 32'hbe373bf9;
    11'b00111100001: data <= 32'hb140b6ea;
    11'b00111100010: data <= 32'h3f01bc72;
    11'b00111100011: data <= 32'h3f8abc22;
    11'b00111100100: data <= 32'h388abc54;
    11'b00111100101: data <= 32'h8fd3bc71;
    11'b00111100110: data <= 32'h3a31b43b;
    11'b00111100111: data <= 32'h3c763bc3;
    11'b00111101000: data <= 32'hb1783b03;
    11'b00111101001: data <= 32'hbf42baa6;
    11'b00111101010: data <= 32'hc01bc033;
    11'b00111101011: data <= 32'hbc6ebd3d;
    11'b00111101100: data <= 32'hb5f7357f;
    11'b00111101101: data <= 32'hb0833949;
    11'b00111101110: data <= 32'h34acb377;
    11'b00111101111: data <= 32'h39eeb306;
    11'b00111110000: data <= 32'h31ac3d80;
    11'b00111110001: data <= 32'hbcb5413e;
    11'b00111110010: data <= 32'hbe333f65;
    11'b00111110011: data <= 32'hb1a324a3;
    11'b00111110100: data <= 32'h3d2ebb0e;
    11'b00111110101: data <= 32'h3c92b8bb;
    11'b00111110110: data <= 32'h323fb481;
    11'b00111110111: data <= 32'h37e5b499;
    11'b00111111000: data <= 32'h3fcb2ef3;
    11'b00111111001: data <= 32'h40903a58;
    11'b00111111010: data <= 32'h3797386a;
    11'b00111111011: data <= 32'hbe65ba99;
    11'b00111111100: data <= 32'hbf33bf0a;
    11'b00111111101: data <= 32'hb87cbcb4;
    11'b00111111110: data <= 32'h32deb447;
    11'b00111111111: data <= 32'h24cbb90d;
    11'b01000000000: data <= 32'hb034be2e;
    11'b01000000001: data <= 32'h2d6cbb55;
    11'b01000000010: data <= 32'hb2a53d49;
    11'b01000000011: data <= 32'hbcae4170;
    11'b01000000100: data <= 32'hbe493eca;
    11'b01000000101: data <= 32'hba17b406;
    11'b01000000110: data <= 32'h2e0fba71;
    11'b01000000111: data <= 32'hae812b45;
    11'b01000001000: data <= 32'hb6843913;
    11'b01000001001: data <= 32'h398235cb;
    11'b01000001010: data <= 32'h40f2347e;
    11'b01000001011: data <= 32'h41323a92;
    11'b01000001100: data <= 32'h38543bb4;
    11'b01000001101: data <= 32'hbd6a2f02;
    11'b01000001110: data <= 32'hbc37ba1d;
    11'b01000001111: data <= 32'h3781ba4f;
    11'b01000010000: data <= 32'h3bc8b9e2;
    11'b01000010001: data <= 32'h325dbe34;
    11'b01000010010: data <= 32'hb436c094;
    11'b01000010011: data <= 32'h31eebd13;
    11'b01000010100: data <= 32'h35ac3c17;
    11'b01000010101: data <= 32'hb8154021;
    11'b01000010110: data <= 32'hbdc93a0e;
    11'b01000010111: data <= 32'hbddcbba0;
    11'b01000011000: data <= 32'hbc65baeb;
    11'b01000011001: data <= 32'hbc86376a;
    11'b01000011010: data <= 32'hbb5b3b7a;
    11'b01000011011: data <= 32'h377832b6;
    11'b01000011100: data <= 32'h402cabf3;
    11'b01000011101: data <= 32'h3fce3b31;
    11'b01000011110: data <= 32'h2a723f32;
    11'b01000011111: data <= 32'hbce73da9;
    11'b01000100000: data <= 32'hb5c935a4;
    11'b01000100001: data <= 32'h3caab4ac;
    11'b01000100010: data <= 32'h3cccb9c3;
    11'b01000100011: data <= 32'h2d51be31;
    11'b01000100100: data <= 32'hb02ac020;
    11'b01000100101: data <= 32'h3bdcbc5c;
    11'b01000100110: data <= 32'h3e643998;
    11'b01000100111: data <= 32'h38233cb0;
    11'b01000101000: data <= 32'hbc80b2fc;
    11'b01000101001: data <= 32'hbf0cbdce;
    11'b01000101010: data <= 32'hbe19bad6;
    11'b01000101011: data <= 32'hbd5e371e;
    11'b01000101100: data <= 32'hbc3635fb;
    11'b01000101101: data <= 32'h1032ba67;
    11'b01000101110: data <= 32'h3c8dbb0f;
    11'b01000101111: data <= 32'h3b283aa1;
    11'b01000110000: data <= 32'hb85740e2;
    11'b01000110001: data <= 32'hbcc2407f;
    11'b01000110010: data <= 32'hb0693b62;
    11'b01000110011: data <= 32'h3bf22a25;
    11'b01000110100: data <= 32'h3874b37f;
    11'b01000110101: data <= 32'hb796b9a1;
    11'b01000110110: data <= 32'h259bbc85;
    11'b01000110111: data <= 32'h3f9bb8c6;
    11'b01000111000: data <= 32'h417c3817;
    11'b01000111001: data <= 32'h3d453929;
    11'b01000111010: data <= 32'hb9f2b7b7;
    11'b01000111011: data <= 32'hbdb8bce6;
    11'b01000111100: data <= 32'hbb91b872;
    11'b01000111101: data <= 32'hb9783187;
    11'b01000111110: data <= 32'hba62b934;
    11'b01000111111: data <= 32'hb6b9c02c;
    11'b01001000000: data <= 32'h34fcbf0e;
    11'b01001000001: data <= 32'h34113876;
    11'b01001000010: data <= 32'hb95240da;
    11'b01001000011: data <= 32'hbc4b4025;
    11'b01001000100: data <= 32'hb6543903;
    11'b01001000101: data <= 32'h2c692c36;
    11'b01001000110: data <= 32'hb944368f;
    11'b01001000111: data <= 32'hbd2135a8;
    11'b01001001000: data <= 32'ha96ab3cd;
    11'b01001001001: data <= 32'h4090b47f;
    11'b01001001010: data <= 32'h421736f7;
    11'b01001001011: data <= 32'h3d9d39fd;
    11'b01001001100: data <= 32'hb8163175;
    11'b01001001101: data <= 32'hb96bb44a;
    11'b01001001110: data <= 32'h32712a40;
    11'b01001001111: data <= 32'h34969904;
    11'b01001010000: data <= 32'hb779bd99;
    11'b01001010001: data <= 32'hb8fec1a9;
    11'b01001010010: data <= 32'h3025c05e;
    11'b01001010011: data <= 32'h3841330d;
    11'b01001010100: data <= 32'habf63efc;
    11'b01001010101: data <= 32'hb9dd3c24;
    11'b01001010110: data <= 32'hba45b421;
    11'b01001010111: data <= 32'hbb73b07e;
    11'b01001011000: data <= 32'hbec83ae7;
    11'b01001011001: data <= 32'hbfa43b46;
    11'b01001011010: data <= 32'hb5b4af20;
    11'b01001011011: data <= 32'h3f65b85a;
    11'b01001011100: data <= 32'h40a43501;
    11'b01001011101: data <= 32'h3a1f3d08;
    11'b01001011110: data <= 32'hb81e3d0d;
    11'b01001011111: data <= 32'h29cf3ae8;
    11'b01001100000: data <= 32'h3c8439a2;
    11'b01001100001: data <= 32'h3a5d3115;
    11'b01001100010: data <= 32'hb7abbd4f;
    11'b01001100011: data <= 32'hb956c119;
    11'b01001100100: data <= 32'h38cdbf99;
    11'b01001100101: data <= 32'h3e2e1b1d;
    11'b01001100110: data <= 32'h3bd43aa8;
    11'b01001100111: data <= 32'hb2fbb0bc;
    11'b01001101000: data <= 32'hbb14bc21;
    11'b01001101001: data <= 32'hbd0fb413;
    11'b01001101010: data <= 32'hbf823bf0;
    11'b01001101011: data <= 32'hbff53956;
    11'b01001101100: data <= 32'hba03bb04;
    11'b01001101101: data <= 32'h3b07bd79;
    11'b01001101110: data <= 32'h3c4e274d;
    11'b01001101111: data <= 32'hae053ea9;
    11'b01001110000: data <= 32'hb8f53fed;
    11'b01001110001: data <= 32'h363e3db6;
    11'b01001110010: data <= 32'h3d0e3c30;
    11'b01001110011: data <= 32'h368f38f3;
    11'b01001110100: data <= 32'hbc19b750;
    11'b01001110101: data <= 32'hb9e2bdd0;
    11'b01001110110: data <= 32'h3d03bca1;
    11'b01001110111: data <= 32'h411ca847;
    11'b01001111000: data <= 32'h3f2d32aa;
    11'b01001111001: data <= 32'h3322b9ab;
    11'b01001111010: data <= 32'hb836bc4f;
    11'b01001111011: data <= 32'hb934212b;
    11'b01001111100: data <= 32'hbc573b7f;
    11'b01001111101: data <= 32'hbe10ac96;
    11'b01001111110: data <= 32'hbc17c006;
    11'b01001111111: data <= 32'ha60fc08f;
    11'b01010000000: data <= 32'h30dab5a2;
    11'b01010000001: data <= 32'hb8053e48;
    11'b01010000010: data <= 32'hb8843f08;
    11'b01010000011: data <= 32'h35653c1e;
    11'b01010000100: data <= 32'h391b3b1b;
    11'b01010000101: data <= 32'hb9163c83;
    11'b01010000110: data <= 32'hbf7d3949;
    11'b01010000111: data <= 32'hbb9cb4c1;
    11'b01010001000: data <= 32'h3e0ab85d;
    11'b01010001001: data <= 32'h4197a4e4;
    11'b01010001010: data <= 32'h3f3f2ffc;
    11'b01010001011: data <= 32'h3546b5d1;
    11'b01010001100: data <= 32'h2f98b4f5;
    11'b01010001101: data <= 32'h3864393d;
    11'b01010001110: data <= 32'h30563b8f;
    11'b01010001111: data <= 32'hbb17b942;
    11'b01010010000: data <= 32'hbc70c15e;
    11'b01010010001: data <= 32'hb5eec154;
    11'b01010010010: data <= 32'h2f62b8f3;
    11'b01010010011: data <= 32'haf3d3bb1;
    11'b01010010100: data <= 32'hb23a395e;
    11'b01010010101: data <= 32'h30e8ad43;
    11'b01010010110: data <= 32'hb1463648;
    11'b01010010111: data <= 32'hbe5f3dca;
    11'b01010011000: data <= 32'hc0ff3d70;
    11'b01010011001: data <= 32'hbd0130da;
    11'b01010011010: data <= 32'h3c6db88a;
    11'b01010011011: data <= 32'h400bb0cf;
    11'b01010011100: data <= 32'h3bc836b7;
    11'b01010011101: data <= 32'h2b493804;
    11'b01010011110: data <= 32'h399d39d5;
    11'b01010011111: data <= 32'h3e683d5a;
    11'b01010100000: data <= 32'h3bae3c97;
    11'b01010100001: data <= 32'hb90eb898;
    11'b01010100010: data <= 32'hbc88c0b5;
    11'b01010100011: data <= 32'haf39c06d;
    11'b01010100100: data <= 32'h3b03b8ca;
    11'b01010100101: data <= 32'h3a8b31cb;
    11'b01010100110: data <= 32'h35e6b901;
    11'b01010100111: data <= 32'h30a5bcad;
    11'b01010101000: data <= 32'hb72aa0be;
    11'b01010101001: data <= 32'hbeea3e1b;
    11'b01010101010: data <= 32'hc0e73d49;
    11'b01010101011: data <= 32'hbdceb578;
    11'b01010101100: data <= 32'h3419bd09;
    11'b01010101101: data <= 32'h3966b7db;
    11'b01010101110: data <= 32'hb224398a;
    11'b01010101111: data <= 32'hb5993c86;
    11'b01010110000: data <= 32'h3bc43d01;
    11'b01010110001: data <= 32'h3fb83e66;
    11'b01010110010: data <= 32'h3aea3ddb;
    11'b01010110011: data <= 32'hbc103252;
    11'b01010110100: data <= 32'hbd03bca8;
    11'b01010110101: data <= 32'h3605bcb9;
    11'b01010110110: data <= 32'h3f0cb53f;
    11'b01010110111: data <= 32'h3e5cb58d;
    11'b01010111000: data <= 32'h3a2fbd7b;
    11'b01010111001: data <= 32'h36aabe15;
    11'b01010111010: data <= 32'h2e2c2c19;
    11'b01010111011: data <= 32'hbad93e0a;
    11'b01010111100: data <= 32'hbed83a1e;
    11'b01010111101: data <= 32'hbdafbd48;
    11'b01010111110: data <= 32'hb84bc03e;
    11'b01010111111: data <= 32'hb6d0bafb;
    11'b01011000000: data <= 32'hbb653908;
    11'b01011000001: data <= 32'hb8283b91;
    11'b01011000010: data <= 32'h3b7e3a47;
    11'b01011000011: data <= 32'h3dfd3cd7;
    11'b01011000100: data <= 32'h1a163ec6;
    11'b01011000101: data <= 32'hbf373ccd;
    11'b01011000110: data <= 32'hbdfe310d;
    11'b01011000111: data <= 32'h38e6b363;
    11'b01011001000: data <= 32'h4004ab2b;
    11'b01011001001: data <= 32'h3e35b6cd;
    11'b01011001010: data <= 32'h398abce7;
    11'b01011001011: data <= 32'h3a88bbbc;
    11'b01011001100: data <= 32'h3cbd390e;
    11'b01011001101: data <= 32'h38293e43;
    11'b01011001110: data <= 32'hb9e933c2;
    11'b01011001111: data <= 32'hbce4bfe0;
    11'b01011010000: data <= 32'hbad3c0ed;
    11'b01011010001: data <= 32'hb959bbfd;
    11'b01011010010: data <= 32'hba3f3310;
    11'b01011010011: data <= 32'hb406a979;
    11'b01011010100: data <= 32'h3a79b785;
    11'b01011010101: data <= 32'h3a593610;
    11'b01011010110: data <= 32'hbb3b3ed7;
    11'b01011010111: data <= 32'hc0cc3f62;
    11'b01011011000: data <= 32'hbed23a86;
    11'b01011011001: data <= 32'h35ce26a7;
    11'b01011011010: data <= 32'h3d43aa70;
    11'b01011011011: data <= 32'h38adb1e9;
    11'b01011011100: data <= 32'h2e81b7d8;
    11'b01011011101: data <= 32'h3c619e61;
    11'b01011011110: data <= 32'h40563d2c;
    11'b01011011111: data <= 32'h3e373ee1;
    11'b01011100000: data <= 32'hb19c3306;
    11'b01011100001: data <= 32'hbc47bed0;
    11'b01011100010: data <= 32'hb91abf9c;
    11'b01011100011: data <= 32'habf7b981;
    11'b01011100100: data <= 32'h290eb43e;
    11'b01011100101: data <= 32'h34a3bd0d;
    11'b01011100110: data <= 32'h3a56bf0f;
    11'b01011100111: data <= 32'h373bb5b6;
    11'b01011101000: data <= 32'hbc5a3e4d;
    11'b01011101001: data <= 32'hc0883f54;
    11'b01011101010: data <= 32'hbe9b37f2;
    11'b01011101011: data <= 32'hb2d7b824;
    11'b01011101100: data <= 32'h2a10b5b7;
    11'b01011101101: data <= 32'hba482c57;
    11'b01011101110: data <= 32'hb94030e0;
    11'b01011101111: data <= 32'h3c783861;
    11'b01011110000: data <= 32'h41023dfb;
    11'b01011110001: data <= 32'h3e993f51;
    11'b01011110010: data <= 32'hb5f939fa;
    11'b01011110011: data <= 32'hbc88b8ba;
    11'b01011110100: data <= 32'hb1f6b95f;
    11'b01011110101: data <= 32'h3a5fab7c;
    11'b01011110110: data <= 32'h3a96b830;
    11'b01011110111: data <= 32'h3945bfff;
    11'b01011111000: data <= 32'h3b41c0a6;
    11'b01011111001: data <= 32'h3a4db814;
    11'b01011111010: data <= 32'hb4a73de1;
    11'b01011111011: data <= 32'hbd5f3d46;
    11'b01011111100: data <= 32'hbd10b6bc;
    11'b01011111101: data <= 32'hb9c8bd79;
    11'b01011111110: data <= 32'hbc23b9c4;
    11'b01011111111: data <= 32'hbef82f23;
    11'b01100000000: data <= 32'hbc5f3057;
    11'b01100000001: data <= 32'h3baf30e7;
    11'b01100000010: data <= 32'h403a3b95;
    11'b01100000011: data <= 32'h3b093ee3;
    11'b01100000100: data <= 32'hbc7c3dd9;
    11'b01100000101: data <= 32'hbd7839a0;
    11'b01100000110: data <= 32'h2f663822;
    11'b01100000111: data <= 32'h3caf3828;
    11'b01100001000: data <= 32'h3ad1b714;
    11'b01100001001: data <= 32'h3733bf94;
    11'b01100001010: data <= 32'h3c02bf92;
    11'b01100001011: data <= 32'h3e62a3fd;
    11'b01100001100: data <= 32'h3c333e0e;
    11'b01100001101: data <= 32'hb00d3a1d;
    11'b01100001110: data <= 32'hb9d5bca3;
    11'b01100001111: data <= 32'hbac1bf16;
    11'b01100010000: data <= 32'hbd3fba01;
    11'b01100010001: data <= 32'hbf03a837;
    11'b01100010010: data <= 32'hbb83b8bb;
    11'b01100010011: data <= 32'h3a79bc3d;
    11'b01100010100: data <= 32'h3d9cb005;
    11'b01100010101: data <= 32'had4b3d84;
    11'b01100010110: data <= 32'hbf143f88;
    11'b01100010111: data <= 32'hbe083d8e;
    11'b01100011000: data <= 32'h2d783bb0;
    11'b01100011001: data <= 32'h39b9397e;
    11'b01100011010: data <= 32'hac5eb0fd;
    11'b01100011011: data <= 32'hb5ecbcae;
    11'b01100011100: data <= 32'h3b52bb49;
    11'b01100011101: data <= 32'h40ab3982;
    11'b01100011110: data <= 32'h40363e83;
    11'b01100011111: data <= 32'h393c3885;
    11'b01100100000: data <= 32'hb5d1bc6c;
    11'b01100100001: data <= 32'hb86bbd0d;
    11'b01100100010: data <= 32'hb9d6b367;
    11'b01100100011: data <= 32'hbb96b12f;
    11'b01100100100: data <= 32'hb5fdbe38;
    11'b01100100101: data <= 32'h3a2dc0be;
    11'b01100100110: data <= 32'h3b68bc6a;
    11'b01100100111: data <= 32'hb7413bdf;
    11'b01100101000: data <= 32'hbeca3f08;
    11'b01100101001: data <= 32'hbd183c69;
    11'b01100101010: data <= 32'hb0e83793;
    11'b01100101011: data <= 32'hb4bd3631;
    11'b01100101100: data <= 32'hbdce2ecf;
    11'b01100101101: data <= 32'hbd8db6e0;
    11'b01100101110: data <= 32'h391ab24d;
    11'b01100101111: data <= 32'h410c3bb0;
    11'b01100110000: data <= 32'h407a3e5d;
    11'b01100110001: data <= 32'h38703a42;
    11'b01100110010: data <= 32'hb611b3db;
    11'b01100110011: data <= 32'hada1a611;
    11'b01100110100: data <= 32'h32393957;
    11'b01100110101: data <= 32'ha865adcb;
    11'b01100110110: data <= 32'h2c98c03e;
    11'b01100110111: data <= 32'h3a38c1f3;
    11'b01100111000: data <= 32'h3be1bd96;
    11'b01100111001: data <= 32'h2e563a45;
    11'b01100111010: data <= 32'hba373cde;
    11'b01100111011: data <= 32'hb8f730a7;
    11'b01100111100: data <= 32'hb504b798;
    11'b01100111101: data <= 32'hbcbfaaae;
    11'b01100111110: data <= 32'hc0eb3333;
    11'b01100111111: data <= 32'hc003b2ab;
    11'b01101000000: data <= 32'h355eb5b2;
    11'b01101000001: data <= 32'h402c36ea;
    11'b01101000010: data <= 32'h3dcc3ceb;
    11'b01101000011: data <= 32'hb4143c91;
    11'b01101000100: data <= 32'hb96b3abc;
    11'b01101000101: data <= 32'h34363ce3;
    11'b01101000110: data <= 32'h3a283dde;
    11'b01101000111: data <= 32'h32f331f2;
    11'b01101001000: data <= 32'hae4cbfc6;
    11'b01101001001: data <= 32'h392ac115;
    11'b01101001010: data <= 32'h3dc6bb0b;
    11'b01101001011: data <= 32'h3ce33af3;
    11'b01101001100: data <= 32'h37fa3905;
    11'b01101001101: data <= 32'h3179ba14;
    11'b01101001110: data <= 32'hb22cbc56;
    11'b01101001111: data <= 32'hbd79b075;
    11'b01101010000: data <= 32'hc0fb3463;
    11'b01101010001: data <= 32'hbf81b8d0;
    11'b01101010010: data <= 32'h3235bd60;
    11'b01101010011: data <= 32'h3d62b98f;
    11'b01101010100: data <= 32'h359938e2;
    11'b01101010101: data <= 32'hbc5f3d1e;
    11'b01101010110: data <= 32'hbb1f3da4;
    11'b01101010111: data <= 32'h36443ed4;
    11'b01101011000: data <= 32'h38ff3ed7;
    11'b01101011001: data <= 32'hb79a3805;
    11'b01101011010: data <= 32'hbbaebcc2;
    11'b01101011011: data <= 32'h3466bdcd;
    11'b01101011100: data <= 32'h3f7aa07e;
    11'b01101011101: data <= 32'h40473c43;
    11'b01101011110: data <= 32'h3d5d34d5;
    11'b01101011111: data <= 32'h3955bbee;
    11'b01101100000: data <= 32'h31aeba72;
    11'b01101100001: data <= 32'hb9ff3675;
    11'b01101100010: data <= 32'hbe6b36c3;
    11'b01101100011: data <= 32'hbcb0bcf3;
    11'b01101100100: data <= 32'h33b6c101;
    11'b01101100101: data <= 32'h3a2abeff;
    11'b01101100110: data <= 32'hb4822883;
    11'b01101100111: data <= 32'hbd023c18;
    11'b01101101000: data <= 32'hb93c3c4d;
    11'b01101101001: data <= 32'h36a03cae;
    11'b01101101010: data <= 32'haafc3d3e;
    11'b01101101011: data <= 32'hbec53986;
    11'b01101101100: data <= 32'hc020b5fa;
    11'b01101101101: data <= 32'hb32db801;
    11'b01101101110: data <= 32'h3f8637f6;
    11'b01101101111: data <= 32'h406b3c35;
    11'b01101110000: data <= 32'h3ce43480;
    11'b01101110001: data <= 32'h38cdb765;
    11'b01101110010: data <= 32'h38ba341b;
    11'b01101110011: data <= 32'h33863d92;
    11'b01101110100: data <= 32'hb7b039fb;
    11'b01101110101: data <= 32'hb7edbe56;
    11'b01101110110: data <= 32'h34bdc20e;
    11'b01101110111: data <= 32'h38f7c01c;
    11'b01101111000: data <= 32'haafeb16a;
    11'b01101111001: data <= 32'hb82b37fd;
    11'b01101111010: data <= 32'h2d5e2c1d;
    11'b01101111011: data <= 32'h38392943;
    11'b01101111100: data <= 32'hb98c3936;
    11'b01101111101: data <= 32'hc13939e9;
    11'b01101111110: data <= 32'hc17426e4;
    11'b01101111111: data <= 32'hb8b3b57e;
    11'b01110000000: data <= 32'h3dab3192;
    11'b01110000001: data <= 32'h3d7838f7;
    11'b01110000010: data <= 32'h343835b9;
    11'b01110000011: data <= 32'h2ebb3596;
    11'b01110000100: data <= 32'h3ae43d9e;
    11'b01110000101: data <= 32'h3bb04088;
    11'b01110000110: data <= 32'h2cc23c8f;
    11'b01110000111: data <= 32'hb717bd5b;
    11'b01110001000: data <= 32'h2fa4c115;
    11'b01110001001: data <= 32'h3a65bdb1;
    11'b01110001010: data <= 32'h3a302d20;
    11'b01110001011: data <= 32'h392ba19c;
    11'b01110001100: data <= 32'h3bcabbc0;
    11'b01110001101: data <= 32'h3a87bada;
    11'b01110001110: data <= 32'hba203542;
    11'b01110001111: data <= 32'hc12d3a6c;
    11'b01110010000: data <= 32'hc109ae81;
    11'b01110010001: data <= 32'hb8d9bc19;
    11'b01110010010: data <= 32'h39f0baa3;
    11'b01110010011: data <= 32'h30f9af12;
    11'b01110010100: data <= 32'hbac3348c;
    11'b01110010101: data <= 32'hb5a13a26;
    11'b01110010110: data <= 32'h3bcf3f5a;
    11'b01110010111: data <= 32'h3c3d40f2;
    11'b01110011000: data <= 32'hb4dd3d89;
    11'b01110011001: data <= 32'hbca5b906;
    11'b01110011010: data <= 32'hb5d1bd65;
    11'b01110011011: data <= 32'h3bdcb4cf;
    11'b01110011100: data <= 32'h3e07382c;
    11'b01110011101: data <= 32'h3dbfb4cb;
    11'b01110011110: data <= 32'h3deabdb1;
    11'b01110011111: data <= 32'h3cafbb2a;
    11'b01110100000: data <= 32'hb13439a7;
    11'b01110100001: data <= 32'hbe763c36;
    11'b01110100010: data <= 32'hbe5cb7a1;
    11'b01110100011: data <= 32'hb529bfe0;
    11'b01110100100: data <= 32'h330dbf51;
    11'b01110100101: data <= 32'hb971b9e4;
    11'b01110100110: data <= 32'hbd4da3f6;
    11'b01110100111: data <= 32'hb4de36a6;
    11'b01110101000: data <= 32'h3c523ce7;
    11'b01110101001: data <= 32'h392f3f89;
    11'b01110101010: data <= 32'hbd233d6c;
    11'b01110101011: data <= 32'hc0683009;
    11'b01110101100: data <= 32'hbb93b2c8;
    11'b01110101101: data <= 32'h3b263839;
    11'b01110101110: data <= 32'h3e1839c3;
    11'b01110101111: data <= 32'h3d07b610;
    11'b01110110000: data <= 32'h3d11bca5;
    11'b01110110001: data <= 32'h3d9cadc1;
    11'b01110110010: data <= 32'h3a173e7e;
    11'b01110110011: data <= 32'hb5223df0;
    11'b01110110100: data <= 32'hb8beb966;
    11'b01110110101: data <= 32'ha829c0d0;
    11'b01110110110: data <= 32'h28e1c02b;
    11'b01110110111: data <= 32'hb9bbbac2;
    11'b01110111000: data <= 32'hbaf5b678;
    11'b01110111001: data <= 32'h3587b85c;
    11'b01110111010: data <= 32'h3d40ab34;
    11'b01110111011: data <= 32'h32373b57;
    11'b01110111100: data <= 32'hc02c3c9e;
    11'b01110111101: data <= 32'hc1a73842;
    11'b01110111110: data <= 32'hbd0e3271;
    11'b01110111111: data <= 32'h38193802;
    11'b01111000000: data <= 32'h39b3366f;
    11'b01111000001: data <= 32'h3127b6c2;
    11'b01111000010: data <= 32'h37c5b882;
    11'b01111000011: data <= 32'h3dae3b55;
    11'b01111000100: data <= 32'h3de240ef;
    11'b01111000101: data <= 32'h37b03f83;
    11'b01111000110: data <= 32'hb32eb758;
    11'b01111000111: data <= 32'hac37bfb7;
    11'b01111001000: data <= 32'h2ed3bd56;
    11'b01111001001: data <= 32'hafe1b572;
    11'b01111001010: data <= 32'h302eb964;
    11'b01111001011: data <= 32'h3cd8be33;
    11'b01111001100: data <= 32'h3e95bcc2;
    11'b01111001101: data <= 32'h309e3432;
    11'b01111001110: data <= 32'hc01a3c2a;
    11'b01111001111: data <= 32'hc10b37ef;
    11'b01111010000: data <= 32'hbc44b35f;
    11'b01111010001: data <= 32'h2b0db4ec;
    11'b01111010010: data <= 32'hb77bb4d1;
    11'b01111010011: data <= 32'hbcb0b89c;
    11'b01111010100: data <= 32'hb4fdb2df;
    11'b01111010101: data <= 32'h3d503d45;
    11'b01111010110: data <= 32'h3e8e4134;
    11'b01111010111: data <= 32'h35c33fd1;
    11'b01111011000: data <= 32'hb9bf2c5a;
    11'b01111011001: data <= 32'hb80dba21;
    11'b01111011010: data <= 32'h31ea16d2;
    11'b01111011011: data <= 32'h37ef3715;
    11'b01111011100: data <= 32'h3af2b9e0;
    11'b01111011101: data <= 32'h3eadc01b;
    11'b01111011110: data <= 32'h3f8cbdf7;
    11'b01111011111: data <= 32'h38d6362b;
    11'b01111100000: data <= 32'hbc683ce6;
    11'b01111100001: data <= 32'hbd95338a;
    11'b01111100010: data <= 32'hb735bc18;
    11'b01111100011: data <= 32'hb345bced;
    11'b01111100100: data <= 32'hbd57bb39;
    11'b01111100101: data <= 32'hbfaeba89;
    11'b01111100110: data <= 32'hb864b788;
    11'b01111100111: data <= 32'h3d5939c6;
    11'b01111101000: data <= 32'h3d5e3f5b;
    11'b01111101001: data <= 32'hb70b3e74;
    11'b01111101010: data <= 32'hbea438a5;
    11'b01111101011: data <= 32'hbc513642;
    11'b01111101100: data <= 32'h2eb93c68;
    11'b01111101101: data <= 32'h387e3ba2;
    11'b01111101110: data <= 32'h3992b97b;
    11'b01111101111: data <= 32'h3d41bf97;
    11'b01111110000: data <= 32'h3f5bbb1d;
    11'b01111110001: data <= 32'h3d2f3cb2;
    11'b01111110010: data <= 32'h328e3e99;
    11'b01111110011: data <= 32'hb00a2c71;
    11'b01111110100: data <= 32'h31aebddc;
    11'b01111110101: data <= 32'hb3f8bdf2;
    11'b01111110110: data <= 32'hbddfbb36;
    11'b01111110111: data <= 32'hbec2bbc7;
    11'b01111111000: data <= 32'hab5bbce2;
    11'b01111111001: data <= 32'h3e3ab887;
    11'b01111111010: data <= 32'h3b9938d6;
    11'b01111111011: data <= 32'hbcd43c3a;
    11'b01111111100: data <= 32'hc08b3a62;
    11'b01111111101: data <= 32'hbd473b21;
    11'b01111111110: data <= 32'hae0d3d4a;
    11'b01111111111: data <= 32'hac793aa4;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    