
module memory_rom_17(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3a193d91;
    11'b00000000001: data <= 32'h371139cb;
    11'b00000000010: data <= 32'hb6bbbb1e;
    11'b00000000011: data <= 32'h947bbf80;
    11'b00000000100: data <= 32'h3df4bb1e;
    11'b00000000101: data <= 32'h40673aea;
    11'b00000000110: data <= 32'h3dd23c3e;
    11'b00000000111: data <= 32'h362ab6a1;
    11'b00000001000: data <= 32'hb18bbd62;
    11'b00000001001: data <= 32'hb9d6b8ab;
    11'b00000001010: data <= 32'hbe263485;
    11'b00000001011: data <= 32'hbe4eb771;
    11'b00000001100: data <= 32'hb45dbfae;
    11'b00000001101: data <= 32'h3bc4bfa3;
    11'b00000001110: data <= 32'h37efb2c9;
    11'b00000001111: data <= 32'hbc163d48;
    11'b00000010000: data <= 32'hbda73e3a;
    11'b00000010001: data <= 32'hb4a33cfe;
    11'b00000010010: data <= 32'h35f53ca7;
    11'b00000010011: data <= 32'hb8e43a53;
    11'b00000010100: data <= 32'hbe90b37a;
    11'b00000010101: data <= 32'hb99cbac2;
    11'b00000010110: data <= 32'h3e26ac48;
    11'b00000010111: data <= 32'h41453c6f;
    11'b00000011000: data <= 32'h3f233bc0;
    11'b00000011001: data <= 32'h382cb361;
    11'b00000011010: data <= 32'h2f42b898;
    11'b00000011011: data <= 32'h26a83680;
    11'b00000011100: data <= 32'hb7353a46;
    11'b00000011101: data <= 32'hb987ba59;
    11'b00000011110: data <= 32'h9dc5c181;
    11'b00000011111: data <= 32'h3a06c14e;
    11'b00000100000: data <= 32'h35cab903;
    11'b00000100001: data <= 32'hb9483b9e;
    11'b00000100010: data <= 32'hba243ae9;
    11'b00000100011: data <= 32'ha44c346e;
    11'b00000100100: data <= 32'hb1483655;
    11'b00000100101: data <= 32'hbee83958;
    11'b00000100110: data <= 32'hc15e331b;
    11'b00000100111: data <= 32'hbd15b588;
    11'b00000101000: data <= 32'h3d029136;
    11'b00000101001: data <= 32'h40653a89;
    11'b00000101010: data <= 32'h3c663b1d;
    11'b00000101011: data <= 32'h970f363b;
    11'b00000101100: data <= 32'h331d3907;
    11'b00000101101: data <= 32'h3a1c3e3e;
    11'b00000101110: data <= 32'h36563d76;
    11'b00000101111: data <= 32'hb459b9c5;
    11'b00000110000: data <= 32'ha977c16f;
    11'b00000110001: data <= 32'h3a0ec0c7;
    11'b00000110010: data <= 32'h3b53b6a2;
    11'b00000110011: data <= 32'h36d73903;
    11'b00000110100: data <= 32'h34aaade0;
    11'b00000110101: data <= 32'h36f6ba9a;
    11'b00000110110: data <= 32'hb5fcb3ef;
    11'b00000110111: data <= 32'hc04838e4;
    11'b00000111000: data <= 32'hc1c834d3;
    11'b00000111001: data <= 32'hbd7fb96c;
    11'b00000111010: data <= 32'h3a61ba8c;
    11'b00000111011: data <= 32'h3cbc1bd8;
    11'b00000111100: data <= 32'had873957;
    11'b00000111101: data <= 32'hb9ba3b1c;
    11'b00000111110: data <= 32'h333a3dbb;
    11'b00000111111: data <= 32'h3c584056;
    11'b00001000000: data <= 32'h36c53ed9;
    11'b00001000001: data <= 32'hb9d3b427;
    11'b00001000010: data <= 32'hb87bbf5e;
    11'b00001000011: data <= 32'h3a30bd58;
    11'b00001000100: data <= 32'h3e993296;
    11'b00001000101: data <= 32'h3df93759;
    11'b00001000110: data <= 32'h3c8db9e9;
    11'b00001000111: data <= 32'h3b06bd22;
    11'b00001001000: data <= 32'ha95fb1d0;
    11'b00001001001: data <= 32'hbe453b03;
    11'b00001001010: data <= 32'hc05130a8;
    11'b00001001011: data <= 32'hbbefbe0f;
    11'b00001001100: data <= 32'h36b7bff0;
    11'b00001001101: data <= 32'h3396bb28;
    11'b00001001110: data <= 32'hbb8234df;
    11'b00001001111: data <= 32'hbbf33a90;
    11'b00001010000: data <= 32'h355e3d0f;
    11'b00001010001: data <= 32'h3ba63f69;
    11'b00001010010: data <= 32'hb52d3e8f;
    11'b00001010011: data <= 32'hbf453515;
    11'b00001010100: data <= 32'hbd6fb99f;
    11'b00001010101: data <= 32'h38fcb39d;
    11'b00001010110: data <= 32'h3fc23996;
    11'b00001010111: data <= 32'h3f123621;
    11'b00001011000: data <= 32'h3ceaba60;
    11'b00001011001: data <= 32'h3c4eba9a;
    11'b00001011010: data <= 32'h393d394a;
    11'b00001011011: data <= 32'hb6343deb;
    11'b00001011100: data <= 32'hbc112a31;
    11'b00001011101: data <= 32'hb78ac055;
    11'b00001011110: data <= 32'h33cec156;
    11'b00001011111: data <= 32'hafa2bd39;
    11'b00001100000: data <= 32'hbb29a83c;
    11'b00001100001: data <= 32'hb81d30fe;
    11'b00001100010: data <= 32'h39a132c3;
    11'b00001100011: data <= 32'h395d3ada;
    11'b00001100100: data <= 32'hbcea3d14;
    11'b00001100101: data <= 32'hc19839af;
    11'b00001100110: data <= 32'hbfda9916;
    11'b00001100111: data <= 32'h34f530cf;
    11'b00001101000: data <= 32'h3dfa38c8;
    11'b00001101001: data <= 32'h3c09332f;
    11'b00001101010: data <= 32'h3816b709;
    11'b00001101011: data <= 32'h3bab3097;
    11'b00001101100: data <= 32'h3d473eff;
    11'b00001101101: data <= 32'h391d4042;
    11'b00001101110: data <= 32'hb4663288;
    11'b00001101111: data <= 32'hb4a8c02d;
    11'b00001110000: data <= 32'h322dc0ae;
    11'b00001110001: data <= 32'h316cbb81;
    11'b00001110010: data <= 32'hac09b147;
    11'b00001110011: data <= 32'h3783b9d2;
    11'b00001110100: data <= 32'h3d01bc36;
    11'b00001110101: data <= 32'h38c1aec1;
    11'b00001110110: data <= 32'hbe423bca;
    11'b00001110111: data <= 32'hc1e63a87;
    11'b00001111000: data <= 32'hbfd3acc8;
    11'b00001111001: data <= 32'h1e38b63f;
    11'b00001111010: data <= 32'h3852afe4;
    11'b00001111011: data <= 32'hb532aeef;
    11'b00001111100: data <= 32'hb816af5f;
    11'b00001111101: data <= 32'h39a93ab6;
    11'b00001111110: data <= 32'h3e8e40a0;
    11'b00001111111: data <= 32'h3b5540d4;
    11'b00010000000: data <= 32'hb6f53883;
    11'b00010000001: data <= 32'hb988bd04;
    11'b00010000010: data <= 32'h2e2ebc9b;
    11'b00010000011: data <= 32'h3991a71a;
    11'b00010000100: data <= 32'h3aeaacbc;
    11'b00010000101: data <= 32'h3d21bd68;
    11'b00010000110: data <= 32'h3ebabf01;
    11'b00010000111: data <= 32'h3b07b5a2;
    11'b00010001000: data <= 32'hbc0d3c5d;
    11'b00010001001: data <= 32'hc0323a1a;
    11'b00010001010: data <= 32'hbd3db976;
    11'b00010001011: data <= 32'hafbbbd8f;
    11'b00010001100: data <= 32'hb5eebbf0;
    11'b00010001101: data <= 32'hbda0b80b;
    11'b00010001110: data <= 32'hbc76b220;
    11'b00010001111: data <= 32'h391e395c;
    11'b00010010000: data <= 32'h3e603f9a;
    11'b00010010001: data <= 32'h3696403a;
    11'b00010010010: data <= 32'hbd523b47;
    11'b00010010011: data <= 32'hbdd2b109;
    11'b00010010100: data <= 32'haff23150;
    11'b00010010101: data <= 32'h3b683a6d;
    11'b00010010110: data <= 32'h3c742b33;
    11'b00010010111: data <= 32'h3d32bde5;
    11'b00010011000: data <= 32'h3ecebe2a;
    11'b00010011001: data <= 32'h3d7f3453;
    11'b00010011010: data <= 32'h2ff43e96;
    11'b00010011011: data <= 32'hb9fd3a12;
    11'b00010011100: data <= 32'hb721bceb;
    11'b00010011101: data <= 32'hac2dc00c;
    11'b00010011110: data <= 32'hba2abd68;
    11'b00010011111: data <= 32'hbe79b9bc;
    11'b00010100000: data <= 32'hbb14b993;
    11'b00010100001: data <= 32'h3b85b58b;
    11'b00010100010: data <= 32'h3da739b2;
    11'b00010100011: data <= 32'hb5a63da1;
    11'b00010100100: data <= 32'hc0793c37;
    11'b00010100101: data <= 32'hc00e3889;
    11'b00010100110: data <= 32'hb5d53a86;
    11'b00010100111: data <= 32'h38ba3bda;
    11'b00010101000: data <= 32'h361d9f79;
    11'b00010101001: data <= 32'h3695bce5;
    11'b00010101010: data <= 32'h3d0fb9f0;
    11'b00010101011: data <= 32'h3f243d0c;
    11'b00010101100: data <= 32'h3ca4408f;
    11'b00010101101: data <= 32'h34213b20;
    11'b00010101110: data <= 32'h29b5bcda;
    11'b00010101111: data <= 32'h223abed8;
    11'b00010110000: data <= 32'hb8adbab8;
    11'b00010110001: data <= 32'hbbdab881;
    11'b00010110010: data <= 32'ha5bebd58;
    11'b00010110011: data <= 32'h3de8be6f;
    11'b00010110100: data <= 32'h3d6cb81c;
    11'b00010110101: data <= 32'hb9a73a33;
    11'b00010110110: data <= 32'hc0c93bf6;
    11'b00010110111: data <= 32'hbf9e38b2;
    11'b00010111000: data <= 32'hb6cb37e7;
    11'b00010111001: data <= 32'hb07e369d;
    11'b00010111010: data <= 32'hbb90b53d;
    11'b00010111011: data <= 32'hbaf2bb9f;
    11'b00010111100: data <= 32'h394aac84;
    11'b00010111101: data <= 32'h3fa43f48;
    11'b00010111110: data <= 32'h3e0e40f6;
    11'b00010111111: data <= 32'h356a3c38;
    11'b00011000000: data <= 32'hb14ab894;
    11'b00011000001: data <= 32'hab50b83b;
    11'b00011000010: data <= 32'hb0573513;
    11'b00011000011: data <= 32'haf6daf5d;
    11'b00011000100: data <= 32'h3a2fbef9;
    11'b00011000101: data <= 32'h3f6cc0bd;
    11'b00011000110: data <= 32'h3dfbbc13;
    11'b00011000111: data <= 32'hb50a394c;
    11'b00011001000: data <= 32'hbe323b1e;
    11'b00011001001: data <= 32'hbc1e2c83;
    11'b00011001010: data <= 32'hb274b680;
    11'b00011001011: data <= 32'hba95b6bd;
    11'b00011001100: data <= 32'hc029b999;
    11'b00011001101: data <= 32'hbefdbb7d;
    11'b00011001110: data <= 32'h352caf61;
    11'b00011001111: data <= 32'h3f203dab;
    11'b00011010000: data <= 32'h3c6c3fe9;
    11'b00011010001: data <= 32'hb6c93c47;
    11'b00011010010: data <= 32'hbaf834b9;
    11'b00011010011: data <= 32'hb4543ab3;
    11'b00011010100: data <= 32'h306c3dbe;
    11'b00011010101: data <= 32'h3309351f;
    11'b00011010110: data <= 32'h3a70beff;
    11'b00011010111: data <= 32'h3ed4c083;
    11'b00011011000: data <= 32'h3ec5b87b;
    11'b00011011001: data <= 32'h38cd3c84;
    11'b00011011010: data <= 32'hb0ff3b11;
    11'b00011011011: data <= 32'h3027b7b4;
    11'b00011011100: data <= 32'h3204bc5c;
    11'b00011011101: data <= 32'hbc4fba61;
    11'b00011011110: data <= 32'hc0c6ba45;
    11'b00011011111: data <= 32'hbed9bcbd;
    11'b00011100000: data <= 32'h37f9bb63;
    11'b00011100001: data <= 32'h3e5d3236;
    11'b00011100010: data <= 32'h35db3bd0;
    11'b00011100011: data <= 32'hbd623ae1;
    11'b00011100100: data <= 32'hbdd53acd;
    11'b00011100101: data <= 32'hb6c13e55;
    11'b00011100110: data <= 32'h224e3f5f;
    11'b00011100111: data <= 32'hb52f36c6;
    11'b00011101000: data <= 32'haee8bde7;
    11'b00011101001: data <= 32'h3beebe04;
    11'b00011101010: data <= 32'h3ef8369a;
    11'b00011101011: data <= 32'h3dca3f13;
    11'b00011101100: data <= 32'h3b923bac;
    11'b00011101101: data <= 32'h3b0fb901;
    11'b00011101110: data <= 32'h37a4bb85;
    11'b00011101111: data <= 32'hbac6b45f;
    11'b00011110000: data <= 32'hbf44b604;
    11'b00011110001: data <= 32'hbb3abde3;
    11'b00011110010: data <= 32'h3c1ebff3;
    11'b00011110011: data <= 32'h3e02bc80;
    11'b00011110100: data <= 32'haebd2ac5;
    11'b00011110101: data <= 32'hbe8e3859;
    11'b00011110110: data <= 32'hbd573a64;
    11'b00011110111: data <= 32'hb42e3d5e;
    11'b00011111000: data <= 32'hb6393d78;
    11'b00011111001: data <= 32'hbdce3037;
    11'b00011111010: data <= 32'hbde8bcc1;
    11'b00011111011: data <= 32'h2d01ba07;
    11'b00011111100: data <= 32'h3e473c56;
    11'b00011111101: data <= 32'h3ed13fee;
    11'b00011111110: data <= 32'h3c7c3b85;
    11'b00011111111: data <= 32'h3a79b48b;
    11'b00100000000: data <= 32'h37862a0b;
    11'b00100000001: data <= 32'hb6383bba;
    11'b00100000010: data <= 32'hbb41363a;
    11'b00100000011: data <= 32'ha4d0be36;
    11'b00100000100: data <= 32'h3dbcc141;
    11'b00100000101: data <= 32'h3dfebef1;
    11'b00100000110: data <= 32'h25a5b3bf;
    11'b00100000111: data <= 32'hbbdb3552;
    11'b00100001000: data <= 32'hb636344f;
    11'b00100001001: data <= 32'h346536dd;
    11'b00100001010: data <= 32'hb9d83793;
    11'b00100001011: data <= 32'hc0e5b45d;
    11'b00100001100: data <= 32'hc0f1bc45;
    11'b00100001101: data <= 32'hb7c4b891;
    11'b00100001110: data <= 32'h3d263ae2;
    11'b00100001111: data <= 32'h3d133db3;
    11'b00100010000: data <= 32'h35fb3940;
    11'b00100010001: data <= 32'h2d1533a4;
    11'b00100010010: data <= 32'h33503d0e;
    11'b00100010011: data <= 32'ha9a1406b;
    11'b00100010100: data <= 32'hb61b3c5b;
    11'b00100010101: data <= 32'h31e0bd70;
    11'b00100010110: data <= 32'h3d03c0f0;
    11'b00100010111: data <= 32'h3db1bd46;
    11'b00100011000: data <= 32'h38ca329c;
    11'b00100011001: data <= 32'h34133568;
    11'b00100011010: data <= 32'h3b37b546;
    11'b00100011011: data <= 32'h3bb0b684;
    11'b00100011100: data <= 32'hb9f5abfb;
    11'b00100011101: data <= 32'hc163b59a;
    11'b00100011110: data <= 32'hc101bc50;
    11'b00100011111: data <= 32'hb5febc39;
    11'b00100100000: data <= 32'h3c54b26a;
    11'b00100100001: data <= 32'h37ea34b5;
    11'b00100100010: data <= 32'hb9523012;
    11'b00100100011: data <= 32'hb9333826;
    11'b00100100100: data <= 32'h2be53fbd;
    11'b00100100101: data <= 32'h26ff416a;
    11'b00100100110: data <= 32'hb8ff3d39;
    11'b00100100111: data <= 32'hb87dbc23;
    11'b00100101000: data <= 32'h36b2bebf;
    11'b00100101001: data <= 32'h3c93b425;
    11'b00100101010: data <= 32'h3c943bbf;
    11'b00100101011: data <= 32'h3d153718;
    11'b00100101100: data <= 32'h3f17b90f;
    11'b00100101101: data <= 32'h3dabb83f;
    11'b00100101110: data <= 32'hb6c034a0;
    11'b00100101111: data <= 32'hc02f30fd;
    11'b00100110000: data <= 32'hbe8dbc2c;
    11'b00100110001: data <= 32'h3402bf35;
    11'b00100110010: data <= 32'h3c1cbdb1;
    11'b00100110011: data <= 32'hae9bba29;
    11'b00100110100: data <= 32'hbcd2b687;
    11'b00100110101: data <= 32'hb9a03551;
    11'b00100110110: data <= 32'h34b73ea5;
    11'b00100110111: data <= 32'hac6c406c;
    11'b00100111000: data <= 32'hbdb83ba5;
    11'b00100111001: data <= 32'hbf49ba39;
    11'b00100111010: data <= 32'hb933baad;
    11'b00100111011: data <= 32'h39a83911;
    11'b00100111100: data <= 32'h3ce43d70;
    11'b00100111101: data <= 32'h3da23613;
    11'b00100111110: data <= 32'h3edfb88e;
    11'b00100111111: data <= 32'h3d96306d;
    11'b00101000000: data <= 32'h25543da4;
    11'b00101000001: data <= 32'hbc683c53;
    11'b00101000010: data <= 32'hb878ba9e;
    11'b00101000011: data <= 32'h3aa7c073;
    11'b00101000100: data <= 32'h3c06bff7;
    11'b00101000101: data <= 32'hb32dbc7e;
    11'b00101000110: data <= 32'hbadcb948;
    11'b00101000111: data <= 32'h2f5db2a8;
    11'b00101001000: data <= 32'h3be33977;
    11'b00101001001: data <= 32'hae223c9c;
    11'b00101001010: data <= 32'hc05c361b;
    11'b00101001011: data <= 32'hc189b94e;
    11'b00101001100: data <= 32'hbd3cb6f1;
    11'b00101001101: data <= 32'h353539ad;
    11'b00101001110: data <= 32'h39ef3b8e;
    11'b00101001111: data <= 32'h38dda9cf;
    11'b00101010000: data <= 32'h3addb5e3;
    11'b00101010001: data <= 32'h3c043c5b;
    11'b00101010010: data <= 32'h357c4134;
    11'b00101010011: data <= 32'hb6373fa3;
    11'b00101010100: data <= 32'hac45b7a9;
    11'b00101010101: data <= 32'h3a7bbfef;
    11'b00101010110: data <= 32'h3a7dbe1c;
    11'b00101010111: data <= 32'h2868b8ae;
    11'b00101011000: data <= 32'h2e5eb846;
    11'b00101011001: data <= 32'h3d65ba3b;
    11'b00101011010: data <= 32'h3f4fb502;
    11'b00101011011: data <= 32'h2e123578;
    11'b00101011100: data <= 32'hc09d301c;
    11'b00101011101: data <= 32'hc185b8ad;
    11'b00101011110: data <= 32'hbc9cb8e7;
    11'b00101011111: data <= 32'h3258abe1;
    11'b00101100000: data <= 32'ha1b4afd1;
    11'b00101100001: data <= 32'hb88bb9fb;
    11'b00101100010: data <= 32'hb01cb557;
    11'b00101100011: data <= 32'h39313e6f;
    11'b00101100100: data <= 32'h378d4224;
    11'b00101100101: data <= 32'hb5854040;
    11'b00101100110: data <= 32'hb81bb1d7;
    11'b00101100111: data <= 32'h2b22bcd1;
    11'b00101101000: data <= 32'h35a3b599;
    11'b00101101001: data <= 32'h34d8368d;
    11'b00101101010: data <= 32'h3b7eb3a5;
    11'b00101101011: data <= 32'h4065bc72;
    11'b00101101100: data <= 32'h40aab999;
    11'b00101101101: data <= 32'h3715363e;
    11'b00101101110: data <= 32'hbebe3842;
    11'b00101101111: data <= 32'hbf2db605;
    11'b00101110000: data <= 32'hb52cbc3e;
    11'b00101110001: data <= 32'h3535bc52;
    11'b00101110010: data <= 32'hb8f4bcb0;
    11'b00101110011: data <= 32'hbd65bd83;
    11'b00101110100: data <= 32'hb7c8b8cf;
    11'b00101110101: data <= 32'h3a0a3d2a;
    11'b00101110110: data <= 32'h383b40fb;
    11'b00101110111: data <= 32'hbac03e6f;
    11'b00101111000: data <= 32'hbe32adaa;
    11'b00101111001: data <= 32'hbbfeb5a4;
    11'b00101111010: data <= 32'hb3033a1c;
    11'b00101111011: data <= 32'h33db3c6b;
    11'b00101111100: data <= 32'h3c06b0dc;
    11'b00101111101: data <= 32'h402abcb5;
    11'b00101111110: data <= 32'h4061b562;
    11'b00101111111: data <= 32'h3a053d12;
    11'b00110000000: data <= 32'hb9963dbf;
    11'b00110000001: data <= 32'hb819196e;
    11'b00110000010: data <= 32'h3876bd33;
    11'b00110000011: data <= 32'h379bbe37;
    11'b00110000100: data <= 32'hbabfbdf2;
    11'b00110000101: data <= 32'hbd34be40;
    11'b00110000110: data <= 32'h2c91bc33;
    11'b00110000111: data <= 32'h3da53501;
    11'b00110001000: data <= 32'h39713cfe;
    11'b00110001001: data <= 32'hbd7e39f5;
    11'b00110001010: data <= 32'hc0c1b11f;
    11'b00110001011: data <= 32'hbe8f300c;
    11'b00110001100: data <= 32'hb8b73c87;
    11'b00110001101: data <= 32'hb2323bbd;
    11'b00110001110: data <= 32'h323ab82d;
    11'b00110001111: data <= 32'h3c40bca0;
    11'b00110010000: data <= 32'h3e1c35de;
    11'b00110010001: data <= 32'h3b0f40a3;
    11'b00110010010: data <= 32'h2ca04086;
    11'b00110010011: data <= 32'h343b364a;
    11'b00110010100: data <= 32'h3aa8bc30;
    11'b00110010101: data <= 32'h35c7bc43;
    11'b00110010110: data <= 32'hba12ba87;
    11'b00110010111: data <= 32'hb8e2bcce;
    11'b00110011000: data <= 32'h3c95bdbe;
    11'b00110011001: data <= 32'h4086b9cb;
    11'b00110011010: data <= 32'h3bac3134;
    11'b00110011011: data <= 32'hbdbf31ba;
    11'b00110011100: data <= 32'hc0a7b226;
    11'b00110011101: data <= 32'hbd852ef4;
    11'b00110011110: data <= 32'hb8343924;
    11'b00110011111: data <= 32'hba442d43;
    11'b00110100000: data <= 32'hbc0cbcf3;
    11'b00110100001: data <= 32'hb1e7bcfd;
    11'b00110100010: data <= 32'h3acd3a3b;
    11'b00110100011: data <= 32'h3af84177;
    11'b00110100100: data <= 32'h342040d0;
    11'b00110100101: data <= 32'h2f163865;
    11'b00110100110: data <= 32'h348eb663;
    11'b00110100111: data <= 32'haeae307c;
    11'b00110101000: data <= 32'hb92636c1;
    11'b00110101001: data <= 32'h2d27b8a9;
    11'b00110101010: data <= 32'h3fb6be6b;
    11'b00110101011: data <= 32'h4173bced;
    11'b00110101100: data <= 32'h3ce3adbb;
    11'b00110101101: data <= 32'hbb433589;
    11'b00110101110: data <= 32'hbd541d53;
    11'b00110101111: data <= 32'hb542b16e;
    11'b00110110000: data <= 32'had98b23f;
    11'b00110110001: data <= 32'hbcdcbb1b;
    11'b00110110010: data <= 32'hbf95bf6e;
    11'b00110110011: data <= 32'hbac7bdf1;
    11'b00110110100: data <= 32'h39833819;
    11'b00110110101: data <= 32'h3b1f403e;
    11'b00110110110: data <= 32'hac3b3ec7;
    11'b00110110111: data <= 32'hb9b635b0;
    11'b00110111000: data <= 32'hb9633469;
    11'b00110111001: data <= 32'hb9843d60;
    11'b00110111010: data <= 32'hb9ce3db2;
    11'b00110111011: data <= 32'h3114b278;
    11'b00110111100: data <= 32'h3f1fbe68;
    11'b00110111101: data <= 32'h40d8bc28;
    11'b00110111110: data <= 32'h3d1c3869;
    11'b00110111111: data <= 32'hada53c85;
    11'b00111000000: data <= 32'h28063692;
    11'b00111000001: data <= 32'h3adeb566;
    11'b00111000010: data <= 32'h360ab918;
    11'b00111000011: data <= 32'hbd5dbcb1;
    11'b00111000100: data <= 32'hc005bfaf;
    11'b00111000101: data <= 32'hb861bee6;
    11'b00111000110: data <= 32'h3cc9b50d;
    11'b00111000111: data <= 32'h3c453a72;
    11'b00111001000: data <= 32'hb7d1383d;
    11'b00111001001: data <= 32'hbde2a9c7;
    11'b00111001010: data <= 32'hbd21390f;
    11'b00111001011: data <= 32'hbbdb3f76;
    11'b00111001100: data <= 32'hbc083e43;
    11'b00111001101: data <= 32'hb837b643;
    11'b00111001110: data <= 32'h3994be63;
    11'b00111001111: data <= 32'h3de6b778;
    11'b00111010000: data <= 32'h3c4c3dfc;
    11'b00111010001: data <= 32'h38553fac;
    11'b00111010010: data <= 32'h3ba43a18;
    11'b00111010011: data <= 32'h3dbbb1e6;
    11'b00111010100: data <= 32'h37acb3c8;
    11'b00111010101: data <= 32'hbd04b72a;
    11'b00111010110: data <= 32'hbdddbd35;
    11'b00111010111: data <= 32'h3638bf27;
    11'b00111011000: data <= 32'h3fffbcce;
    11'b00111011001: data <= 32'h3d5ab6ba;
    11'b00111011010: data <= 32'hb8ccb5b0;
    11'b00111011011: data <= 32'hbdeeb54a;
    11'b00111011100: data <= 32'hbbd338b7;
    11'b00111011101: data <= 32'hb9933e22;
    11'b00111011110: data <= 32'hbd343acb;
    11'b00111011111: data <= 32'hbe53bc2c;
    11'b00111100000: data <= 32'hb975bece;
    11'b00111100001: data <= 32'h3770aadd;
    11'b00111100010: data <= 32'h3a333fc2;
    11'b00111100011: data <= 32'h3967400f;
    11'b00111100100: data <= 32'h3bbb39e9;
    11'b00111100101: data <= 32'h3c5a3284;
    11'b00111100110: data <= 32'h2e7d3a8a;
    11'b00111100111: data <= 32'hbca93b4d;
    11'b00111101000: data <= 32'hba81b58f;
    11'b00111101001: data <= 32'h3cb1be92;
    11'b00111101010: data <= 32'h40e1be86;
    11'b00111101011: data <= 32'h3dddbabe;
    11'b00111101100: data <= 32'hb495b6d5;
    11'b00111101101: data <= 32'hb8f1b411;
    11'b00111101110: data <= 32'h31ea356c;
    11'b00111101111: data <= 32'h2c6e3a23;
    11'b00111110000: data <= 32'hbd9fae09;
    11'b00111110001: data <= 32'hc0bbbe98;
    11'b00111110010: data <= 32'hbe12bf65;
    11'b00111110011: data <= 32'h27acb0cd;
    11'b00111110100: data <= 32'h390f3dc6;
    11'b00111110101: data <= 32'h35ec3cdf;
    11'b00111110110: data <= 32'h33be338c;
    11'b00111110111: data <= 32'h320f3869;
    11'b00111111000: data <= 32'hb78d3fa4;
    11'b00111111001: data <= 32'hbcc9402e;
    11'b00111111010: data <= 32'hb8e3356a;
    11'b00111111011: data <= 32'h3c7dbdbe;
    11'b00111111100: data <= 32'h401dbdc2;
    11'b00111111101: data <= 32'h3cf7b533;
    11'b00111111110: data <= 32'h3301342d;
    11'b00111111111: data <= 32'h390b302f;
    11'b01000000000: data <= 32'h3e3130e9;
    11'b01000000001: data <= 32'h3aea33e8;
    11'b01000000010: data <= 32'hbd27b756;
    11'b01000000011: data <= 32'hc0ecbea0;
    11'b01000000100: data <= 32'hbd71bf62;
    11'b01000000101: data <= 32'h366db97c;
    11'b01000000110: data <= 32'h3a2733c4;
    11'b01000000111: data <= 32'haa34afa7;
    11'b01000001000: data <= 32'hb869b819;
    11'b01000001001: data <= 32'hb7b03914;
    11'b01000001010: data <= 32'hb9da40cb;
    11'b01000001011: data <= 32'hbd2240c8;
    11'b01000001100: data <= 32'hbc23353c;
    11'b01000001101: data <= 32'h30ebbd70;
    11'b01000001110: data <= 32'h3b90bb0c;
    11'b01000001111: data <= 32'h397938f5;
    11'b01000010000: data <= 32'h386a3c58;
    11'b01000010001: data <= 32'h3e05377e;
    11'b01000010010: data <= 32'h4099310b;
    11'b01000010011: data <= 32'h3cc036a3;
    11'b01000010100: data <= 32'hbc6230e9;
    11'b01000010101: data <= 32'hbfbabb1f;
    11'b01000010110: data <= 32'hb74bbe3f;
    11'b01000010111: data <= 32'h3cdbbd0b;
    11'b01000011000: data <= 32'h3c25bb64;
    11'b01000011001: data <= 32'hb43ebccd;
    11'b01000011010: data <= 32'hba00bc41;
    11'b01000011011: data <= 32'hb4903722;
    11'b01000011100: data <= 32'hb5334026;
    11'b01000011101: data <= 32'hbd003ef2;
    11'b01000011110: data <= 32'hbf1cb4d9;
    11'b01000011111: data <= 32'hbca0bdd9;
    11'b01000100000: data <= 32'hb45eb659;
    11'b01000100001: data <= 32'h2d033cda;
    11'b01000100010: data <= 32'h38003d34;
    11'b01000100011: data <= 32'h3e1635a4;
    11'b01000100100: data <= 32'h40193410;
    11'b01000100101: data <= 32'h3af53cb3;
    11'b01000100110: data <= 32'hbbf53dc0;
    11'b01000100111: data <= 32'hbcf0346c;
    11'b01000101000: data <= 32'h3719bc51;
    11'b01000101001: data <= 32'h3f01bde0;
    11'b01000101010: data <= 32'h3c66bd60;
    11'b01000101011: data <= 32'hb28cbd9a;
    11'b01000101100: data <= 32'hb152bc5f;
    11'b01000101101: data <= 32'h3a5e3146;
    11'b01000101110: data <= 32'h392f3d23;
    11'b01000101111: data <= 32'hbc0039b0;
    11'b01000110000: data <= 32'hc09fbbf7;
    11'b01000110001: data <= 32'hbfeebe49;
    11'b01000110010: data <= 32'hbaf5b480;
    11'b01000110011: data <= 32'hb3213bcc;
    11'b01000110100: data <= 32'h3056389d;
    11'b01000110101: data <= 32'h3a4bb57f;
    11'b01000110110: data <= 32'h3c6a33d9;
    11'b01000110111: data <= 32'h33333ffe;
    11'b01000111000: data <= 32'hbc0a4132;
    11'b01000111001: data <= 32'hbae13c9d;
    11'b01000111010: data <= 32'h3907b948;
    11'b01000111011: data <= 32'h3ddabcba;
    11'b01000111100: data <= 32'h39a0ba99;
    11'b01000111101: data <= 32'ha9eeb9a3;
    11'b01000111110: data <= 32'h3a6db94d;
    11'b01000111111: data <= 32'h4046a608;
    11'b01001000000: data <= 32'h3ea13908;
    11'b01001000001: data <= 32'hb900304f;
    11'b01001000010: data <= 32'hc08bbc6e;
    11'b01001000011: data <= 32'hbf50bdb4;
    11'b01001000100: data <= 32'hb83fb7d3;
    11'b01001000101: data <= 32'hacfe2adf;
    11'b01001000110: data <= 32'hb491b9e2;
    11'b01001000111: data <= 32'haf02bd4a;
    11'b01001001000: data <= 32'h33f427f0;
    11'b01001001001: data <= 32'hb0bb40a3;
    11'b01001001010: data <= 32'hbbe841d0;
    11'b01001001011: data <= 32'hbbdd3cde;
    11'b01001001100: data <= 32'hac0cb85e;
    11'b01001001101: data <= 32'h3628b8de;
    11'b01001001110: data <= 32'hadd7324d;
    11'b01001001111: data <= 32'ha9023470;
    11'b01001010000: data <= 32'h3df0b2b6;
    11'b01001010001: data <= 32'h41ceae01;
    11'b01001010010: data <= 32'h4032383c;
    11'b01001010011: data <= 32'hb57d379b;
    11'b01001010100: data <= 32'hbed5b63a;
    11'b01001010101: data <= 32'hbaefbb46;
    11'b01001010110: data <= 32'h367bb9c5;
    11'b01001010111: data <= 32'h34c1bb30;
    11'b01001011000: data <= 32'hb863bf57;
    11'b01001011001: data <= 32'hb853c011;
    11'b01001011010: data <= 32'h31cfb4cb;
    11'b01001011011: data <= 32'h32273fbf;
    11'b01001011100: data <= 32'hb9ee406c;
    11'b01001011101: data <= 32'hbd8237ff;
    11'b01001011110: data <= 32'hbc92b9e9;
    11'b01001011111: data <= 32'hbadaae23;
    11'b01001100000: data <= 32'hbb2c3beb;
    11'b01001100001: data <= 32'hb48e39ef;
    11'b01001100010: data <= 32'h3da9b3aa;
    11'b01001100011: data <= 32'h4143b1e2;
    11'b01001100100: data <= 32'h3ef13b98;
    11'b01001100101: data <= 32'hb4e33e11;
    11'b01001100110: data <= 32'hbbec3a62;
    11'b01001100111: data <= 32'h328ab250;
    11'b01001101000: data <= 32'h3cb6b980;
    11'b01001101001: data <= 32'h376abcd4;
    11'b01001101010: data <= 32'hb923c011;
    11'b01001101011: data <= 32'hb47ec022;
    11'b01001101100: data <= 32'h3c0cb870;
    11'b01001101101: data <= 32'h3cb43c80;
    11'b01001101110: data <= 32'hb3da3c29;
    11'b01001101111: data <= 32'hbe86b697;
    11'b01001110000: data <= 32'hbf54bbb6;
    11'b01001110001: data <= 32'hbde33092;
    11'b01001110010: data <= 32'hbd063c38;
    11'b01001110011: data <= 32'hb95c345e;
    11'b01001110100: data <= 32'h393abb74;
    11'b01001110101: data <= 32'h3e42b70e;
    11'b01001110110: data <= 32'h3b283ddd;
    11'b01001110111: data <= 32'hb715410a;
    11'b01001111000: data <= 32'hb8293ed6;
    11'b01001111001: data <= 32'h39603557;
    11'b01001111010: data <= 32'h3c99b53a;
    11'b01001111011: data <= 32'h2dcfb92e;
    11'b01001111100: data <= 32'hb9cabcfb;
    11'b01001111101: data <= 32'h35e8bde5;
    11'b01001111110: data <= 32'h405cb900;
    11'b01001111111: data <= 32'h4076365b;
    11'b01010000000: data <= 32'h34a43278;
    11'b01010000001: data <= 32'hbdddba50;
    11'b01010000010: data <= 32'hbe7bbaed;
    11'b01010000011: data <= 32'hbc46310c;
    11'b01010000100: data <= 32'hbbee3758;
    11'b01010000101: data <= 32'hbbecbacf;
    11'b01010000110: data <= 32'hb4c5bfda;
    11'b01010000111: data <= 32'h3783bad4;
    11'b01010001000: data <= 32'h340e3e72;
    11'b01010001001: data <= 32'hb7eb4181;
    11'b01010001010: data <= 32'hb7193ef4;
    11'b01010001011: data <= 32'h34e23611;
    11'b01010001100: data <= 32'h346331a5;
    11'b01010001101: data <= 32'hba0c36bb;
    11'b01010001110: data <= 32'hbb8caa2e;
    11'b01010001111: data <= 32'h3ab3ba0f;
    11'b01010010000: data <= 32'h41b6b8c6;
    11'b01010010001: data <= 32'h41563006;
    11'b01010010010: data <= 32'h38793314;
    11'b01010010011: data <= 32'hbb74b4a8;
    11'b01010010100: data <= 32'hb8e9b4ed;
    11'b01010010101: data <= 32'h2b1d316a;
    11'b01010010110: data <= 32'hb5e1b3f0;
    11'b01010010111: data <= 32'hbc8ebf66;
    11'b01010011000: data <= 32'hbafdc166;
    11'b01010011001: data <= 32'h2da4bce9;
    11'b01010011010: data <= 32'h35a93cdd;
    11'b01010011011: data <= 32'hb3434005;
    11'b01010011100: data <= 32'hb8b73ae5;
    11'b01010011101: data <= 32'hb808a8b3;
    11'b01010011110: data <= 32'hbad43891;
    11'b01010011111: data <= 32'hbe733d57;
    11'b01010100000: data <= 32'hbd2639c2;
    11'b01010100001: data <= 32'h39adb83b;
    11'b01010100010: data <= 32'h4110b970;
    11'b01010100011: data <= 32'h405b34dd;
    11'b01010100100: data <= 32'h368c3bc8;
    11'b01010100101: data <= 32'hb52c3a21;
    11'b01010100110: data <= 32'h38803798;
    11'b01010100111: data <= 32'h3c7b359d;
    11'b01010101000: data <= 32'h2c84b74a;
    11'b01010101001: data <= 32'hbcc8bffb;
    11'b01010101010: data <= 32'hbab7c14b;
    11'b01010101011: data <= 32'h38eebd5c;
    11'b01010101100: data <= 32'h3cc037f1;
    11'b01010101101: data <= 32'h358839f3;
    11'b01010101110: data <= 32'hb93eb53b;
    11'b01010101111: data <= 32'hbc35b852;
    11'b01010110000: data <= 32'hbda739fa;
    11'b01010110001: data <= 32'hbfb63e6e;
    11'b01010110010: data <= 32'hbe55387f;
    11'b01010110011: data <= 32'h22d2bc31;
    11'b01010110100: data <= 32'h3d85bc08;
    11'b01010110101: data <= 32'h3c5238da;
    11'b01010110110: data <= 32'h9eaf3f31;
    11'b01010110111: data <= 32'h2c153e79;
    11'b01010111000: data <= 32'h3ce13c03;
    11'b01010111001: data <= 32'h3da33974;
    11'b01010111010: data <= 32'haea52c88;
    11'b01010111011: data <= 32'hbd55bc86;
    11'b01010111100: data <= 32'hb6b0bf49;
    11'b01010111101: data <= 32'h3e4fbc92;
    11'b01010111110: data <= 32'h405ab058;
    11'b01010111111: data <= 32'h3b51b451;
    11'b01011000000: data <= 32'hb764bc1d;
    11'b01011000001: data <= 32'hbab1b957;
    11'b01011000010: data <= 32'hbb913a5e;
    11'b01011000011: data <= 32'hbde03cfa;
    11'b01011000100: data <= 32'hbea5b54c;
    11'b01011000101: data <= 32'hbab6c001;
    11'b01011000110: data <= 32'h2fe8bdec;
    11'b01011000111: data <= 32'h2f0b395f;
    11'b01011001000: data <= 32'hb4f93ff6;
    11'b01011001001: data <= 32'h30c33e5e;
    11'b01011001010: data <= 32'h3c593b31;
    11'b01011001011: data <= 32'h3a4d3bdc;
    11'b01011001100: data <= 32'hbadc3c2f;
    11'b01011001101: data <= 32'hbe8432d1;
    11'b01011001110: data <= 32'hacbeba3a;
    11'b01011001111: data <= 32'h405bbab9;
    11'b01011010000: data <= 32'h4122b638;
    11'b01011010001: data <= 32'h3c53b7b4;
    11'b01011010010: data <= 32'had2fba77;
    11'b01011010011: data <= 32'h2e06b339;
    11'b01011010100: data <= 32'h34fc3b20;
    11'b01011010101: data <= 32'hb8413992;
    11'b01011010110: data <= 32'hbe19bce8;
    11'b01011010111: data <= 32'hbd7cc166;
    11'b01011011000: data <= 32'hb7b9bf33;
    11'b01011011001: data <= 32'hadd73605;
    11'b01011011010: data <= 32'hb2103d35;
    11'b01011011011: data <= 32'h2d4138c6;
    11'b01011011100: data <= 32'h376c322a;
    11'b01011011101: data <= 32'hb2b13c5f;
    11'b01011011110: data <= 32'hbeba3f9a;
    11'b01011011111: data <= 32'hbfda3ccb;
    11'b01011100000: data <= 32'hb0eab344;
    11'b01011100001: data <= 32'h3f8bb9ee;
    11'b01011100010: data <= 32'h3fe6b466;
    11'b01011100011: data <= 32'h39622c24;
    11'b01011100100: data <= 32'h34262dab;
    11'b01011100101: data <= 32'h3ccf382f;
    11'b01011100110: data <= 32'h3e573c67;
    11'b01011100111: data <= 32'h33d937db;
    11'b01011101000: data <= 32'hbd75bd86;
    11'b01011101001: data <= 32'hbd85c120;
    11'b01011101010: data <= 32'hb18dbec6;
    11'b01011101011: data <= 32'h3867ae85;
    11'b01011101100: data <= 32'h35672e9b;
    11'b01011101101: data <= 32'h2cc5ba59;
    11'b01011101110: data <= 32'ha86db946;
    11'b01011101111: data <= 32'hba0b3c18;
    11'b01011110000: data <= 32'hbfbf4063;
    11'b01011110001: data <= 32'hc02d3d12;
    11'b01011110010: data <= 32'hb926b829;
    11'b01011110011: data <= 32'h3a5fbc01;
    11'b01011110100: data <= 32'h3978a9fa;
    11'b01011110101: data <= 32'haddf3a65;
    11'b01011110110: data <= 32'h361a3b3b;
    11'b01011110111: data <= 32'h3f733c0e;
    11'b01011111000: data <= 32'h40383d42;
    11'b01011111001: data <= 32'h35483ad4;
    11'b01011111010: data <= 32'hbd9db893;
    11'b01011111011: data <= 32'hbc24be41;
    11'b01011111100: data <= 32'h394fbca1;
    11'b01011111101: data <= 32'h3de8b75a;
    11'b01011111110: data <= 32'h3b15bb31;
    11'b01011111111: data <= 32'h3274bef3;
    11'b01100000000: data <= 32'h2c12bc50;
    11'b01100000001: data <= 32'hb55b3b88;
    11'b01100000010: data <= 32'hbd503f9d;
    11'b01100000011: data <= 32'hbf683834;
    11'b01100000100: data <= 32'hbce3bd88;
    11'b01100000101: data <= 32'hb705bdd6;
    11'b01100000110: data <= 32'hb8462922;
    11'b01100000111: data <= 32'hb9c13c3f;
    11'b01100001000: data <= 32'h34cf3b4f;
    11'b01100001001: data <= 32'h3f2d3a50;
    11'b01100001010: data <= 32'h3ea73d58;
    11'b01100001011: data <= 32'hb4d43e46;
    11'b01100001100: data <= 32'hbebb39f3;
    11'b01100001101: data <= 32'hb9a2b459;
    11'b01100001110: data <= 32'h3d2bb80c;
    11'b01100001111: data <= 32'h3f8fb81a;
    11'b01100010000: data <= 32'h3bb2bca8;
    11'b01100010001: data <= 32'h359abede;
    11'b01100010010: data <= 32'h3a12ba5c;
    11'b01100010011: data <= 32'h3b1f3c06;
    11'b01100010100: data <= 32'hb0c13d91;
    11'b01100010101: data <= 32'hbd67b5c2;
    11'b01100010110: data <= 32'hbe1bc02f;
    11'b01100010111: data <= 32'hbc5abede;
    11'b01100011000: data <= 32'hbbafac98;
    11'b01100011001: data <= 32'hba63389d;
    11'b01100011010: data <= 32'h31d4aa19;
    11'b01100011011: data <= 32'h3ce5b098;
    11'b01100011100: data <= 32'h39b03c56;
    11'b01100011101: data <= 32'hbc7e405a;
    11'b01100011110: data <= 32'hbfeb3f0c;
    11'b01100011111: data <= 32'hb9303837;
    11'b01100100000: data <= 32'h3cacb125;
    11'b01100100001: data <= 32'h3d54b511;
    11'b01100100010: data <= 32'h3598b974;
    11'b01100100011: data <= 32'h3578bb34;
    11'b01100100100: data <= 32'h3e75ac6f;
    11'b01100100101: data <= 32'h40603ccd;
    11'b01100100110: data <= 32'h3b253c62;
    11'b01100100111: data <= 32'hbb38b932;
    11'b01100101000: data <= 32'hbdabbffa;
    11'b01100101001: data <= 32'hbac3bdbf;
    11'b01100101010: data <= 32'hb6f9b346;
    11'b01100101011: data <= 32'hb52fb5f8;
    11'b01100101100: data <= 32'h315bbdd4;
    11'b01100101101: data <= 32'h3967bd15;
    11'b01100101110: data <= 32'h2be63988;
    11'b01100101111: data <= 32'hbdae40a2;
    11'b01100110000: data <= 32'hbfdd3f97;
    11'b01100110001: data <= 32'hbace362f;
    11'b01100110010: data <= 32'h3511b546;
    11'b01100110011: data <= 32'h2735acf8;
    11'b01100110100: data <= 32'hb98d2c6e;
    11'b01100110101: data <= 32'h2f7da42b;
    11'b01100110110: data <= 32'h40303774;
    11'b01100110111: data <= 32'h418e3d3f;
    11'b01100111000: data <= 32'h3caa3cd8;
    11'b01100111001: data <= 32'hba70ac03;
    11'b01100111010: data <= 32'hbc30bbe8;
    11'b01100111011: data <= 32'ha474b905;
    11'b01100111100: data <= 32'h3830b332;
    11'b01100111101: data <= 32'h3433bcb4;
    11'b01100111110: data <= 32'h334dc0ef;
    11'b01100111111: data <= 32'h3892bfa7;
    11'b01101000000: data <= 32'h347636ce;
    11'b01101000001: data <= 32'hba8a3fe9;
    11'b01101000010: data <= 32'hbde43cba;
    11'b01101000011: data <= 32'hbc45b792;
    11'b01101000100: data <= 32'hb9a7ba80;
    11'b01101000101: data <= 32'hbd092a39;
    11'b01101000110: data <= 32'hbe4f37d8;
    11'b01101000111: data <= 32'hb23b31a0;
    11'b01101001000: data <= 32'h3fcd3435;
    11'b01101001001: data <= 32'h40be3c6e;
    11'b01101001010: data <= 32'h389b3e50;
    11'b01101001011: data <= 32'hbc573c22;
    11'b01101001100: data <= 32'hb98835f3;
    11'b01101001101: data <= 32'h39d834e8;
    11'b01101001110: data <= 32'h3c629b5f;
    11'b01101001111: data <= 32'h3604bd5d;
    11'b01101010000: data <= 32'h31fbc101;
    11'b01101010001: data <= 32'h3b8abeda;
    11'b01101010010: data <= 32'h3d22375d;
    11'b01101010011: data <= 32'h36c73dc9;
    11'b01101010100: data <= 32'hb96332b6;
    11'b01101010101: data <= 32'hbc3ebd44;
    11'b01101010110: data <= 32'hbcecbc79;
    11'b01101010111: data <= 32'hbf072d9f;
    11'b01101011000: data <= 32'hbf2534c1;
    11'b01101011001: data <= 32'hb622b88d;
    11'b01101011010: data <= 32'h3d6fb9c2;
    11'b01101011011: data <= 32'h3d73386e;
    11'b01101011100: data <= 32'hb5a93f65;
    11'b01101011101: data <= 32'hbdbf3f9e;
    11'b01101011110: data <= 32'hb8293d06;
    11'b01101011111: data <= 32'h3aea3aa6;
    11'b01101100000: data <= 32'h39fd34f6;
    11'b01101100001: data <= 32'hb453ba9c;
    11'b01101100010: data <= 32'haf1bbea0;
    11'b01101100011: data <= 32'h3dcdbb46;
    11'b01101100100: data <= 32'h40d639a9;
    11'b01101100101: data <= 32'h3e3f3c44;
    11'b01101100110: data <= 32'h8b27b4df;
    11'b01101100111: data <= 32'hba45bdaf;
    11'b01101101000: data <= 32'hbb86ba96;
    11'b01101101001: data <= 32'hbceb326c;
    11'b01101101010: data <= 32'hbd18b4ef;
    11'b01101101011: data <= 32'hb5b2bf38;
    11'b01101101100: data <= 32'h39ffbfcc;
    11'b01101101101: data <= 32'h3828ae72;
    11'b01101101110: data <= 32'hbac73f18;
    11'b01101101111: data <= 32'hbdb93fe6;
    11'b01101110000: data <= 32'hb7b73c91;
    11'b01101110001: data <= 32'h358d3960;
    11'b01101110010: data <= 32'hb604383f;
    11'b01101110011: data <= 32'hbdaaa7ee;
    11'b01101110100: data <= 32'hb8ffb8e2;
    11'b01101110101: data <= 32'h3eb4b201;
    11'b01101110110: data <= 32'h41d93ace;
    11'b01101110111: data <= 32'h3f8c3bce;
    11'b01101111000: data <= 32'h311ca8bc;
    11'b01101111001: data <= 32'hb653b8d0;
    11'b01101111010: data <= 32'haccc2d4b;
    11'b01101111011: data <= 32'hb082380e;
    11'b01101111100: data <= 32'hb823ba9c;
    11'b01101111101: data <= 32'hb3d1c170;
    11'b01101111110: data <= 32'h3798c156;
    11'b01101111111: data <= 32'h36fcb7bd;
    11'b01110000000: data <= 32'hb7073d7e;
    11'b01110000001: data <= 32'hbada3ce1;
    11'b01110000010: data <= 32'hb64931e9;
    11'b01110000011: data <= 32'hb5ed29d0;
    11'b01110000100: data <= 32'hbe3938c7;
    11'b01110000101: data <= 32'hc0cd3837;
    11'b01110000110: data <= 32'hbc6bb080;
    11'b01110000111: data <= 32'h3db3b1fa;
    11'b01110001000: data <= 32'h40f238b5;
    11'b01110001001: data <= 32'h3ced3c2d;
    11'b01110001010: data <= 32'hb35339ee;
    11'b01110001011: data <= 32'hae223921;
    11'b01110001100: data <= 32'h3a443c8e;
    11'b01110001101: data <= 32'h397b3b8f;
    11'b01110001110: data <= 32'hb231babb;
    11'b01110001111: data <= 32'hb504c168;
    11'b01110010000: data <= 32'h388dc0e1;
    11'b01110010001: data <= 32'h3c78b623;
    11'b01110010010: data <= 32'h39603b11;
    11'b01110010011: data <= 32'h2cda3100;
    11'b01110010100: data <= 32'hb020bb1b;
    11'b01110010101: data <= 32'hb9a4b78b;
    11'b01110010110: data <= 32'hc0003917;
    11'b01110010111: data <= 32'hc13d38aa;
    11'b01110011000: data <= 32'hbd1db883;
    11'b01110011001: data <= 32'h3accbc19;
    11'b01110011010: data <= 32'h3d8aae2b;
    11'b01110011011: data <= 32'h2e473c1f;
    11'b01110011100: data <= 32'hba4b3d8d;
    11'b01110011101: data <= 32'h2a973de1;
    11'b01110011110: data <= 32'h3c8c3edb;
    11'b01110011111: data <= 32'h39373d34;
    11'b01110100000: data <= 32'hb96db4ff;
    11'b01110100001: data <= 32'hb9d8bf28;
    11'b01110100010: data <= 32'h3a3bbdd8;
    11'b01110100011: data <= 32'h40002b46;
    11'b01110100100: data <= 32'h3eff3857;
    11'b01110100101: data <= 32'h3ab3b86b;
    11'b01110100110: data <= 32'h33febd32;
    11'b01110100111: data <= 32'hb5d5b5b0;
    11'b01110101000: data <= 32'hbda93ac6;
    11'b01110101001: data <= 32'hbfe0346b;
    11'b01110101010: data <= 32'hbc54be1e;
    11'b01110101011: data <= 32'h349ac05e;
    11'b01110101100: data <= 32'h35efbaf4;
    11'b01110101101: data <= 32'hb98d3a63;
    11'b01110101110: data <= 32'hbbd23d79;
    11'b01110101111: data <= 32'h312f3d38;
    11'b01110110000: data <= 32'h3b493dd6;
    11'b01110110001: data <= 32'hb2083d8e;
    11'b01110110010: data <= 32'hbefc3703;
    11'b01110110011: data <= 32'hbd86b8bc;
    11'b01110110100: data <= 32'h3a67b738;
    11'b01110110101: data <= 32'h40c2369b;
    11'b01110110110: data <= 32'h400f3683;
    11'b01110110111: data <= 32'h3b9ab881;
    11'b01110111000: data <= 32'h3870ba32;
    11'b01110111001: data <= 32'h37833752;
    11'b01110111010: data <= 32'hb2383d33;
    11'b01110111011: data <= 32'hbb899bbb;
    11'b01110111100: data <= 32'hb9fbc092;
    11'b01110111101: data <= 32'h9bffc1bc;
    11'b01110111110: data <= 32'h2679bd03;
    11'b01110111111: data <= 32'hb8bc36d0;
    11'b01111000000: data <= 32'hb82138fb;
    11'b01111000001: data <= 32'h36583378;
    11'b01111000010: data <= 32'h374838b6;
    11'b01111000011: data <= 32'hbcbd3cf0;
    11'b01111000100: data <= 32'hc1663beb;
    11'b01111000101: data <= 32'hbfa22fd9;
    11'b01111000110: data <= 32'h382db04f;
    11'b01111000111: data <= 32'h3fa634a4;
    11'b01111001000: data <= 32'h3d1c357c;
    11'b01111001001: data <= 32'h35a3ac00;
    11'b01111001010: data <= 32'h39303433;
    11'b01111001011: data <= 32'h3d3b3df2;
    11'b01111001100: data <= 32'h3ade3f4d;
    11'b01111001101: data <= 32'hb4be2c04;
    11'b01111001110: data <= 32'hb930c074;
    11'b01111001111: data <= 32'ha565c11d;
    11'b01111010000: data <= 32'h36bdbbe2;
    11'b01111010001: data <= 32'h34a52f3a;
    11'b01111010010: data <= 32'h362cb6ae;
    11'b01111010011: data <= 32'h3a41bc31;
    11'b01111010100: data <= 32'h3405b400;
    11'b01111010101: data <= 32'hbe3f3c51;
    11'b01111010110: data <= 32'hc1b83c85;
    11'b01111010111: data <= 32'hbfdaa3eb;
    11'b01111011000: data <= 32'h2d78b9c2;
    11'b01111011001: data <= 32'h3abcb59d;
    11'b01111011010: data <= 32'haa4331f2;
    11'b01111011011: data <= 32'hb82a3692;
    11'b01111011100: data <= 32'h38ad3bfe;
    11'b01111011101: data <= 32'h3ee2400c;
    11'b01111011110: data <= 32'h3c6c403b;
    11'b01111011111: data <= 32'hb80c37f6;
    11'b01111100000: data <= 32'hbbfebd47;
    11'b01111100001: data <= 32'h28eebd9e;
    11'b01111100010: data <= 32'h3c62b3d1;
    11'b01111100011: data <= 32'h3d00a02d;
    11'b01111100100: data <= 32'h3c85bca9;
    11'b01111100101: data <= 32'h3c99bef1;
    11'b01111100110: data <= 32'h3862b6e1;
    11'b01111100111: data <= 32'hbbc83cc8;
    11'b01111101000: data <= 32'hc01c3bc2;
    11'b01111101001: data <= 32'hbdf6b9fa;
    11'b01111101010: data <= 32'hb425bef5;
    11'b01111101011: data <= 32'hb254bc79;
    11'b01111101100: data <= 32'hbc72ad8b;
    11'b01111101101: data <= 32'hbc1c3620;
    11'b01111101110: data <= 32'h388f3a8a;
    11'b01111101111: data <= 32'h3e833e96;
    11'b01111110000: data <= 32'h38203fdd;
    11'b01111110001: data <= 32'hbda23c2e;
    11'b01111110010: data <= 32'hbe97aed4;
    11'b01111110011: data <= 32'ha568b027;
    11'b01111110100: data <= 32'h3dac371a;
    11'b01111110101: data <= 32'h3e022161;
    11'b01111110110: data <= 32'h3c9abd2d;
    11'b01111110111: data <= 32'h3d10bde6;
    11'b01111111000: data <= 32'h3cd2321c;
    11'b01111111001: data <= 32'h34243e8e;
    11'b01111111010: data <= 32'hba333a66;
    11'b01111111011: data <= 32'hba85bd9d;
    11'b01111111100: data <= 32'hb5ebc0c1;
    11'b01111111101: data <= 32'hb92abdc4;
    11'b01111111110: data <= 32'hbd26b533;
    11'b01111111111: data <= 32'hba4db31c;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    