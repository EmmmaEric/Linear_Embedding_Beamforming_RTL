
module memory_rom_10(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbd723a8b;
    11'b00000000001: data <= 32'hb98d3750;
    11'b00000000010: data <= 32'h3b22b755;
    11'b00000000011: data <= 32'h3f80ab3c;
    11'b00000000100: data <= 32'h3b663de2;
    11'b00000000101: data <= 32'hba604076;
    11'b00000000110: data <= 32'hbbfa3dec;
    11'b00000000111: data <= 32'h372135c2;
    11'b00000001000: data <= 32'h3d5ab346;
    11'b00000001001: data <= 32'h3857ba11;
    11'b00000001010: data <= 32'hb573be21;
    11'b00000001011: data <= 32'h36c6be57;
    11'b00000001100: data <= 32'h3faeb535;
    11'b00000001101: data <= 32'h3fba3b3f;
    11'b00000001110: data <= 32'h32a73794;
    11'b00000001111: data <= 32'hbd78bbe3;
    11'b00000010000: data <= 32'hbe6bbd65;
    11'b00000010001: data <= 32'hbd05b358;
    11'b00000010010: data <= 32'hbc973699;
    11'b00000010011: data <= 32'hba70b8c9;
    11'b00000010100: data <= 32'h31ebbe9a;
    11'b00000010101: data <= 32'h3a8cb9ae;
    11'b00000010110: data <= 32'h2f063e3a;
    11'b00000010111: data <= 32'hbc134159;
    11'b00000011000: data <= 32'hbb243f36;
    11'b00000011001: data <= 32'h342d3805;
    11'b00000011010: data <= 32'h38942de0;
    11'b00000011011: data <= 32'hb6ad28e8;
    11'b00000011100: data <= 32'hba59b6d8;
    11'b00000011101: data <= 32'h3a57b9be;
    11'b00000011110: data <= 32'h4187ae2b;
    11'b00000011111: data <= 32'h41533945;
    11'b00000100000: data <= 32'h38ea3542;
    11'b00000100001: data <= 32'hbbdfb910;
    11'b00000100010: data <= 32'hbb13b9d6;
    11'b00000100011: data <= 32'hb4618636;
    11'b00000100100: data <= 32'hb681b12c;
    11'b00000100101: data <= 32'hb9d9bee1;
    11'b00000100110: data <= 32'hb4ffc158;
    11'b00000100111: data <= 32'h34d4bd05;
    11'b00000101000: data <= 32'h28f23d19;
    11'b00000101001: data <= 32'hb9f04072;
    11'b00000101010: data <= 32'hbac13c75;
    11'b00000101011: data <= 32'hb62d1fca;
    11'b00000101100: data <= 32'hb907340d;
    11'b00000101101: data <= 32'hbe283a94;
    11'b00000101110: data <= 32'hbd5836fe;
    11'b00000101111: data <= 32'h39e9b4d8;
    11'b00000110000: data <= 32'h4173b051;
    11'b00000110001: data <= 32'h40cc3968;
    11'b00000110010: data <= 32'h36d43b2d;
    11'b00000110011: data <= 32'hb8e33720;
    11'b00000110100: data <= 32'h2f5934a2;
    11'b00000110101: data <= 32'h3abb3671;
    11'b00000110110: data <= 32'h3319b663;
    11'b00000110111: data <= 32'hb98fc045;
    11'b00000111000: data <= 32'hb65cc1bf;
    11'b00000111001: data <= 32'h3917bd7d;
    11'b00000111010: data <= 32'h3abd3a46;
    11'b00000111011: data <= 32'h27773cb3;
    11'b00000111100: data <= 32'hb966ace4;
    11'b00000111101: data <= 32'hbb57b970;
    11'b00000111110: data <= 32'hbdba34b0;
    11'b00000111111: data <= 32'hc0433caa;
    11'b00001000000: data <= 32'hbeb9378a;
    11'b00001000001: data <= 32'h341cb9f6;
    11'b00001000010: data <= 32'h3f4fb8ef;
    11'b00001000011: data <= 32'h3d6439eb;
    11'b00001000100: data <= 32'hb10f3ea3;
    11'b00001000101: data <= 32'hb6573e04;
    11'b00001000110: data <= 32'h3a5a3c6e;
    11'b00001000111: data <= 32'h3d3e3a9a;
    11'b00001001000: data <= 32'h3135ac10;
    11'b00001001001: data <= 32'hbb7fbe32;
    11'b00001001010: data <= 32'hb2a2c04b;
    11'b00001001011: data <= 32'h3df9bc1d;
    11'b00001001100: data <= 32'h3ff935af;
    11'b00001001101: data <= 32'h3b18322f;
    11'b00001001110: data <= 32'hb593bb7e;
    11'b00001001111: data <= 32'hbae1bba0;
    11'b00001010000: data <= 32'hbd08365b;
    11'b00001010001: data <= 32'hbf483c13;
    11'b00001010010: data <= 32'hbe91b48b;
    11'b00001010011: data <= 32'hb5e4bf40;
    11'b00001010100: data <= 32'h3940bd77;
    11'b00001010101: data <= 32'h34003917;
    11'b00001010110: data <= 32'hb90e3fe1;
    11'b00001010111: data <= 32'hb4e73f18;
    11'b00001011000: data <= 32'h3ad03cc7;
    11'b00001011001: data <= 32'h3ad43c2e;
    11'b00001011010: data <= 32'hb93d395d;
    11'b00001011011: data <= 32'hbdf6b586;
    11'b00001011100: data <= 32'habb7bc10;
    11'b00001011101: data <= 32'h4055b854;
    11'b00001011110: data <= 32'h415630c2;
    11'b00001011111: data <= 32'h3d20b1a2;
    11'b00001100000: data <= 32'h9fd3bb32;
    11'b00001100001: data <= 32'hb18ab7f1;
    11'b00001100010: data <= 32'hb20d39c5;
    11'b00001100011: data <= 32'hbab83983;
    11'b00001100100: data <= 32'hbd42bcd3;
    11'b00001100101: data <= 32'hba6ec18d;
    11'b00001100110: data <= 32'hac2bbfc2;
    11'b00001100111: data <= 32'hb09a356a;
    11'b00001101000: data <= 32'hb8593e11;
    11'b00001101001: data <= 32'hb1b93c08;
    11'b00001101010: data <= 32'h375f37ea;
    11'b00001101011: data <= 32'hafe23bc5;
    11'b00001101100: data <= 32'hbedc3d86;
    11'b00001101101: data <= 32'hc03139a4;
    11'b00001101110: data <= 32'hb1edb463;
    11'b00001101111: data <= 32'h402fb5d1;
    11'b00001110000: data <= 32'h40ac2f17;
    11'b00001110001: data <= 32'h3b6c3039;
    11'b00001110010: data <= 32'h3137ac60;
    11'b00001110011: data <= 32'h3a07373d;
    11'b00001110100: data <= 32'h3c613cdc;
    11'b00001110101: data <= 32'h2f293893;
    11'b00001110110: data <= 32'hbc26be36;
    11'b00001110111: data <= 32'hbb52c1d7;
    11'b00001111000: data <= 32'h221bbfbe;
    11'b00001111001: data <= 32'h363d205f;
    11'b00001111010: data <= 32'h307d383e;
    11'b00001111011: data <= 32'h2e42b569;
    11'b00001111100: data <= 32'h2deab80f;
    11'b00001111101: data <= 32'hbaa03a0a;
    11'b00001111110: data <= 32'hc0873ee6;
    11'b00001111111: data <= 32'hc0bc3be9;
    11'b00010000000: data <= 32'hb870b6cf;
    11'b00010000001: data <= 32'h3cf4b9dc;
    11'b00010000010: data <= 32'h3c932c1c;
    11'b00010000011: data <= 32'h29b13996;
    11'b00010000100: data <= 32'h2f6e3ae7;
    11'b00010000101: data <= 32'h3da53cf3;
    11'b00010000110: data <= 32'h3f383e77;
    11'b00010000111: data <= 32'h35ce3ac9;
    11'b00010001000: data <= 32'hbc8bbbf1;
    11'b00010001001: data <= 32'hba9bc024;
    11'b00010001010: data <= 32'h3931bd46;
    11'b00010001011: data <= 32'h3d8ab148;
    11'b00010001100: data <= 32'h3bc3b6af;
    11'b00010001101: data <= 32'h3731bdb9;
    11'b00010001110: data <= 32'h30a7bc6e;
    11'b00010001111: data <= 32'hb9453979;
    11'b00010010000: data <= 32'hbf683ea5;
    11'b00010010001: data <= 32'hc02f377b;
    11'b00010010010: data <= 32'hbb89bd3c;
    11'b00010010011: data <= 32'h2ef1bdce;
    11'b00010010100: data <= 32'hb1bbae7e;
    11'b00010010101: data <= 32'hba273baf;
    11'b00010010110: data <= 32'h14fd3c75;
    11'b00010010111: data <= 32'h3e223cfe;
    11'b00010011000: data <= 32'h3e5d3e95;
    11'b00010011001: data <= 32'hb3c73d7f;
    11'b00010011010: data <= 32'hbe953171;
    11'b00010011011: data <= 32'hba1fb9ca;
    11'b00010011100: data <= 32'h3cedb7bf;
    11'b00010011101: data <= 32'h4009b082;
    11'b00010011110: data <= 32'h3d3fbaa7;
    11'b00010011111: data <= 32'h393bbe95;
    11'b00010100000: data <= 32'h3951bb22;
    11'b00010100001: data <= 32'h35f63b8d;
    11'b00010100010: data <= 32'hb9613db9;
    11'b00010100011: data <= 32'hbdb0b53b;
    11'b00010100100: data <= 32'hbc84c06a;
    11'b00010100101: data <= 32'hb91dbff6;
    11'b00010100110: data <= 32'hbaaab50f;
    11'b00010100111: data <= 32'hbba43907;
    11'b00010101000: data <= 32'h28c43609;
    11'b00010101001: data <= 32'h3cfb35f2;
    11'b00010101010: data <= 32'h3a2c3cfd;
    11'b00010101011: data <= 32'hbcde3f52;
    11'b00010101100: data <= 32'hc0773ced;
    11'b00010101101: data <= 32'hbad93487;
    11'b00010101110: data <= 32'h3cec057c;
    11'b00010101111: data <= 32'h3ed1aae5;
    11'b00010110000: data <= 32'h3a77b8fc;
    11'b00010110001: data <= 32'h3840bbfe;
    11'b00010110010: data <= 32'h3d61aaf7;
    11'b00010110011: data <= 32'h3ea13db6;
    11'b00010110100: data <= 32'h385e3d49;
    11'b00010110101: data <= 32'hba7cb9a1;
    11'b00010110110: data <= 32'hbc51c0b9;
    11'b00010110111: data <= 32'hb938bf77;
    11'b00010111000: data <= 32'hb813b64c;
    11'b00010111001: data <= 32'hb6a1b032;
    11'b00010111010: data <= 32'h34d8bbb8;
    11'b00010111011: data <= 32'h3b5dbb23;
    11'b00010111100: data <= 32'h2ce8396d;
    11'b00010111101: data <= 32'hbf113fed;
    11'b00010111110: data <= 32'hc0d63e5e;
    11'b00010111111: data <= 32'hbc1435d8;
    11'b00011000000: data <= 32'h389bb1fc;
    11'b00011000001: data <= 32'h3823acd0;
    11'b00011000010: data <= 32'hb53cb006;
    11'b00011000011: data <= 32'h3004af70;
    11'b00011000100: data <= 32'h3f2639c6;
    11'b00011000101: data <= 32'h40dd3f19;
    11'b00011000110: data <= 32'h3c343dc6;
    11'b00011000111: data <= 32'hb97db4fa;
    11'b00011001000: data <= 32'hbb85be13;
    11'b00011001001: data <= 32'hae53bc0f;
    11'b00011001010: data <= 32'h3667b2d9;
    11'b00011001011: data <= 32'h3641bad2;
    11'b00011001100: data <= 32'h3905c03a;
    11'b00011001101: data <= 32'h3af6bf0e;
    11'b00011001110: data <= 32'h2f303581;
    11'b00011001111: data <= 32'hbd763f59;
    11'b00011010000: data <= 32'hbfbb3ca4;
    11'b00011010001: data <= 32'hbc49b65f;
    11'b00011010010: data <= 32'hb536badb;
    11'b00011010011: data <= 32'hbadbb36b;
    11'b00011010100: data <= 32'hbdb63227;
    11'b00011010101: data <= 32'hb4a23376;
    11'b00011010110: data <= 32'h3f2f39ff;
    11'b00011010111: data <= 32'h409e3e86;
    11'b00011011000: data <= 32'h38c83ea7;
    11'b00011011001: data <= 32'hbc763906;
    11'b00011011010: data <= 32'hbb01b007;
    11'b00011011011: data <= 32'h37fe2f7b;
    11'b00011011100: data <= 32'h3c623083;
    11'b00011011101: data <= 32'h3a06bc80;
    11'b00011011110: data <= 32'h3998c0d7;
    11'b00011011111: data <= 32'h3c7fbef0;
    11'b00011100000: data <= 32'h3b7637ce;
    11'b00011100001: data <= 32'hb0c13e62;
    11'b00011100010: data <= 32'hbbbb3615;
    11'b00011100011: data <= 32'hbb40bd4d;
    11'b00011100100: data <= 32'hbb43bdab;
    11'b00011100101: data <= 32'hbe6cb5a4;
    11'b00011100110: data <= 32'hbf572d05;
    11'b00011100111: data <= 32'hb698b4fe;
    11'b00011101000: data <= 32'h3df0b0ed;
    11'b00011101001: data <= 32'h3e1b3b97;
    11'b00011101010: data <= 32'hb5f33f09;
    11'b00011101011: data <= 32'hbede3e05;
    11'b00011101100: data <= 32'hbb3e3bd1;
    11'b00011101101: data <= 32'h395c3add;
    11'b00011101110: data <= 32'h3b9c36ec;
    11'b00011101111: data <= 32'h338abafb;
    11'b00011110000: data <= 32'h3514bf53;
    11'b00011110001: data <= 32'h3dcebb7f;
    11'b00011110010: data <= 32'h400b3bc8;
    11'b00011110011: data <= 32'h3ca93dce;
    11'b00011110100: data <= 32'hac4eb004;
    11'b00011110101: data <= 32'hb8d9be80;
    11'b00011110110: data <= 32'hbad0bd2b;
    11'b00011110111: data <= 32'hbd6cb289;
    11'b00011111000: data <= 32'hbd7fb593;
    11'b00011111001: data <= 32'hb159bdd3;
    11'b00011111010: data <= 32'h3c90be09;
    11'b00011111011: data <= 32'h39ed2c99;
    11'b00011111100: data <= 32'hbc2e3e79;
    11'b00011111101: data <= 32'hbfaa3f15;
    11'b00011111110: data <= 32'hbb0c3c98;
    11'b00011111111: data <= 32'h351c3a5e;
    11'b00100000000: data <= 32'ha94b3772;
    11'b00100000001: data <= 32'hbbe0b5cf;
    11'b00100000010: data <= 32'hb67bbb21;
    11'b00100000011: data <= 32'h3e4aabae;
    11'b00100000100: data <= 32'h415b3d63;
    11'b00100000101: data <= 32'h3f173db2;
    11'b00100000110: data <= 32'h33579c84;
    11'b00100000111: data <= 32'hb5e8bbc3;
    11'b00100001000: data <= 32'hb486b5dd;
    11'b00100001001: data <= 32'hb6bf34a2;
    11'b00100001010: data <= 32'hb7f3b9dc;
    11'b00100001011: data <= 32'h3232c0f1;
    11'b00100001100: data <= 32'h3bd7c0fd;
    11'b00100001101: data <= 32'h3852b7ad;
    11'b00100001110: data <= 32'hba9c3d51;
    11'b00100001111: data <= 32'hbd803d3f;
    11'b00100010000: data <= 32'hb90e363b;
    11'b00100010001: data <= 32'hb3aa2db8;
    11'b00100010010: data <= 32'hbd153468;
    11'b00100010011: data <= 32'hc06b2813;
    11'b00100010100: data <= 32'hbc4fb578;
    11'b00100010101: data <= 32'h3d8f309d;
    11'b00100010110: data <= 32'h41063caf;
    11'b00100010111: data <= 32'h3d663d79;
    11'b00100011000: data <= 32'hb23d38c6;
    11'b00100011001: data <= 32'hb5273451;
    11'b00100011010: data <= 32'h35e63b2c;
    11'b00100011011: data <= 32'h37043b7d;
    11'b00100011100: data <= 32'h2824ba2c;
    11'b00100011101: data <= 32'h3421c170;
    11'b00100011110: data <= 32'h3bf0c10c;
    11'b00100011111: data <= 32'h3c24b635;
    11'b00100100000: data <= 32'h33613c50;
    11'b00100100001: data <= 32'hb46e37db;
    11'b00100100010: data <= 32'hb0d0b958;
    11'b00100100011: data <= 32'hb86db8fc;
    11'b00100100100: data <= 32'hbfca3072;
    11'b00100100101: data <= 32'hc1672fba;
    11'b00100100110: data <= 32'hbd36b8a9;
    11'b00100100111: data <= 32'h3c23b8bc;
    11'b00100101000: data <= 32'h3ec735e4;
    11'b00100101001: data <= 32'h34803c8c;
    11'b00100101010: data <= 32'hbb6f3cb7;
    11'b00100101011: data <= 32'hb6213d29;
    11'b00100101100: data <= 32'h39a23f01;
    11'b00100101101: data <= 32'h38973d89;
    11'b00100101110: data <= 32'hb4fcb6f5;
    11'b00100101111: data <= 32'hb327c030;
    11'b00100110000: data <= 32'h3bf9bea2;
    11'b00100110001: data <= 32'h3f403281;
    11'b00100110010: data <= 32'h3dce3bc4;
    11'b00100110011: data <= 32'h3a14b0c0;
    11'b00100110100: data <= 32'h35bebce4;
    11'b00100110101: data <= 32'hb5ecb96b;
    11'b00100110110: data <= 32'hbea635c8;
    11'b00100110111: data <= 32'hc06b91f0;
    11'b00100111000: data <= 32'hbbe5bda1;
    11'b00100111001: data <= 32'h39c9bf60;
    11'b00100111010: data <= 32'h3a66b94c;
    11'b00100111011: data <= 32'hb8fc39ee;
    11'b00100111100: data <= 32'hbd3e3d18;
    11'b00100111101: data <= 32'hb4fe3db2;
    11'b00100111110: data <= 32'h39123eca;
    11'b00100111111: data <= 32'hae933d91;
    11'b00101000000: data <= 32'hbdab2b18;
    11'b00101000001: data <= 32'hbc6cbc43;
    11'b00101000010: data <= 32'h3aa2b899;
    11'b00101000011: data <= 32'h40853a16;
    11'b00101000100: data <= 32'h40093b64;
    11'b00101000101: data <= 32'h3c6cb479;
    11'b00101000110: data <= 32'h3900bb06;
    11'b00101000111: data <= 32'h328e2fda;
    11'b00101001000: data <= 32'hb9413c0b;
    11'b00101001001: data <= 32'hbc9eacd7;
    11'b00101001010: data <= 32'hb72ec05e;
    11'b00101001011: data <= 32'h388ac192;
    11'b00101001100: data <= 32'h3602bd35;
    11'b00101001101: data <= 32'hb9a835d1;
    11'b00101001110: data <= 32'hbb483a33;
    11'b00101001111: data <= 32'h2d1138d8;
    11'b00101010000: data <= 32'h36473ac9;
    11'b00101010001: data <= 32'hbc4b3c2a;
    11'b00101010010: data <= 32'hc13036d9;
    11'b00101010011: data <= 32'hbf9ab527;
    11'b00101010100: data <= 32'h3805acda;
    11'b00101010101: data <= 32'h400839f2;
    11'b00101010110: data <= 32'h3e2d39fc;
    11'b00101010111: data <= 32'h38a21e6f;
    11'b00101011000: data <= 32'h38552db1;
    11'b00101011001: data <= 32'h3a9f3d56;
    11'b00101011010: data <= 32'h35f03f3b;
    11'b00101011011: data <= 32'hb57b2d10;
    11'b00101011100: data <= 32'hb29bc0a4;
    11'b00101011101: data <= 32'h37d2c18a;
    11'b00101011110: data <= 32'h3887bc9c;
    11'b00101011111: data <= 32'h2c203277;
    11'b00101100000: data <= 32'h3013a617;
    11'b00101100001: data <= 32'h39d8b8c6;
    11'b00101100010: data <= 32'h3508b02c;
    11'b00101100011: data <= 32'hbe6e39b5;
    11'b00101100100: data <= 32'hc21c389d;
    11'b00101100101: data <= 32'hc03bb466;
    11'b00101100110: data <= 32'h31f6b822;
    11'b00101100111: data <= 32'h3cd12497;
    11'b00101101000: data <= 32'h3596356f;
    11'b00101101001: data <= 32'hb660351b;
    11'b00101101010: data <= 32'h34933b84;
    11'b00101101011: data <= 32'h3cc84055;
    11'b00101101100: data <= 32'h3a2f4096;
    11'b00101101101: data <= 32'hb62336df;
    11'b00101101110: data <= 32'hb8b5beb8;
    11'b00101101111: data <= 32'h3525bf2f;
    11'b00101110000: data <= 32'h3c35b58b;
    11'b00101110001: data <= 32'h3c5c3484;
    11'b00101110010: data <= 32'h3c9bb968;
    11'b00101110011: data <= 32'h3d4ebd97;
    11'b00101110100: data <= 32'h3888b7dd;
    11'b00101110101: data <= 32'hbd233a7c;
    11'b00101110110: data <= 32'hc0f238de;
    11'b00101110111: data <= 32'hbe7bba65;
    11'b00101111000: data <= 32'h29cabe34;
    11'b00101111001: data <= 32'h34eebc01;
    11'b00101111010: data <= 32'hba44b1e3;
    11'b00101111011: data <= 32'hbc5a34a8;
    11'b00101111100: data <= 32'h329c3c0b;
    11'b00101111101: data <= 32'h3d054018;
    11'b00101111110: data <= 32'h36604056;
    11'b00101111111: data <= 32'hbd023a3b;
    11'b00110000000: data <= 32'hbdcfb93a;
    11'b00110000001: data <= 32'h9905b803;
    11'b00110000010: data <= 32'h3d503824;
    11'b00110000011: data <= 32'h3e473685;
    11'b00110000100: data <= 32'h3dd1bb4a;
    11'b00110000101: data <= 32'h3e0dbd67;
    11'b00110000110: data <= 32'h3c2a2ad4;
    11'b00110000111: data <= 32'hb46c3db6;
    11'b00110001000: data <= 32'hbce739a6;
    11'b00110001001: data <= 32'hba45bd77;
    11'b00110001010: data <= 32'h2cf6c0c3;
    11'b00110001011: data <= 32'hb24bbe7c;
    11'b00110001100: data <= 32'hbca4b850;
    11'b00110001101: data <= 32'hbbb2b0fd;
    11'b00110001110: data <= 32'h385d31d4;
    11'b00110001111: data <= 32'h3cc23c1e;
    11'b00110010000: data <= 32'hb55d3e28;
    11'b00110010001: data <= 32'hc0983ba7;
    11'b00110010010: data <= 32'hc07d30d2;
    11'b00110010011: data <= 32'hb5c4348f;
    11'b00110010100: data <= 32'h3c563a5c;
    11'b00110010101: data <= 32'h3c4b34f5;
    11'b00110010110: data <= 32'h3a4eba60;
    11'b00110010111: data <= 32'h3cbcb922;
    11'b00110011000: data <= 32'h3de63c74;
    11'b00110011001: data <= 32'h3a5d4077;
    11'b00110011010: data <= 32'hb0493b82;
    11'b00110011011: data <= 32'hb34dbdce;
    11'b00110011100: data <= 32'h2ee8c0a9;
    11'b00110011101: data <= 32'hb150bd71;
    11'b00110011110: data <= 32'hb94db7fc;
    11'b00110011111: data <= 32'hae40ba4a;
    11'b00110100000: data <= 32'h3cd7bc37;
    11'b00110100001: data <= 32'h3ce9b2ed;
    11'b00110100010: data <= 32'hba323b16;
    11'b00110100011: data <= 32'hc16b3bba;
    11'b00110100100: data <= 32'hc0c23570;
    11'b00110100101: data <= 32'hb8343039;
    11'b00110100110: data <= 32'h368e3450;
    11'b00110100111: data <= 32'hb0e1aed1;
    11'b00110101000: data <= 32'hb70eb908;
    11'b00110101001: data <= 32'h38cf2cd7;
    11'b00110101010: data <= 32'h3eb83f8c;
    11'b00110101011: data <= 32'h3d474159;
    11'b00110101100: data <= 32'h2fdd3cc5;
    11'b00110101101: data <= 32'hb60fbb4a;
    11'b00110101110: data <= 32'haa5bbd4c;
    11'b00110101111: data <= 32'h310ab52f;
    11'b00110110000: data <= 32'h323aae7d;
    11'b00110110001: data <= 32'h3ad6bd0c;
    11'b00110110010: data <= 32'h3f2cbfd8;
    11'b00110110011: data <= 32'h3dc2bb0e;
    11'b00110110100: data <= 32'hb81739c2;
    11'b00110110101: data <= 32'hc0303bb1;
    11'b00110110110: data <= 32'hbebaa3f6;
    11'b00110110111: data <= 32'hb5f0b9a0;
    11'b00110111000: data <= 32'hb4f1b949;
    11'b00110111001: data <= 32'hbd83b921;
    11'b00110111010: data <= 32'hbdc2b95c;
    11'b00110111011: data <= 32'h335d3155;
    11'b00110111100: data <= 32'h3eb03ef2;
    11'b00110111101: data <= 32'h3c7240c2;
    11'b00110111110: data <= 32'hb8283d1e;
    11'b00110111111: data <= 32'hbc85ab04;
    11'b00111000000: data <= 32'hb6602b14;
    11'b00111000001: data <= 32'h35fc3acd;
    11'b00111000010: data <= 32'h39393569;
    11'b00111000011: data <= 32'h3c85bd9b;
    11'b00111000100: data <= 32'h3f67c025;
    11'b00111000101: data <= 32'h3ec7b8b2;
    11'b00111000110: data <= 32'h357a3cc9;
    11'b00111000111: data <= 32'hba2b3c56;
    11'b00111001000: data <= 32'hb851b7c8;
    11'b00111001001: data <= 32'ha04bbde6;
    11'b00111001010: data <= 32'hb98cbd02;
    11'b00111001011: data <= 32'hbfa3bb4b;
    11'b00111001100: data <= 32'hbe58bb9a;
    11'b00111001101: data <= 32'h3652b840;
    11'b00111001110: data <= 32'h3e7d3937;
    11'b00111001111: data <= 32'h37f93dd6;
    11'b00111010000: data <= 32'hbde33c7c;
    11'b00111010001: data <= 32'hbf8f38e2;
    11'b00111010010: data <= 32'hb9b03bec;
    11'b00111010011: data <= 32'h33ba3db2;
    11'b00111010100: data <= 32'h34253739;
    11'b00111010101: data <= 32'h3685bd24;
    11'b00111010110: data <= 32'h3d07be02;
    11'b00111010111: data <= 32'h3f353590;
    11'b00111011000: data <= 32'h3d0e3fd7;
    11'b00111011001: data <= 32'h376b3d36;
    11'b00111011010: data <= 32'h355ab90c;
    11'b00111011011: data <= 32'h3456bdf9;
    11'b00111011100: data <= 32'hb91bbb95;
    11'b00111011101: data <= 32'hbe3fb924;
    11'b00111011110: data <= 32'hbb07bd1c;
    11'b00111011111: data <= 32'h3c03be76;
    11'b00111100000: data <= 32'h3eadb9d7;
    11'b00111100001: data <= 32'h29cb378f;
    11'b00111100010: data <= 32'hbfb23ac3;
    11'b00111100011: data <= 32'hbff939ff;
    11'b00111100100: data <= 32'hb9843bfa;
    11'b00111100101: data <= 32'hb1513c5c;
    11'b00111100110: data <= 32'hba922f65;
    11'b00111100111: data <= 32'hbb96bc8e;
    11'b00111101000: data <= 32'h355fba7a;
    11'b00111101001: data <= 32'h3ec63c8a;
    11'b00111101010: data <= 32'h3eda40c2;
    11'b00111101011: data <= 32'h3b1a3da8;
    11'b00111101100: data <= 32'h369fb50d;
    11'b00111101101: data <= 32'h3349b8f6;
    11'b00111101110: data <= 32'hb56f328c;
    11'b00111101111: data <= 32'hba1b2d88;
    11'b00111110000: data <= 32'h2b83bdb4;
    11'b00111110001: data <= 32'h3e4bc0da;
    11'b00111110010: data <= 32'h3f20be45;
    11'b00111110011: data <= 32'h301b28fc;
    11'b00111110100: data <= 32'hbdb5397b;
    11'b00111110101: data <= 32'hbcc53693;
    11'b00111110110: data <= 32'hb3103403;
    11'b00111110111: data <= 32'hb875329c;
    11'b00111111000: data <= 32'hbfc2b694;
    11'b00111111001: data <= 32'hc03ebc7d;
    11'b00111111010: data <= 32'hb55fb8ab;
    11'b00111111011: data <= 32'h3df33c59;
    11'b00111111100: data <= 32'h3e054001;
    11'b00111111101: data <= 32'h35bb3cdb;
    11'b00111111110: data <= 32'hb410332b;
    11'b00111111111: data <= 32'haebb392c;
    11'b01000000000: data <= 32'hae4e3e3a;
    11'b01000000001: data <= 32'hb2d53ad4;
    11'b01000000010: data <= 32'h36c5bd50;
    11'b01000000011: data <= 32'h3e4cc10a;
    11'b01000000100: data <= 32'h3f27bda0;
    11'b01000000101: data <= 32'h397b3640;
    11'b01000000110: data <= 32'hb2f43a2e;
    11'b01000000111: data <= 32'h3004ac04;
    11'b01000001000: data <= 32'h37d0b891;
    11'b01000001001: data <= 32'hb961b74a;
    11'b01000001010: data <= 32'hc0dfb930;
    11'b01000001011: data <= 32'hc0d8bccb;
    11'b01000001100: data <= 32'hb56abc0d;
    11'b01000001101: data <= 32'h3d7d2f7f;
    11'b01000001110: data <= 32'h3b323b52;
    11'b01000001111: data <= 32'hb8dc399d;
    11'b01000010000: data <= 32'hbc4038c5;
    11'b01000010001: data <= 32'hb67a3e23;
    11'b01000010010: data <= 32'hacbe409b;
    11'b01000010011: data <= 32'hb5fb3cb7;
    11'b01000010100: data <= 32'hb1f3bc72;
    11'b01000010101: data <= 32'h3aa5bfd5;
    11'b01000010110: data <= 32'h3e2fb7d7;
    11'b01000010111: data <= 32'h3d333cb5;
    11'b01000011000: data <= 32'h3bb03bea;
    11'b01000011001: data <= 32'h3cc6b526;
    11'b01000011010: data <= 32'h3c1aba4b;
    11'b01000011011: data <= 32'hb7a5b434;
    11'b01000011100: data <= 32'hc031b414;
    11'b01000011101: data <= 32'hbf0fbcca;
    11'b01000011110: data <= 32'h342abf26;
    11'b01000011111: data <= 32'h3dadbccc;
    11'b01000100000: data <= 32'h35dfb47a;
    11'b01000100001: data <= 32'hbce13005;
    11'b01000100010: data <= 32'hbd183872;
    11'b01000100011: data <= 32'hb4993e2e;
    11'b01000100100: data <= 32'hb1ee401c;
    11'b01000100101: data <= 32'hbc9d3b22;
    11'b01000100110: data <= 32'hbddfbba7;
    11'b01000100111: data <= 32'hb4dcbcdb;
    11'b01000101000: data <= 32'h3c6c36cc;
    11'b01000101001: data <= 32'h3e213ecd;
    11'b01000101010: data <= 32'h3d873c22;
    11'b01000101011: data <= 32'h3d92b43d;
    11'b01000101100: data <= 32'h3c4fb24e;
    11'b01000101101: data <= 32'hb0dc3a7b;
    11'b01000101110: data <= 32'hbd0f3976;
    11'b01000101111: data <= 32'hb9dabbf6;
    11'b01000110000: data <= 32'h3b69c0b4;
    11'b01000110001: data <= 32'h3df7c00e;
    11'b01000110010: data <= 32'h3361baf2;
    11'b01000110011: data <= 32'hbbe6b1d7;
    11'b01000110100: data <= 32'hb87a312c;
    11'b01000110101: data <= 32'h36073a40;
    11'b01000110110: data <= 32'hb3143c71;
    11'b01000110111: data <= 32'hc003348a;
    11'b01000111000: data <= 32'hc141bb62;
    11'b01000111001: data <= 32'hbca5ba73;
    11'b01000111010: data <= 32'h399438f6;
    11'b01000111011: data <= 32'h3cef3dac;
    11'b01000111100: data <= 32'h3ac43947;
    11'b01000111101: data <= 32'h39a0aca1;
    11'b01000111110: data <= 32'h39833a5d;
    11'b01000111111: data <= 32'h2df04049;
    11'b01001000000: data <= 32'hb8903ea4;
    11'b01001000001: data <= 32'hb0adb92d;
    11'b01001000010: data <= 32'h3c23c0a3;
    11'b01001000011: data <= 32'h3d69bf76;
    11'b01001000100: data <= 32'h3753b84b;
    11'b01001000101: data <= 32'haaf8aceb;
    11'b01001000110: data <= 32'h39e4b506;
    11'b01001000111: data <= 32'h3d41b0e6;
    11'b01001001000: data <= 32'ha9fd3405;
    11'b01001001001: data <= 32'hc0afac8a;
    11'b01001001010: data <= 32'hc1ddbb19;
    11'b01001001011: data <= 32'hbce9bb73;
    11'b01001001100: data <= 32'h3870acb3;
    11'b01001001101: data <= 32'h38eb35c7;
    11'b01001001110: data <= 32'hb2a0adbb;
    11'b01001001111: data <= 32'hb461a50a;
    11'b01001010000: data <= 32'h344c3dfd;
    11'b01001010001: data <= 32'h323a41ce;
    11'b01001010010: data <= 32'hb7534030;
    11'b01001010011: data <= 32'hb7b6b5a0;
    11'b01001010100: data <= 32'h3560bee5;
    11'b01001010101: data <= 32'h3b07bb11;
    11'b01001010110: data <= 32'h39de362d;
    11'b01001010111: data <= 32'h3b543414;
    11'b01001011000: data <= 32'h3f4cb8fb;
    11'b01001011001: data <= 32'h4002b8de;
    11'b01001011010: data <= 32'h347731b0;
    11'b01001011011: data <= 32'hbfc8341d;
    11'b01001011100: data <= 32'hc074b95e;
    11'b01001011101: data <= 32'hb83bbd71;
    11'b01001011110: data <= 32'h3999bca8;
    11'b01001011111: data <= 32'h2a6fbade;
    11'b01001100000: data <= 32'hbc1dbade;
    11'b01001100001: data <= 32'hb9eeb3cb;
    11'b01001100010: data <= 32'h34cb3db4;
    11'b01001100011: data <= 32'h34584140;
    11'b01001100100: data <= 32'hbb2f3eff;
    11'b01001100101: data <= 32'hbe1bb44c;
    11'b01001100110: data <= 32'hba92bba5;
    11'b01001100111: data <= 32'h32d532d5;
    11'b01001101000: data <= 32'h39e03c9d;
    11'b01001101001: data <= 32'h3ced3676;
    11'b01001101010: data <= 32'h4008b9c8;
    11'b01001101011: data <= 32'h4018b57f;
    11'b01001101100: data <= 32'h388f3c03;
    11'b01001101101: data <= 32'hbc5e3cd5;
    11'b01001101110: data <= 32'hbc26b341;
    11'b01001101111: data <= 32'h35ddbe9e;
    11'b01001110000: data <= 32'h3b21bf74;
    11'b01001110001: data <= 32'hb2cdbdd8;
    11'b01001110010: data <= 32'hbc67bcda;
    11'b01001110011: data <= 32'hb481b931;
    11'b01001110100: data <= 32'h3bb23912;
    11'b01001110101: data <= 32'h37b43e33;
    11'b01001110110: data <= 32'hbdd03b78;
    11'b01001110111: data <= 32'hc112b5c3;
    11'b01001111000: data <= 32'hbed8b72e;
    11'b01001111001: data <= 32'hb4be3992;
    11'b01001111010: data <= 32'h35f53c87;
    11'b01001111011: data <= 32'h393d2a9b;
    11'b01001111100: data <= 32'h3ce6ba26;
    11'b01001111101: data <= 32'h3def3560;
    11'b01001111110: data <= 32'h39894056;
    11'b01001111111: data <= 32'hb5244076;
    11'b01010000000: data <= 32'hb1d93459;
    11'b01010000001: data <= 32'h39f1be05;
    11'b01010000010: data <= 32'h3a63be95;
    11'b01010000011: data <= 32'hb2a8bc3b;
    11'b01010000100: data <= 32'hb7d1bbce;
    11'b01010000101: data <= 32'h3aa9bc12;
    11'b01010000110: data <= 32'h3fd0b5c1;
    11'b01010000111: data <= 32'h3ac43715;
    11'b01010001000: data <= 32'hbe8134e4;
    11'b01010001001: data <= 32'hc189b663;
    11'b01010001010: data <= 32'hbef1b5f9;
    11'b01010001011: data <= 32'hb5bb3534;
    11'b01010001100: data <= 32'hb16d345d;
    11'b01010001101: data <= 32'hb72bba02;
    11'b01010001110: data <= 32'h25dbbb7b;
    11'b01010001111: data <= 32'h3a573aae;
    11'b01010010000: data <= 32'h398f41b0;
    11'b01010010001: data <= 32'ha867414f;
    11'b01010010010: data <= 32'hb2503856;
    11'b01010010011: data <= 32'h342dbb95;
    11'b01010010100: data <= 32'h347fb8eb;
    11'b01010010101: data <= 32'hb1702c17;
    11'b01010010110: data <= 32'h33e9b62f;
    11'b01010010111: data <= 32'h3f4cbcd8;
    11'b01010011000: data <= 32'h4153bbb4;
    11'b01010011001: data <= 32'h3cd02ac2;
    11'b01010011010: data <= 32'hbce53655;
    11'b01010011011: data <= 32'hc006b121;
    11'b01010011100: data <= 32'hbaf0b878;
    11'b01010011101: data <= 32'h24f3b80a;
    11'b01010011110: data <= 32'hb8eabab7;
    11'b01010011111: data <= 32'hbd94be46;
    11'b01010100000: data <= 32'hba05bcfb;
    11'b01010100001: data <= 32'h388639b9;
    11'b01010100010: data <= 32'h3a204107;
    11'b01010100011: data <= 32'hb38f4058;
    11'b01010100100: data <= 32'hbbad36d4;
    11'b01010100101: data <= 32'hba2fb4ac;
    11'b01010100110: data <= 32'hb73a38bc;
    11'b01010100111: data <= 32'hb4e63c84;
    11'b01010101000: data <= 32'h378e289a;
    11'b01010101001: data <= 32'h3fdcbd1a;
    11'b01010101010: data <= 32'h4138bb61;
    11'b01010101011: data <= 32'h3d5c38a7;
    11'b01010101100: data <= 32'hb7763cd0;
    11'b01010101101: data <= 32'hb9c935c0;
    11'b01010101110: data <= 32'h3503b966;
    11'b01010101111: data <= 32'h37e5bc4b;
    11'b01010110000: data <= 32'hba85bd8f;
    11'b01010110001: data <= 32'hbeb4bf7b;
    11'b01010110010: data <= 32'hb8cdbe33;
    11'b01010110011: data <= 32'h3c3d9d6a;
    11'b01010110100: data <= 32'h3c2f3d65;
    11'b01010110101: data <= 32'hb8b03c5d;
    11'b01010110110: data <= 32'hbf362a9a;
    11'b01010110111: data <= 32'hbe6e303f;
    11'b01010111000: data <= 32'hbb9d3d12;
    11'b01010111001: data <= 32'hb9023db3;
    11'b01010111010: data <= 32'hac1eafcd;
    11'b01010111011: data <= 32'h3c60bd82;
    11'b01010111100: data <= 32'h3f39b76b;
    11'b01010111101: data <= 32'h3cc13e35;
    11'b01010111110: data <= 32'h32b34054;
    11'b01010111111: data <= 32'h34f83b15;
    11'b01011000000: data <= 32'h3c10b813;
    11'b01011000001: data <= 32'h38fdbae2;
    11'b01011000010: data <= 32'hbac3bb5a;
    11'b01011000011: data <= 32'hbd2abdb7;
    11'b01011000100: data <= 32'h34b2beae;
    11'b01011000101: data <= 32'h3feabb32;
    11'b01011000110: data <= 32'h3ddc2cd9;
    11'b01011000111: data <= 32'hb986302c;
    11'b01011001000: data <= 32'hc002b3a1;
    11'b01011001001: data <= 32'hbe4d32f6;
    11'b01011001010: data <= 32'hbad73c81;
    11'b01011001011: data <= 32'hbba73a7a;
    11'b01011001100: data <= 32'hbc4bbab2;
    11'b01011001101: data <= 32'hb428be77;
    11'b01011001110: data <= 32'h3a43ace2;
    11'b01011001111: data <= 32'h3b544054;
    11'b01011010000: data <= 32'h37ab4115;
    11'b01011010001: data <= 32'h38333c2d;
    11'b01011010010: data <= 32'h3a6faf62;
    11'b01011010011: data <= 32'h32f12de1;
    11'b01011010100: data <= 32'hbb193575;
    11'b01011010101: data <= 32'hb99db828;
    11'b01011010110: data <= 32'h3cc6be4d;
    11'b01011010111: data <= 32'h414dbdd8;
    11'b01011011000: data <= 32'h3f09b850;
    11'b01011011001: data <= 32'hb667ace6;
    11'b01011011010: data <= 32'hbd3ab088;
    11'b01011011011: data <= 32'hb8aa2eff;
    11'b01011011100: data <= 32'hb1ba3788;
    11'b01011011101: data <= 32'hbc74b1db;
    11'b01011011110: data <= 32'hbfd9be7f;
    11'b01011011111: data <= 32'hbd04bfa2;
    11'b01011100000: data <= 32'h3386b057;
    11'b01011100001: data <= 32'h3a793f7b;
    11'b01011100010: data <= 32'h35733fcf;
    11'b01011100011: data <= 32'ha949394b;
    11'b01011100100: data <= 32'had233447;
    11'b01011100101: data <= 32'hb7c53cee;
    11'b01011100110: data <= 32'hbc2d3e7a;
    11'b01011100111: data <= 32'hb77633bb;
    11'b01011101000: data <= 32'h3d67bdb4;
    11'b01011101001: data <= 32'h4106bddb;
    11'b01011101010: data <= 32'h3eacb317;
    11'b01011101011: data <= 32'h2f073863;
    11'b01011101100: data <= 32'had5a3563;
    11'b01011101101: data <= 32'h3a6e29a1;
    11'b01011101110: data <= 32'h3929abe5;
    11'b01011101111: data <= 32'hbc49b9d6;
    11'b01011110000: data <= 32'hc087bf76;
    11'b01011110001: data <= 32'hbd4cc010;
    11'b01011110010: data <= 32'h3819b924;
    11'b01011110011: data <= 32'h3c1a3a24;
    11'b01011110100: data <= 32'h2b813963;
    11'b01011110101: data <= 32'hba75ac3c;
    11'b01011110110: data <= 32'hbb1b36dc;
    11'b01011110111: data <= 32'hbb953fa6;
    11'b01011111000: data <= 32'hbcf3404b;
    11'b01011111001: data <= 32'hbaa3355f;
    11'b01011111010: data <= 32'h384abdbc;
    11'b01011111011: data <= 32'h3e1dbc4f;
    11'b01011111100: data <= 32'h3cb0391b;
    11'b01011111101: data <= 32'h38163dd5;
    11'b01011111110: data <= 32'h3b873abb;
    11'b01011111111: data <= 32'h3efd3046;
    11'b01100000000: data <= 32'h3c3f2604;
    11'b01100000001: data <= 32'hbbcdb4ed;
    11'b01100000010: data <= 32'hbfcbbd12;
    11'b01100000011: data <= 32'hb88ebf52;
    11'b01100000100: data <= 32'h3d68bd0c;
    11'b01100000101: data <= 32'h3db9b7cc;
    11'b01100000110: data <= 32'hacf4b84b;
    11'b01100000111: data <= 32'hbc5db969;
    11'b01100001000: data <= 32'hbb2d35a0;
    11'b01100001001: data <= 32'hb9ce3f55;
    11'b01100001010: data <= 32'hbd203ec9;
    11'b01100001011: data <= 32'hbe4eb449;
    11'b01100001100: data <= 32'hba56bea1;
    11'b01100001101: data <= 32'h3410b98a;
    11'b01100001110: data <= 32'h386c3d29;
    11'b01100001111: data <= 32'h38ae3f76;
    11'b01100010000: data <= 32'h3cd53b40;
    11'b01100010001: data <= 32'h3ee93496;
    11'b01100010010: data <= 32'h3a6e39e3;
    11'b01100010011: data <= 32'hbbea3b5f;
    11'b01100010100: data <= 32'hbd8caf3e;
    11'b01100010101: data <= 32'h355abd7d;
    11'b01100010110: data <= 32'h4016be65;
    11'b01100010111: data <= 32'h3ea4bc95;
    11'b01100011000: data <= 32'h253abbb3;
    11'b01100011001: data <= 32'hb8d3ba2b;
    11'b01100011010: data <= 32'h2bfd3238;
    11'b01100011011: data <= 32'h31cd3ce4;
    11'b01100011100: data <= 32'hbc4c39e1;
    11'b01100011101: data <= 32'hc071bc3f;
    11'b01100011110: data <= 32'hbf48bfa5;
    11'b01100011111: data <= 32'hb84cb8da;
    11'b01100100000: data <= 32'h32a23cb2;
    11'b01100100001: data <= 32'h35e13d3f;
    11'b01100100010: data <= 32'h3997350c;
    11'b01100100011: data <= 32'h3b483516;
    11'b01100100100: data <= 32'h2f513e80;
    11'b01100100101: data <= 32'hbc844074;
    11'b01100100110: data <= 32'hbc343b49;
    11'b01100100111: data <= 32'h3918bb87;
    11'b01100101000: data <= 32'h3fc8bdf3;
    11'b01100101001: data <= 32'h3d90bb1e;
    11'b01100101010: data <= 32'h3281b712;
    11'b01100101011: data <= 32'h35f2b55d;
    11'b01100101100: data <= 32'h3de22fbf;
    11'b01100101101: data <= 32'h3d1f390a;
    11'b01100101110: data <= 32'hb9b72cb8;
    11'b01100101111: data <= 32'hc0c0bd64;
    11'b01100110000: data <= 32'hbfd0bf90;
    11'b01100110001: data <= 32'hb66fba8e;
    11'b01100110010: data <= 32'h357934f5;
    11'b01100110011: data <= 32'h2cc12402;
    11'b01100110100: data <= 32'hae01b98a;
    11'b01100110101: data <= 32'h252e3057;
    11'b01100110110: data <= 32'hb65b4042;
    11'b01100110111: data <= 32'hbcdc41a2;
    11'b01100111000: data <= 32'hbca33cbc;
    11'b01100111001: data <= 32'h2a2aba92;
    11'b01100111010: data <= 32'h3b9ebc4c;
    11'b01100111011: data <= 32'h38f3a763;
    11'b01100111100: data <= 32'h33e2381f;
    11'b01100111101: data <= 32'h3cce32e1;
    11'b01100111110: data <= 32'h40f6307c;
    11'b01100111111: data <= 32'h3fa73807;
    11'b01101000000: data <= 32'hb7123493;
    11'b01101000001: data <= 32'hc005ba0d;
    11'b01101000010: data <= 32'hbcddbdb8;
    11'b01101000011: data <= 32'h3728bc50;
    11'b01101000100: data <= 32'h3a3eb9e5;
    11'b01101000101: data <= 32'haeb8bd0e;
    11'b01101000110: data <= 32'hb860be36;
    11'b01101000111: data <= 32'hb1b5b141;
    11'b01101001000: data <= 32'hb24b3fe9;
    11'b01101001001: data <= 32'hbc1e40cd;
    11'b01101001010: data <= 32'hbe3938de;
    11'b01101001011: data <= 32'hbc41bc38;
    11'b01101001100: data <= 32'hb649b94e;
    11'b01101001101: data <= 32'hb4793a08;
    11'b01101001110: data <= 32'h2acd3c5d;
    11'b01101001111: data <= 32'h3d7c3517;
    11'b01101010000: data <= 32'h41062e5b;
    11'b01101010001: data <= 32'h3ee73b1b;
    11'b01101010010: data <= 32'hb6f63d2f;
    11'b01101010011: data <= 32'hbdb63768;
    11'b01101010100: data <= 32'hb2dab966;
    11'b01101010101: data <= 32'h3d25bc71;
    11'b01101010110: data <= 32'h3c3dbd19;
    11'b01101010111: data <= 32'hb139bf08;
    11'b01101011000: data <= 32'hb5b3bf11;
    11'b01101011001: data <= 32'h3883b620;
    11'b01101011010: data <= 32'h3a193d60;
    11'b01101011011: data <= 32'hb82c3d7a;
    11'b01101011100: data <= 32'hbf7ab4e4;
    11'b01101011101: data <= 32'hbfcdbd77;
    11'b01101011110: data <= 32'hbd12b74e;
    11'b01101011111: data <= 32'hba5b3b39;
    11'b01101100000: data <= 32'hb45f39fe;
    11'b01101100001: data <= 32'h3aa2b4f1;
    11'b01101100010: data <= 32'h3e9db11d;
    11'b01101100011: data <= 32'h3b913dbe;
    11'b01101100100: data <= 32'hb90f40e3;
    11'b01101100101: data <= 32'hbc013e54;
    11'b01101100110: data <= 32'h3528a6c9;
    11'b01101100111: data <= 32'h3d93bab7;
    11'b01101101000: data <= 32'h3a32bbc6;
    11'b01101101001: data <= 32'hb402bce6;
    11'b01101101010: data <= 32'h346dbd1f;
    11'b01101101011: data <= 32'h3f37b688;
    11'b01101101100: data <= 32'h3fdb397a;
    11'b01101101101: data <= 32'h2e02380a;
    11'b01101101110: data <= 32'hbf44ba5d;
    11'b01101101111: data <= 32'hc009bd6b;
    11'b01101110000: data <= 32'hbc99b6d1;
    11'b01101110001: data <= 32'hb94135f5;
    11'b01101110010: data <= 32'hb856b5ee;
    11'b01101110011: data <= 32'ha291bdaf;
    11'b01101110100: data <= 32'h38b8b901;
    11'b01101110101: data <= 32'h33a93ec5;
    11'b01101110110: data <= 32'hba0341e8;
    11'b01101110111: data <= 32'hbb323f9a;
    11'b01101111000: data <= 32'h2af83098;
    11'b01101111001: data <= 32'h38aeb6a7;
    11'b01101111010: data <= 32'hae1fac62;
    11'b01101111011: data <= 32'hb80fb00d;
    11'b01101111100: data <= 32'h3aa2b866;
    11'b01101111101: data <= 32'h4171b564;
    11'b01101111110: data <= 32'h4156361e;
    11'b01101111111: data <= 32'h378b369a;
    11'b01110000000: data <= 32'hbd98b65d;
    11'b01110000001: data <= 32'hbcf5ba7b;
    11'b01110000010: data <= 32'hb218b616;
    11'b01110000011: data <= 32'hac19b603;
    11'b01110000100: data <= 32'hb946be31;
    11'b01110000101: data <= 32'hb8dfc0c2;
    11'b01110000110: data <= 32'h2ed6bc55;
    11'b01110000111: data <= 32'h33813dc4;
    11'b01110001000: data <= 32'hb80d40fb;
    11'b01110001001: data <= 32'hbbfe3cff;
    11'b01110001010: data <= 32'hb9f5b2b7;
    11'b01110001011: data <= 32'hb92dac03;
    11'b01110001100: data <= 32'hbc753aa6;
    11'b01110001101: data <= 32'hbb4339b0;
    11'b01110001110: data <= 32'h3adeb376;
    11'b01110001111: data <= 32'h4168b684;
    11'b01110010000: data <= 32'h40e237d8;
    11'b01110010001: data <= 32'h366b3c6a;
    11'b01110010010: data <= 32'hbae23991;
    11'b01110010011: data <= 32'hb0722cec;
    11'b01110010100: data <= 32'h3b19b140;
    11'b01110010101: data <= 32'h36ecb9dd;
    11'b01110010110: data <= 32'hb9bebff6;
    11'b01110010111: data <= 32'hb95bc130;
    11'b01110011000: data <= 32'h383dbd1a;
    11'b01110011001: data <= 32'h3c353aa3;
    11'b01110011010: data <= 32'h303e3d7f;
    11'b01110011011: data <= 32'hbc242fa5;
    11'b01110011100: data <= 32'hbdabb9e1;
    11'b01110011101: data <= 32'hbde02fbc;
    11'b01110011110: data <= 32'hbeb03cd1;
    11'b01110011111: data <= 32'hbd0e397b;
    11'b01110100000: data <= 32'h34edb99b;
    11'b01110100001: data <= 32'h3f13ba49;
    11'b01110100010: data <= 32'h3de739f4;
    11'b01110100011: data <= 32'h18784004;
    11'b01110100100: data <= 32'hb7913f08;
    11'b01110100101: data <= 32'h38c73a75;
    11'b01110100110: data <= 32'h3d39324c;
    11'b01110100111: data <= 32'h3533b62f;
    11'b01110101000: data <= 32'hbb3cbd93;
    11'b01110101001: data <= 32'hb54dbfd3;
    11'b01110101010: data <= 32'h3e07bc7d;
    11'b01110101011: data <= 32'h406132f7;
    11'b01110101100: data <= 32'h3ae3354c;
    11'b01110101101: data <= 32'hbab2b966;
    11'b01110101110: data <= 32'hbd9dbb5d;
    11'b01110101111: data <= 32'hbd303332;
    11'b01110110000: data <= 32'hbdb63bb2;
    11'b01110110001: data <= 32'hbd90b108;
    11'b01110110010: data <= 32'hb7d1bef4;
    11'b01110110011: data <= 32'h3861bd8a;
    11'b01110110100: data <= 32'h37913a7a;
    11'b01110110101: data <= 32'hb54f40cd;
    11'b01110110110: data <= 32'hb5324010;
    11'b01110110111: data <= 32'h38db3b5a;
    11'b01110111000: data <= 32'h3a4c3834;
    11'b01110111001: data <= 32'hb74d37bb;
    11'b01110111010: data <= 32'hbd38b103;
    11'b01110111011: data <= 32'h9e37bb93;
    11'b01110111100: data <= 32'h408dba98;
    11'b01110111101: data <= 32'h41b7ae98;
    11'b01110111110: data <= 32'h3ceba679;
    11'b01110111111: data <= 32'hb755b8a5;
    11'b01111000000: data <= 32'hb917b7c5;
    11'b01111000001: data <= 32'hb2f3369f;
    11'b01111000010: data <= 32'hb8a43778;
    11'b01111000011: data <= 32'hbd20bca5;
    11'b01111000100: data <= 32'hbc52c156;
    11'b01111000101: data <= 32'hb1e2bf86;
    11'b01111000110: data <= 32'h30de3857;
    11'b01111000111: data <= 32'hb32b3fb3;
    11'b01111001000: data <= 32'hb4ae3d1b;
    11'b01111001001: data <= 32'h2cfc3587;
    11'b01111001010: data <= 32'hb3f63956;
    11'b01111001011: data <= 32'hbdcd3d75;
    11'b01111001100: data <= 32'hbf243b4d;
    11'b01111001101: data <= 32'ha9eab4e3;
    11'b01111001110: data <= 32'h4070b9d2;
    11'b01111001111: data <= 32'h4117aed2;
    11'b01111010000: data <= 32'h3bd8362e;
    11'b01111010001: data <= 32'haeb034ae;
    11'b01111010010: data <= 32'h371435fc;
    11'b01111010011: data <= 32'h3c4e39f4;
    11'b01111010100: data <= 32'h33c6334a;
    11'b01111010101: data <= 32'hbc96be2b;
    11'b01111010110: data <= 32'hbce8c1a3;
    11'b01111010111: data <= 32'ha978bfc4;
    11'b01111011000: data <= 32'h39cb2cff;
    11'b01111011001: data <= 32'h35fd3a9b;
    11'b01111011010: data <= 32'hb221aae5;
    11'b01111011011: data <= 32'hb6ebb802;
    11'b01111011100: data <= 32'hbbe5391b;
    11'b01111011101: data <= 32'hbfe03f32;
    11'b01111011110: data <= 32'hc0213caa;
    11'b01111011111: data <= 32'hb7e3b806;
    11'b01111100000: data <= 32'h3d2ebc2b;
    11'b01111100001: data <= 32'h3d951842;
    11'b01111100010: data <= 32'h345f3c5f;
    11'b01111100011: data <= 32'h2bda3cfd;
    11'b01111100100: data <= 32'h3ce13c58;
    11'b01111100101: data <= 32'h3f163c56;
    11'b01111100110: data <= 32'h36da3828;
    11'b01111100111: data <= 32'hbcf6bb90;
    11'b01111101000: data <= 32'hbc1fc00b;
    11'b01111101001: data <= 32'h39b1be04;
    11'b01111101010: data <= 32'h3eecb504;
    11'b01111101011: data <= 32'h3c64b3e0;
    11'b01111101100: data <= 32'h28b7bc7d;
    11'b01111101101: data <= 32'hb6c5bc01;
    11'b01111101110: data <= 32'hba6c38f5;
    11'b01111101111: data <= 32'hbe603ec0;
    11'b01111110000: data <= 32'hbfc53886;
    11'b01111110001: data <= 32'hbc54bd89;
    11'b01111110010: data <= 32'h2aecbe8f;
    11'b01111110011: data <= 32'h2fea9c93;
    11'b01111110100: data <= 32'hb64e3dc4;
    11'b01111110101: data <= 32'h2b4e3dfc;
    11'b01111110110: data <= 32'h3d643c67;
    11'b01111110111: data <= 32'h3e0a3cda;
    11'b01111111000: data <= 32'hb16c3cd3;
    11'b01111111001: data <= 32'hbe8934e3;
    11'b01111111010: data <= 32'hba73ba05;
    11'b01111111011: data <= 32'h3d94bae5;
    11'b01111111100: data <= 32'h40b8b747;
    11'b01111111101: data <= 32'h3d9bb9a5;
    11'b01111111110: data <= 32'h3453bd34;
    11'b01111111111: data <= 32'h3246ba40;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    