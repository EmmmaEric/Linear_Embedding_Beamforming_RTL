
module memory_rom_31(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hb92bbdc9;
    11'b00000000001: data <= 32'hb67fba45;
    11'b00000000010: data <= 32'h358e3b0b;
    11'b00000000011: data <= 32'haf0b3f7c;
    11'b00000000100: data <= 32'hbe163a8f;
    11'b00000000101: data <= 32'hc046bbf7;
    11'b00000000110: data <= 32'hbd97bcbf;
    11'b00000000111: data <= 32'hb6e23590;
    11'b00000001000: data <= 32'h2c253d69;
    11'b00000001001: data <= 32'h3953394b;
    11'b00000001010: data <= 32'h3e28b14e;
    11'b00000001011: data <= 32'h3e393862;
    11'b00000001100: data <= 32'h31683fa8;
    11'b00000001101: data <= 32'hbc643f6d;
    11'b00000001110: data <= 32'hb85732ee;
    11'b00000001111: data <= 32'h3c58bce5;
    11'b00000010000: data <= 32'h3e25bdcf;
    11'b00000010001: data <= 32'h368ebce8;
    11'b00000010010: data <= 32'hb4a3bcc2;
    11'b00000010011: data <= 32'h3918ba19;
    11'b00000010100: data <= 32'h3e763544;
    11'b00000010101: data <= 32'h39713b2f;
    11'b00000010110: data <= 32'hbdfaa332;
    11'b00000010111: data <= 32'hc118bd22;
    11'b00000011000: data <= 32'hbef4bc7a;
    11'b00000011001: data <= 32'hb8713150;
    11'b00000011010: data <= 32'hb1093899;
    11'b00000011011: data <= 32'h9ba4b622;
    11'b00000011100: data <= 32'h37eeba1a;
    11'b00000011101: data <= 32'h391c3a58;
    11'b00000011110: data <= 32'hb1884170;
    11'b00000011111: data <= 32'hbb88413d;
    11'b00000100000: data <= 32'hb6e8392b;
    11'b00000100001: data <= 32'h39aebb17;
    11'b00000100010: data <= 32'h3abcba8c;
    11'b00000100011: data <= 32'h2a8cb47d;
    11'b00000100100: data <= 32'h3179b601;
    11'b00000100101: data <= 32'h3eeeb858;
    11'b00000100110: data <= 32'h4164a922;
    11'b00000100111: data <= 32'h3d2e3700;
    11'b00000101000: data <= 32'hbcd0ac81;
    11'b00000101001: data <= 32'hc047bbb5;
    11'b00000101010: data <= 32'hbc41bbd5;
    11'b00000101011: data <= 32'h2545b657;
    11'b00000101100: data <= 32'hb12eb8ff;
    11'b00000101101: data <= 32'hb927be62;
    11'b00000101110: data <= 32'hb4f3bdad;
    11'b00000101111: data <= 32'h32de3976;
    11'b00000110000: data <= 32'hb0774162;
    11'b00000110001: data <= 32'hbb5940b9;
    11'b00000110010: data <= 32'hbba13636;
    11'b00000110011: data <= 32'hb640b93f;
    11'b00000110100: data <= 32'hb4ac29df;
    11'b00000110101: data <= 32'hb7f43a4e;
    11'b00000110110: data <= 32'h352034b9;
    11'b00000110111: data <= 32'h4049b725;
    11'b00000111000: data <= 32'h41d5aee3;
    11'b00000111001: data <= 32'h3d7e3a1c;
    11'b00000111010: data <= 32'hba923a2a;
    11'b00000111011: data <= 32'hbccbac93;
    11'b00000111100: data <= 32'h2eb4b93b;
    11'b00000111101: data <= 32'h3a46ba9f;
    11'b00000111110: data <= 32'hadf0bdb3;
    11'b00000111111: data <= 32'hbb5dc078;
    11'b00001000000: data <= 32'hb526bf15;
    11'b00001000001: data <= 32'h398f3432;
    11'b00001000010: data <= 32'h37233f76;
    11'b00001000011: data <= 32'hbabc3d3c;
    11'b00001000100: data <= 32'hbe80b4c9;
    11'b00001000101: data <= 32'hbddab8ac;
    11'b00001000110: data <= 32'hbcc538ff;
    11'b00001000111: data <= 32'hbbd83ce4;
    11'b00001001000: data <= 32'h9caf32e3;
    11'b00001001001: data <= 32'h3e63ba0a;
    11'b00001001010: data <= 32'h4058a531;
    11'b00001001011: data <= 32'h3b563e3a;
    11'b00001001100: data <= 32'hb8613fd6;
    11'b00001001101: data <= 32'hb53a3b3d;
    11'b00001001110: data <= 32'h3b7eb2f6;
    11'b00001001111: data <= 32'h3c47b9e4;
    11'b00001010000: data <= 32'hb2c7bd15;
    11'b00001010001: data <= 32'hba9bbfa4;
    11'b00001010010: data <= 32'h3676be89;
    11'b00001010011: data <= 32'h3f49b2f7;
    11'b00001010100: data <= 32'h3d5a3a5e;
    11'b00001010101: data <= 32'hb8c532f7;
    11'b00001010110: data <= 32'hbf7dba9e;
    11'b00001010111: data <= 32'hbefcb849;
    11'b00001011000: data <= 32'hbd293978;
    11'b00001011001: data <= 32'hbc8e3a1c;
    11'b00001011010: data <= 32'hb8ffb962;
    11'b00001011011: data <= 32'h378dbdd1;
    11'b00001011100: data <= 32'h3c15a62d;
    11'b00001011101: data <= 32'h35574052;
    11'b00001011110: data <= 32'hb6f34151;
    11'b00001011111: data <= 32'h16393d62;
    11'b00001100000: data <= 32'h3b0b2f4a;
    11'b00001100001: data <= 32'h3863af95;
    11'b00001100010: data <= 32'hb953b40c;
    11'b00001100011: data <= 32'hb90dbb1c;
    11'b00001100100: data <= 32'h3d14bcb9;
    11'b00001100101: data <= 32'h41aab830;
    11'b00001100110: data <= 32'h4000308c;
    11'b00001100111: data <= 32'hb40ab10b;
    11'b00001101000: data <= 32'hbdc4b99e;
    11'b00001101001: data <= 32'hbc07b510;
    11'b00001101010: data <= 32'hb8553654;
    11'b00001101011: data <= 32'hbb76b1d6;
    11'b00001101100: data <= 32'hbcc5bf3e;
    11'b00001101101: data <= 32'hb806c062;
    11'b00001101110: data <= 32'h347fb3bf;
    11'b00001101111: data <= 32'h30c34024;
    11'b00001110000: data <= 32'hb5bd40ae;
    11'b00001110001: data <= 32'hb3e83ba4;
    11'b00001110010: data <= 32'h2aa13169;
    11'b00001110011: data <= 32'hb8003967;
    11'b00001110100: data <= 32'hbd463bbb;
    11'b00001110101: data <= 32'hb91b2da8;
    11'b00001110110: data <= 32'h3e54bac6;
    11'b00001110111: data <= 32'h41ffb8e9;
    11'b00001111000: data <= 32'h3ff4328b;
    11'b00001111001: data <= 32'h92a5364d;
    11'b00001111010: data <= 32'hb8752da1;
    11'b00001111011: data <= 32'h34bf300f;
    11'b00001111100: data <= 32'h381d3128;
    11'b00001111101: data <= 32'hb8eabad4;
    11'b00001111110: data <= 32'hbddac0ce;
    11'b00001111111: data <= 32'hba1fc100;
    11'b00010000000: data <= 32'h374eb8aa;
    11'b00010000001: data <= 32'h38df3d1f;
    11'b00010000010: data <= 32'hb1383ca9;
    11'b00010000011: data <= 32'hb9879cb7;
    11'b00010000100: data <= 32'hbae5a0ca;
    11'b00010000101: data <= 32'hbd743ce9;
    11'b00010000110: data <= 32'hbf3b3e8a;
    11'b00010000111: data <= 32'hbb843533;
    11'b00010001000: data <= 32'h3c31bc01;
    11'b00010001001: data <= 32'h404bb910;
    11'b00010001010: data <= 32'h3d2739ff;
    11'b00010001011: data <= 32'h282a3d94;
    11'b00010001100: data <= 32'h34633c1d;
    11'b00010001101: data <= 32'h3d6638e8;
    11'b00010001110: data <= 32'h3c803491;
    11'b00010001111: data <= 32'hb868b97b;
    11'b00010010000: data <= 32'hbdd1bff7;
    11'b00010010001: data <= 32'hb4bdc04f;
    11'b00010010010: data <= 32'h3d7abac1;
    11'b00010010011: data <= 32'h3dd63419;
    11'b00010010100: data <= 32'h3159b058;
    11'b00010010101: data <= 32'hbad1baec;
    11'b00010010110: data <= 32'hbc69b173;
    11'b00010010111: data <= 32'hbd933d66;
    11'b00010011000: data <= 32'hbf3a3dbe;
    11'b00010011001: data <= 32'hbd7fb536;
    11'b00010011010: data <= 32'ha83abe96;
    11'b00010011011: data <= 32'h3a65b9f2;
    11'b00010011100: data <= 32'h35ef3ce4;
    11'b00010011101: data <= 32'had82400c;
    11'b00010011110: data <= 32'h39253db1;
    11'b00010011111: data <= 32'h3e383ab6;
    11'b00010100000: data <= 32'h3aef3a19;
    11'b00010100001: data <= 32'hbb6f34bd;
    11'b00010100010: data <= 32'hbd81ba53;
    11'b00010100011: data <= 32'h3675bd83;
    11'b00010100100: data <= 32'h4092bb3a;
    11'b00010100101: data <= 32'h402fb6af;
    11'b00010100110: data <= 32'h3756ba31;
    11'b00010100111: data <= 32'hb817bc1e;
    11'b00010101000: data <= 32'hb631aad1;
    11'b00010101001: data <= 32'hb7ce3cb6;
    11'b00010101010: data <= 32'hbd303976;
    11'b00010101011: data <= 32'hbec5bd62;
    11'b00010101100: data <= 32'hbc0bc0ba;
    11'b00010101101: data <= 32'hb276bba9;
    11'b00010101110: data <= 32'hb0263cb0;
    11'b00010101111: data <= 32'hb0a33edc;
    11'b00010110000: data <= 32'h38073b31;
    11'b00010110001: data <= 32'h3b893900;
    11'b00010110010: data <= 32'ha9193d46;
    11'b00010110011: data <= 32'hbe473e08;
    11'b00010110100: data <= 32'hbdaf3719;
    11'b00010110101: data <= 32'h39aab9a5;
    11'b00010110110: data <= 32'h40e3ba98;
    11'b00010110111: data <= 32'h3fe5b735;
    11'b00010111000: data <= 32'h37c2b753;
    11'b00010111001: data <= 32'h311bb694;
    11'b00010111010: data <= 32'h3b3e35fb;
    11'b00010111011: data <= 32'h3a893c0f;
    11'b00010111100: data <= 32'hb9062bed;
    11'b00010111101: data <= 32'hbf0dbfac;
    11'b00010111110: data <= 32'hbd67c131;
    11'b00010111111: data <= 32'hb475bc7d;
    11'b00011000000: data <= 32'h2fdf387f;
    11'b00011000001: data <= 32'h24d73866;
    11'b00011000010: data <= 32'h30eab4bd;
    11'b00011000011: data <= 32'h2f8e2e19;
    11'b00011000100: data <= 32'hbaf33e99;
    11'b00011000101: data <= 32'hc0064079;
    11'b00011000110: data <= 32'hbe643b92;
    11'b00011000111: data <= 32'h3518b8ed;
    11'b00011001000: data <= 32'h3e69ba49;
    11'b00011001001: data <= 32'h3c3aa1ba;
    11'b00011001010: data <= 32'h31a936ae;
    11'b00011001011: data <= 32'h3a1737a2;
    11'b00011001100: data <= 32'h40043ab8;
    11'b00011001101: data <= 32'h3ed23c45;
    11'b00011001110: data <= 32'hb48a3007;
    11'b00011001111: data <= 32'hbea8be0e;
    11'b00011010000: data <= 32'hbbebc020;
    11'b00011010001: data <= 32'h37a2bc41;
    11'b00011010010: data <= 32'h3b2cb373;
    11'b00011010011: data <= 32'h3585ba58;
    11'b00011010100: data <= 32'ha785bdc6;
    11'b00011010101: data <= 32'hb202b60e;
    11'b00011010110: data <= 32'hbb443e99;
    11'b00011010111: data <= 32'hbf6c4049;
    11'b00011011000: data <= 32'hbefe37b4;
    11'b00011011001: data <= 32'hb859bc9c;
    11'b00011011010: data <= 32'h32fdbb28;
    11'b00011011011: data <= 32'hb0de371c;
    11'b00011011100: data <= 32'hb47d3c4a;
    11'b00011011101: data <= 32'h3bd33b08;
    11'b00011011110: data <= 32'h40a03b98;
    11'b00011011111: data <= 32'h3ea43d38;
    11'b00011100000: data <= 32'hb8273b3e;
    11'b00011100001: data <= 32'hbe4fb48d;
    11'b00011100010: data <= 32'hb562bbfb;
    11'b00011100011: data <= 32'h3d86ba23;
    11'b00011100100: data <= 32'h3e21b9d8;
    11'b00011100101: data <= 32'h3875be1c;
    11'b00011100110: data <= 32'h2fc8bf67;
    11'b00011100111: data <= 32'h359fb71d;
    11'b00011101000: data <= 32'h24af3dcf;
    11'b00011101001: data <= 32'hbc4d3dd3;
    11'b00011101010: data <= 32'hbed3b7e0;
    11'b00011101011: data <= 32'hbd4fbf75;
    11'b00011101100: data <= 32'hbb03bc3f;
    11'b00011101101: data <= 32'hbb663843;
    11'b00011101110: data <= 32'hb8873b49;
    11'b00011101111: data <= 32'h3a523582;
    11'b00011110000: data <= 32'h3f2037dc;
    11'b00011110001: data <= 32'h3aac3e0d;
    11'b00011110010: data <= 32'hbc8c3fa7;
    11'b00011110011: data <= 32'hbe653c28;
    11'b00011110100: data <= 32'h2bf8a759;
    11'b00011110101: data <= 32'h3ea2b6af;
    11'b00011110110: data <= 32'h3da7b980;
    11'b00011110111: data <= 32'h35fbbd3a;
    11'b00011111000: data <= 32'h3786bd66;
    11'b00011111001: data <= 32'h3dc3abf7;
    11'b00011111010: data <= 32'h3da03d1f;
    11'b00011111011: data <= 32'hae063a3f;
    11'b00011111100: data <= 32'hbde0bca0;
    11'b00011111101: data <= 32'hbe41c036;
    11'b00011111110: data <= 32'hbc3bbc38;
    11'b00011111111: data <= 32'hbaa632c1;
    11'b00100000000: data <= 32'hb7b1abc0;
    11'b00100000001: data <= 32'h36febb6a;
    11'b00100000010: data <= 32'h3b81b5ae;
    11'b00100000011: data <= 32'hab953e0a;
    11'b00100000100: data <= 32'hbe664107;
    11'b00100000101: data <= 32'hbe943e9d;
    11'b00100000110: data <= 32'hacfb3435;
    11'b00100000111: data <= 32'h3bffb420;
    11'b00100001000: data <= 32'h36e1b3a5;
    11'b00100001001: data <= 32'hb3ceb714;
    11'b00100001010: data <= 32'h39cdb6da;
    11'b00100001011: data <= 32'h40cb36d6;
    11'b00100001100: data <= 32'h40d33cf7;
    11'b00100001101: data <= 32'h37de3915;
    11'b00100001110: data <= 32'hbccebb61;
    11'b00100001111: data <= 32'hbcb5be15;
    11'b00100010000: data <= 32'hb56fb9a2;
    11'b00100010001: data <= 32'habb6b393;
    11'b00100010010: data <= 32'hb060bcfc;
    11'b00100010011: data <= 32'h323fc065;
    11'b00100010100: data <= 32'h376dbc6c;
    11'b00100010101: data <= 32'hb41a3d2e;
    11'b00100010110: data <= 32'hbda740bf;
    11'b00100010111: data <= 32'hbe1e3cfe;
    11'b00100011000: data <= 32'hb8d1b35e;
    11'b00100011001: data <= 32'hb320b5df;
    11'b00100011010: data <= 32'hbb413409;
    11'b00100011011: data <= 32'hbc073575;
    11'b00100011100: data <= 32'h397f2f78;
    11'b00100011101: data <= 32'h4146383e;
    11'b00100011110: data <= 32'h40e63d00;
    11'b00100011111: data <= 32'h35863c63;
    11'b00100100000: data <= 32'hbc583081;
    11'b00100100001: data <= 32'hb7ffb54a;
    11'b00100100010: data <= 32'h3942ad41;
    11'b00100100011: data <= 32'h3997b724;
    11'b00100100100: data <= 32'h2dbcbf9a;
    11'b00100100101: data <= 32'h3121c16b;
    11'b00100100110: data <= 32'h39b1bd3c;
    11'b00100100111: data <= 32'h38013c21;
    11'b00100101000: data <= 32'hb8263eaa;
    11'b00100101001: data <= 32'hbc9f32dc;
    11'b00100101010: data <= 32'hbc4bbc2a;
    11'b00100101011: data <= 32'hbce5b87c;
    11'b00100101100: data <= 32'hbf3937ca;
    11'b00100101101: data <= 32'hbdeb3707;
    11'b00100101110: data <= 32'h3648b3f1;
    11'b00100101111: data <= 32'h4029a585;
    11'b00100110000: data <= 32'h3e5f3c8a;
    11'b00100110001: data <= 32'hb57f3f1d;
    11'b00100110010: data <= 32'hbc8c3d6f;
    11'b00100110011: data <= 32'h21c63a45;
    11'b00100110100: data <= 32'h3ca73807;
    11'b00100110101: data <= 32'h39fdb40a;
    11'b00100110110: data <= 32'hb132be99;
    11'b00100110111: data <= 32'h329ec06c;
    11'b00100111000: data <= 32'h3de4bb23;
    11'b00100111001: data <= 32'h3f173b14;
    11'b00100111010: data <= 32'h38f53b3c;
    11'b00100111011: data <= 32'hb91eb931;
    11'b00100111100: data <= 32'hbc75bdcc;
    11'b00100111101: data <= 32'hbd79b819;
    11'b00100111110: data <= 32'hbf0036ff;
    11'b00100111111: data <= 32'hbd9fb2c5;
    11'b00101000000: data <= 32'h29f6bd93;
    11'b00101000001: data <= 32'h3cb0bc1c;
    11'b00101000010: data <= 32'h383a3a96;
    11'b00101000011: data <= 32'hbbbf404b;
    11'b00101000100: data <= 32'hbcab3fb7;
    11'b00101000101: data <= 32'h2f183c9a;
    11'b00101000110: data <= 32'h3a7d39d5;
    11'b00101000111: data <= 32'hae7732ef;
    11'b00101001000: data <= 32'hbb78b9de;
    11'b00101001001: data <= 32'h305fbc98;
    11'b00101001010: data <= 32'h4055b400;
    11'b00101001011: data <= 32'h41743ad3;
    11'b00101001100: data <= 32'h3d42386c;
    11'b00101001101: data <= 32'hb3ffb9aa;
    11'b00101001110: data <= 32'hb95fbc08;
    11'b00101001111: data <= 32'hb8dda5c4;
    11'b00101010000: data <= 32'hbb003516;
    11'b00101010001: data <= 32'hbb6fbc78;
    11'b00101010010: data <= 32'hb184c137;
    11'b00101010011: data <= 32'h3831bfab;
    11'b00101010100: data <= 32'h2ae036e5;
    11'b00101010101: data <= 32'hbb833fa3;
    11'b00101010110: data <= 32'hbb7d3df1;
    11'b00101010111: data <= 32'hade738bd;
    11'b00101011000: data <= 32'hafac3829;
    11'b00101011001: data <= 32'hbd7f3972;
    11'b00101011010: data <= 32'hbf703236;
    11'b00101011011: data <= 32'hb00bb584;
    11'b00101011100: data <= 32'h408b261b;
    11'b00101011101: data <= 32'h41753a34;
    11'b00101011110: data <= 32'h3c9539ab;
    11'b00101011111: data <= 32'hb2172b50;
    11'b00101100000: data <= 32'ha2842f06;
    11'b00101100001: data <= 32'h38123a3a;
    11'b00101100010: data <= 32'h2fb835f7;
    11'b00101100011: data <= 32'hb82fbe6a;
    11'b00101100100: data <= 32'hb42ec22d;
    11'b00101100101: data <= 32'h37d2c048;
    11'b00101100110: data <= 32'h38123197;
    11'b00101100111: data <= 32'hb0323ccd;
    11'b00101101000: data <= 32'hb6113599;
    11'b00101101001: data <= 32'hb44fb6dc;
    11'b00101101010: data <= 32'hbb6630b3;
    11'b00101101011: data <= 32'hc0803b87;
    11'b00101101100: data <= 32'hc0cc3862;
    11'b00101101101: data <= 32'hb781b684;
    11'b00101101110: data <= 32'h3ec4b6bc;
    11'b00101101111: data <= 32'h3f2537c8;
    11'b00101110000: data <= 32'h346f3c4f;
    11'b00101110001: data <= 32'hb6903c38;
    11'b00101110010: data <= 32'h38093cd3;
    11'b00101110011: data <= 32'h3cfa3de7;
    11'b00101110100: data <= 32'h3785395d;
    11'b00101110101: data <= 32'hb92abd32;
    11'b00101110110: data <= 32'hb5e5c10a;
    11'b00101110111: data <= 32'h3b77be54;
    11'b00101111000: data <= 32'h3e293192;
    11'b00101111001: data <= 32'h3be93711;
    11'b00101111010: data <= 32'h3493b9c3;
    11'b00101111011: data <= 32'hb0ddbc86;
    11'b00101111100: data <= 32'hbbe829b1;
    11'b00101111101: data <= 32'hc0493c12;
    11'b00101111110: data <= 32'hc07432b1;
    11'b00101111111: data <= 32'hb999bd2f;
    11'b00110000000: data <= 32'h3a4abd9a;
    11'b00110000001: data <= 32'h384791d2;
    11'b00110000010: data <= 32'hb9113cf5;
    11'b00110000011: data <= 32'hb8df3e0f;
    11'b00110000100: data <= 32'h39a03e2a;
    11'b00110000101: data <= 32'h3cc63ea0;
    11'b00110000110: data <= 32'haf033c45;
    11'b00110000111: data <= 32'hbd81b621;
    11'b00110001000: data <= 32'hb902bd2c;
    11'b00110001001: data <= 32'h3d89b957;
    11'b00110001010: data <= 32'h40b7352e;
    11'b00110001011: data <= 32'h3eae2451;
    11'b00110001100: data <= 32'h397dbc46;
    11'b00110001101: data <= 32'h3454bbc9;
    11'b00110001110: data <= 32'hb2e33796;
    11'b00110001111: data <= 32'hbc813c58;
    11'b00110010000: data <= 32'hbe02b6dd;
    11'b00110010001: data <= 32'hb9dfc0b4;
    11'b00110010010: data <= 32'h2d97c094;
    11'b00110010011: data <= 32'hb2f4b74a;
    11'b00110010100: data <= 32'hbb353bbf;
    11'b00110010101: data <= 32'hb7673c2c;
    11'b00110010110: data <= 32'h396f3af0;
    11'b00110010111: data <= 32'h385f3cee;
    11'b00110011000: data <= 32'hbcd23d6c;
    11'b00110011001: data <= 32'hc09f38a1;
    11'b00110011010: data <= 32'hbbf8b32f;
    11'b00110011011: data <= 32'h3d9cad6a;
    11'b00110011100: data <= 32'h409f35c2;
    11'b00110011101: data <= 32'h3da520c8;
    11'b00110011110: data <= 32'h389eb8c9;
    11'b00110011111: data <= 32'h3a38aaa5;
    11'b00110100000: data <= 32'h3b693d24;
    11'b00110100001: data <= 32'h2f7d3d23;
    11'b00110100010: data <= 32'hba3eba43;
    11'b00110100011: data <= 32'hb971c189;
    11'b00110100100: data <= 32'hadb3c0e8;
    11'b00110100101: data <= 32'hac0fb8c3;
    11'b00110100110: data <= 32'hb5043603;
    11'b00110100111: data <= 32'h2e45af71;
    11'b00110101000: data <= 32'h395eb61e;
    11'b00110101001: data <= 32'had953862;
    11'b00110101010: data <= 32'hc0003dcf;
    11'b00110101011: data <= 32'hc1a33c33;
    11'b00110101100: data <= 32'hbd1c2475;
    11'b00110101101: data <= 32'h3b2db486;
    11'b00110101110: data <= 32'h3d5e2d71;
    11'b00110101111: data <= 32'h35643242;
    11'b00110110000: data <= 32'h2bb9323a;
    11'b00110110001: data <= 32'h3c7a3b99;
    11'b00110110010: data <= 32'h3f093feb;
    11'b00110110011: data <= 32'h3a293e4e;
    11'b00110110100: data <= 32'hb909b815;
    11'b00110110101: data <= 32'hb9f8c055;
    11'b00110110110: data <= 32'h316fbedc;
    11'b00110110111: data <= 32'h39e0b52f;
    11'b00110111000: data <= 32'h398cb2ab;
    11'b00110111001: data <= 32'h3a41bd13;
    11'b00110111010: data <= 32'h3ab0bd8b;
    11'b00110111011: data <= 32'hb06930c4;
    11'b00110111100: data <= 32'hbf713dd4;
    11'b00110111101: data <= 32'hc1003b1d;
    11'b00110111110: data <= 32'hbd17b8ee;
    11'b00110111111: data <= 32'h30f2bc81;
    11'b00111000000: data <= 32'h24b5b6e8;
    11'b00111000001: data <= 32'hbaf73439;
    11'b00111000010: data <= 32'hb73f38ca;
    11'b00111000011: data <= 32'h3cde3cfe;
    11'b00111000100: data <= 32'h3f7f401b;
    11'b00111000101: data <= 32'h376c3f23;
    11'b00111000110: data <= 32'hbcc93439;
    11'b00111000111: data <= 32'hbc20bafe;
    11'b00111001000: data <= 32'h37e2b818;
    11'b00111001001: data <= 32'h3dd330d1;
    11'b00111001010: data <= 32'h3d55b80f;
    11'b00111001011: data <= 32'h3c77bf16;
    11'b00111001100: data <= 32'h3c7fbe11;
    11'b00111001101: data <= 32'h382b3629;
    11'b00111001110: data <= 32'hba473e2a;
    11'b00111001111: data <= 32'hbe05366d;
    11'b00111010000: data <= 32'hbbd8be28;
    11'b00111010001: data <= 32'hb669bfdd;
    11'b00111010010: data <= 32'hbb05bade;
    11'b00111010011: data <= 32'hbdc62c67;
    11'b00111010100: data <= 32'hb844329b;
    11'b00111010101: data <= 32'h3cc23830;
    11'b00111010110: data <= 32'h3d8f3d8d;
    11'b00111010111: data <= 32'hb7833f0a;
    11'b00111011000: data <= 32'hc0243c4a;
    11'b00111011001: data <= 32'hbd9d3541;
    11'b00111011010: data <= 32'h38453644;
    11'b00111011011: data <= 32'h3dd0372b;
    11'b00111011100: data <= 32'h3c20b7cc;
    11'b00111011101: data <= 32'h3a6abde2;
    11'b00111011110: data <= 32'h3d63ba4d;
    11'b00111011111: data <= 32'h3e0a3c79;
    11'b00111100000: data <= 32'h38a93f0c;
    11'b00111100001: data <= 32'hb7412c9a;
    11'b00111100010: data <= 32'hb912bfdb;
    11'b00111100011: data <= 32'hb82cc030;
    11'b00111100100: data <= 32'hbb30baad;
    11'b00111100101: data <= 32'hbc50b477;
    11'b00111100110: data <= 32'hacbdba7b;
    11'b00111100111: data <= 32'h3cdbbab8;
    11'b00111101000: data <= 32'h3a8d35f8;
    11'b00111101001: data <= 32'hbcf93e28;
    11'b00111101010: data <= 32'hc11a3dd8;
    11'b00111101011: data <= 32'hbe4239f8;
    11'b00111101100: data <= 32'h3338372c;
    11'b00111101101: data <= 32'h38de34ea;
    11'b00111101110: data <= 32'hb0abb558;
    11'b00111101111: data <= 32'ha850ba31;
    11'b00111110000: data <= 32'h3d72312b;
    11'b00111110001: data <= 32'h407a3f2a;
    11'b00111110010: data <= 32'h3da43fe8;
    11'b00111110011: data <= 32'ha4403244;
    11'b00111110100: data <= 32'hb835bddf;
    11'b00111110101: data <= 32'hb490bd0f;
    11'b00111110110: data <= 32'hb31db440;
    11'b00111110111: data <= 32'hb103b851;
    11'b00111111000: data <= 32'h38b5bf63;
    11'b00111111001: data <= 32'h3d5fc008;
    11'b00111111010: data <= 32'h3959b56d;
    11'b00111111011: data <= 32'hbcbe3d51;
    11'b00111111100: data <= 32'hc0513d37;
    11'b00111111101: data <= 32'hbd2b3411;
    11'b00111111110: data <= 32'hb2acb464;
    11'b00111111111: data <= 32'hb8c5b1b9;
    11'b01000000000: data <= 32'hbe18b430;
    11'b01000000001: data <= 32'hbb0cb512;
    11'b01000000010: data <= 32'h3cd3382f;
    11'b01000000011: data <= 32'h40ab3f3f;
    11'b01000000100: data <= 32'h3d0b3fd4;
    11'b01000000101: data <= 32'hb6cc397e;
    11'b01000000110: data <= 32'hba14b4b0;
    11'b01000000111: data <= 32'h257c2eba;
    11'b01000001000: data <= 32'h38133874;
    11'b01000001001: data <= 32'h3831b875;
    11'b01000001010: data <= 32'h3b22c09f;
    11'b01000001011: data <= 32'h3dcdc0a2;
    11'b01000001100: data <= 32'h3c50b4d3;
    11'b01000001101: data <= 32'hb32d3d53;
    11'b01000001110: data <= 32'hbc053ab8;
    11'b01000001111: data <= 32'hb932b922;
    11'b01000010000: data <= 32'hb761bc84;
    11'b01000010001: data <= 32'hbdc0b8b9;
    11'b01000010010: data <= 32'hc090b52f;
    11'b01000010011: data <= 32'hbccdb800;
    11'b01000010100: data <= 32'h3c3eadec;
    11'b01000010101: data <= 32'h3f7e3c06;
    11'b01000010110: data <= 32'h362c3e5d;
    11'b01000010111: data <= 32'hbd233cba;
    11'b01000011000: data <= 32'hbc803abf;
    11'b01000011001: data <= 32'h30d93cd4;
    11'b01000011010: data <= 32'h39613c89;
    11'b01000011011: data <= 32'h352fb613;
    11'b01000011100: data <= 32'h3764c00d;
    11'b01000011101: data <= 32'h3d6cbeb2;
    11'b01000011110: data <= 32'h3f053631;
    11'b01000011111: data <= 32'h3c453e2d;
    11'b01000100000: data <= 32'h3412374e;
    11'b01000100001: data <= 32'h231abcc4;
    11'b01000100010: data <= 32'hb62bbd65;
    11'b01000100011: data <= 32'hbdddb7aa;
    11'b01000100100: data <= 32'hc010b641;
    11'b01000100101: data <= 32'hba98bce0;
    11'b01000100110: data <= 32'h3c45bd7f;
    11'b01000100111: data <= 32'h3d19b2f7;
    11'b01000101000: data <= 32'hb7a03c1a;
    11'b01000101001: data <= 32'hbf633d5a;
    11'b01000101010: data <= 32'hbce73d09;
    11'b01000101011: data <= 32'h2d4a3da3;
    11'b01000101100: data <= 32'h2e863c7c;
    11'b01000101101: data <= 32'hba26b206;
    11'b01000101110: data <= 32'hb89bbd48;
    11'b01000101111: data <= 32'h3c0bb95d;
    11'b01000110000: data <= 32'h40713c83;
    11'b01000110001: data <= 32'h3f883ee6;
    11'b01000110010: data <= 32'h3aee3624;
    11'b01000110011: data <= 32'h34d1bb8d;
    11'b01000110100: data <= 32'had25b8dc;
    11'b01000110101: data <= 32'hba5a346f;
    11'b01000110110: data <= 32'hbc5cb4b2;
    11'b01000110111: data <= 32'haf0ebfe8;
    11'b01000111000: data <= 32'h3cbac10f;
    11'b01000111001: data <= 32'h3bc0bc85;
    11'b01000111010: data <= 32'hb91d38af;
    11'b01000111011: data <= 32'hbe303c4c;
    11'b01000111100: data <= 32'hba4e3a37;
    11'b01000111101: data <= 32'h9e8a39a3;
    11'b01000111110: data <= 32'hba8a38e3;
    11'b01000111111: data <= 32'hc03daf3f;
    11'b01001000000: data <= 32'hbe92b9fa;
    11'b01001000001: data <= 32'h38a7af7a;
    11'b01001000010: data <= 32'h40583cfd;
    11'b01001000011: data <= 32'h3efb3e45;
    11'b01001000100: data <= 32'h381e386b;
    11'b01001000101: data <= 32'h2d2aaa99;
    11'b01001000110: data <= 32'h335839d7;
    11'b01001000111: data <= 32'h256d3d55;
    11'b01001001000: data <= 32'hb3e90eba;
    11'b01001001001: data <= 32'h34c0c086;
    11'b01001001010: data <= 32'h3cbfc1af;
    11'b01001001011: data <= 32'h3c59bcc1;
    11'b01001001100: data <= 32'h29ce383a;
    11'b01001001101: data <= 32'hb6eb38bf;
    11'b01001001110: data <= 32'h2deeb1a9;
    11'b01001001111: data <= 32'h2cffb47f;
    11'b01001010000: data <= 32'hbdd02e20;
    11'b01001010001: data <= 32'hc1c8aed9;
    11'b01001010010: data <= 32'hc032b966;
    11'b01001010011: data <= 32'h3536b774;
    11'b01001010100: data <= 32'h3eb037e5;
    11'b01001010101: data <= 32'h3aa53bc5;
    11'b01001010110: data <= 32'hb7103991;
    11'b01001010111: data <= 32'hb60d3ade;
    11'b01001011000: data <= 32'h36683f66;
    11'b01001011001: data <= 32'h366b402b;
    11'b01001011010: data <= 32'hb2363571;
    11'b01001011011: data <= 32'hac2abfa5;
    11'b01001011100: data <= 32'h3b0cc059;
    11'b01001011101: data <= 32'h3da4b70c;
    11'b01001011110: data <= 32'h3c623a85;
    11'b01001011111: data <= 32'h3ac531f8;
    11'b01001100000: data <= 32'h3bbdbb45;
    11'b01001100001: data <= 32'h35e1b9e5;
    11'b01001100010: data <= 32'hbd8c2fd6;
    11'b01001100011: data <= 32'hc144200d;
    11'b01001100100: data <= 32'hbed1bc35;
    11'b01001100101: data <= 32'h360bbdfb;
    11'b01001100110: data <= 32'h3c3ab9f8;
    11'b01001100111: data <= 32'hb1de315c;
    11'b01001101000: data <= 32'hbce238bb;
    11'b01001101001: data <= 32'hb8a03c9b;
    11'b01001101010: data <= 32'h37ae401e;
    11'b01001101011: data <= 32'h30dd4034;
    11'b01001101100: data <= 32'hbc1f3832;
    11'b01001101101: data <= 32'hbc6fbcbf;
    11'b01001101110: data <= 32'h348dbc2f;
    11'b01001101111: data <= 32'h3e5137fb;
    11'b01001110000: data <= 32'h3f0c3c6b;
    11'b01001110001: data <= 32'h3dee987c;
    11'b01001110010: data <= 32'h3d57bba7;
    11'b01001110011: data <= 32'h39b4b40a;
    11'b01001110100: data <= 32'hb9803af6;
    11'b01001110101: data <= 32'hbe5d35bb;
    11'b01001110110: data <= 32'hba89bdf4;
    11'b01001110111: data <= 32'h38d7c0f5;
    11'b01001111000: data <= 32'h3950bec9;
    11'b01001111001: data <= 32'hb8f0b67a;
    11'b01001111010: data <= 32'hbcb73379;
    11'b01001111011: data <= 32'hb15d3904;
    11'b01001111100: data <= 32'h390f3d20;
    11'b01001111101: data <= 32'hb6f83dcf;
    11'b01001111110: data <= 32'hc06337e1;
    11'b01001111111: data <= 32'hc072b865;
    11'b01010000000: data <= 32'hb52cb3da;
    11'b01010000001: data <= 32'h3d883b01;
    11'b01010000010: data <= 32'h3e3f3bfc;
    11'b01010000011: data <= 32'h3c56ab1d;
    11'b01010000100: data <= 32'h3c14b65e;
    11'b01010000101: data <= 32'h3b7a3b14;
    11'b01010000110: data <= 32'h31953fe9;
    11'b01010000111: data <= 32'hb8353aed;
    11'b01010001000: data <= 32'hb0eabe50;
    11'b01010001001: data <= 32'h3979c16c;
    11'b01010001010: data <= 32'h38b0bef1;
    11'b01010001011: data <= 32'hb430b6b3;
    11'b01010001100: data <= 32'hb46cb21e;
    11'b01010001101: data <= 32'h3a1ab5db;
    11'b01010001110: data <= 32'h3ba72e77;
    11'b01010001111: data <= 32'hbab23982;
    11'b01010010000: data <= 32'hc1bb366c;
    11'b01010010001: data <= 32'hc15fb4fb;
    11'b01010010010: data <= 32'hb8bab45f;
    11'b01010010011: data <= 32'h3b2c3592;
    11'b01010010100: data <= 32'h38dc35cc;
    11'b01010010101: data <= 32'ha8f9b153;
    11'b01010010110: data <= 32'h354a33e9;
    11'b01010010111: data <= 32'h3bf43f90;
    11'b01010011000: data <= 32'h39874187;
    11'b01010011001: data <= 32'hb1403d17;
    11'b01010011010: data <= 32'hb45ebcc8;
    11'b01010011011: data <= 32'h35c4bffd;
    11'b01010011100: data <= 32'h3939bac9;
    11'b01010011101: data <= 32'h38012c86;
    11'b01010011110: data <= 32'h3b01b7c2;
    11'b01010011111: data <= 32'h3ec8bcd6;
    11'b01010100000: data <= 32'h3d77b931;
    11'b01010100001: data <= 32'hb98a3757;
    11'b01010100010: data <= 32'hc11c380d;
    11'b01010100011: data <= 32'hc05eb712;
    11'b01010100100: data <= 32'hb5f7bbfe;
    11'b01010100101: data <= 32'h3627b9fe;
    11'b01010100110: data <= 32'hb802b820;
    11'b01010100111: data <= 32'hbc62b707;
    11'b01010101000: data <= 32'hb05b36ad;
    11'b01010101001: data <= 32'h3c234017;
    11'b01010101010: data <= 32'h395a416b;
    11'b01010101011: data <= 32'hb97f3d59;
    11'b01010101100: data <= 32'hbc9fb86f;
    11'b01010101101: data <= 32'hb50aba47;
    11'b01010101110: data <= 32'h38ed359d;
    11'b01010101111: data <= 32'h3c02390c;
    11'b01010110000: data <= 32'h3dcdb8de;
    11'b01010110001: data <= 32'h4011bdda;
    11'b01010110010: data <= 32'h3e96b7b4;
    11'b01010110011: data <= 32'haa213c18;
    11'b01010110100: data <= 32'hbdc03b6d;
    11'b01010110101: data <= 32'hbc3bb92d;
    11'b01010110110: data <= 32'h2fbebf22;
    11'b01010110111: data <= 32'h2cd2be86;
    11'b01010111000: data <= 32'hbc7abc65;
    11'b01010111001: data <= 32'hbd7dba55;
    11'b01010111010: data <= 32'h2c74ad9b;
    11'b01010111011: data <= 32'h3cf83ccb;
    11'b01010111100: data <= 32'h35303f66;
    11'b01010111101: data <= 32'hbe7d3c35;
    11'b01010111110: data <= 32'hc062a261;
    11'b01010111111: data <= 32'hbbbd31dc;
    11'b01011000000: data <= 32'h35db3c32;
    11'b01011000001: data <= 32'h3a423a05;
    11'b01011000010: data <= 32'h3bf0b98e;
    11'b01011000011: data <= 32'h3e2ebc98;
    11'b01011000100: data <= 32'h3e92367e;
    11'b01011000101: data <= 32'h39ba4015;
    11'b01011000110: data <= 32'hb31d3e06;
    11'b01011000111: data <= 32'hacbcb90c;
    11'b01011001000: data <= 32'h373fbfd1;
    11'b01011001001: data <= 32'ha097be77;
    11'b01011001010: data <= 32'hbc05bbdd;
    11'b01011001011: data <= 32'hb9ecbc21;
    11'b01011001100: data <= 32'h3b2abbed;
    11'b01011001101: data <= 32'h3e9aaf86;
    11'b01011001110: data <= 32'h2c843a2d;
    11'b01011001111: data <= 32'hc0653984;
    11'b01011010000: data <= 32'hc1363289;
    11'b01011010001: data <= 32'hbc9b3639;
    11'b01011010010: data <= 32'h21e73a7c;
    11'b01011010011: data <= 32'hae7733c9;
    11'b01011010100: data <= 32'hb40cbb28;
    11'b01011010101: data <= 32'h3874b979;
    11'b01011010110: data <= 32'h3db03d25;
    11'b01011010111: data <= 32'h3cbe4192;
    11'b01011011000: data <= 32'h35d13f80;
    11'b01011011001: data <= 32'h2f6ab539;
    11'b01011011010: data <= 32'h348cbd25;
    11'b01011011011: data <= 32'ha676b8f7;
    11'b01011011100: data <= 32'hb72db308;
    11'b01011011101: data <= 32'h3420bc33;
    11'b01011011110: data <= 32'h3f27bf15;
    11'b01011011111: data <= 32'h4022bc51;
    11'b01011100000: data <= 32'h322032e7;
    11'b01011100001: data <= 32'hbfa038d8;
    11'b01011100010: data <= 32'hc005307d;
    11'b01011100011: data <= 32'hb98baf4c;
    11'b01011100100: data <= 32'hb3c3aea6;
    11'b01011100101: data <= 32'hbc8eb8be;
    11'b01011100110: data <= 32'hbe0cbcd8;
    11'b01011100111: data <= 32'hb3ecb856;
    11'b01011101000: data <= 32'h3cf63dbb;
    11'b01011101001: data <= 32'h3cd4414f;
    11'b01011101010: data <= 32'h2caa3ef5;
    11'b01011101011: data <= 32'hb86f2d8c;
    11'b01011101100: data <= 32'hb564b08f;
    11'b01011101101: data <= 32'hb0463a28;
    11'b01011101110: data <= 32'ha5a73977;
    11'b01011101111: data <= 32'h3a68bb68;
    11'b01011110000: data <= 32'h4024c015;
    11'b01011110001: data <= 32'h4064bc98;
    11'b01011110010: data <= 32'h392c384e;
    11'b01011110011: data <= 32'hbad03b9b;
    11'b01011110100: data <= 32'hb9a32552;
    11'b01011110101: data <= 32'h3083ba41;
    11'b01011110110: data <= 32'hb493bb6d;
    11'b01011110111: data <= 32'hbf06bc8f;
    11'b01011111000: data <= 32'hc00ebddc;
    11'b01011111001: data <= 32'hb508bb38;
    11'b01011111010: data <= 32'h3d5e391b;
    11'b01011111011: data <= 32'h3b983e86;
    11'b01011111100: data <= 32'hb9b43c83;
    11'b01011111101: data <= 32'hbe0735af;
    11'b01011111110: data <= 32'hbbbc3a78;
    11'b01011111111: data <= 32'hb5623ed7;
    11'b01100000000: data <= 32'hb0b73c6d;
    11'b01100000001: data <= 32'h361fbafb;
    11'b01100000010: data <= 32'h3dc5bf3b;
    11'b01100000011: data <= 32'h3f8fb6f7;
    11'b01100000100: data <= 32'h3c903dc6;
    11'b01100000101: data <= 32'h35663e0a;
    11'b01100000110: data <= 32'h38312853;
    11'b01100000111: data <= 32'h3a6abbfc;
    11'b01100001000: data <= 32'hb24ebb83;
    11'b01100001001: data <= 32'hbed6bb4b;
    11'b01100001010: data <= 32'hbe5bbdc6;
    11'b01100001011: data <= 32'h35e5be36;
    11'b01100001100: data <= 32'h3eeab927;
    11'b01100001101: data <= 32'h39cf34f9;
    11'b01100001110: data <= 32'hbd29369f;
    11'b01100001111: data <= 32'hbfb935d9;
    11'b01100010000: data <= 32'hbc453c47;
    11'b01100010001: data <= 32'hb79d3ec0;
    11'b01100010010: data <= 32'hba723a33;
    11'b01100010011: data <= 32'hba9cbc26;
    11'b01100010100: data <= 32'h3311bd97;
    11'b01100010101: data <= 32'h3d3a3684;
    11'b01100010110: data <= 32'h3d82405c;
    11'b01100010111: data <= 32'h3bb73f4b;
    11'b01100011000: data <= 32'h3b993195;
    11'b01100011001: data <= 32'h3aceb828;
    11'b01100011010: data <= 32'hb0f92557;
    11'b01100011011: data <= 32'hbce22c5c;
    11'b01100011100: data <= 32'hb94fbc68;
    11'b01100011101: data <= 32'h3cf5c029;
    11'b01100011110: data <= 32'h4039be8a;
    11'b01100011111: data <= 32'h39dcb7fd;
    11'b01100100000: data <= 32'hbc992c7b;
    11'b01100100001: data <= 32'hbd7932ce;
    11'b01100100010: data <= 32'hb6a83923;
    11'b01100100011: data <= 32'hb63a3b08;
    11'b01100100100: data <= 32'hbe5aa4a1;
    11'b01100100101: data <= 32'hc035bd5b;
    11'b01100100110: data <= 32'hbacebcbf;
    11'b01100100111: data <= 32'h3a9b3958;
    11'b01100101000: data <= 32'h3d17402a;
    11'b01100101001: data <= 32'h3a003e19;
    11'b01100101010: data <= 32'h36b83468;
    11'b01100101011: data <= 32'h34d53603;
    11'b01100101100: data <= 32'hb41e3db2;
    11'b01100101101: data <= 32'hba223cfb;
    11'b01100101110: data <= 32'ha970b92c;
    11'b01100101111: data <= 32'h3e39c063;
    11'b01100110000: data <= 32'h4038bf1a;
    11'b01100110001: data <= 32'h3b4db59b;
    11'b01100110010: data <= 32'hb54134de;
    11'b01100110011: data <= 32'haadf2d3d;
    11'b01100110100: data <= 32'h398ba525;
    11'b01100110101: data <= 32'had212245;
    11'b01100110110: data <= 32'hc009b8c7;
    11'b01100110111: data <= 32'hc15fbe00;
    11'b01100111000: data <= 32'hbc7dbd43;
    11'b01100111001: data <= 32'h3a2c2da5;
    11'b01100111010: data <= 32'h3be53c3b;
    11'b01100111011: data <= 32'h9f4a3928;
    11'b01100111100: data <= 32'hb84e31d0;
    11'b01100111101: data <= 32'hb5a53c7b;
    11'b01100111110: data <= 32'hb66e40dc;
    11'b01100111111: data <= 32'hb9ab3f9e;
    11'b01101000000: data <= 32'hb44db645;
    11'b01101000001: data <= 32'h3b7bbf9f;
    11'b01101000010: data <= 32'h3e3abc6d;
    11'b01101000011: data <= 32'h3c303831;
    11'b01101000100: data <= 32'h39233afb;
    11'b01101000101: data <= 32'h3cf62c01;
    11'b01101000110: data <= 32'h3e79b5fa;
    11'b01101000111: data <= 32'h3415b145;
    11'b01101001000: data <= 32'hbf8fb63f;
    11'b01101001001: data <= 32'hc09cbd0a;
    11'b01101001010: data <= 32'hb80fbe7c;
    11'b01101001011: data <= 32'h3c92bbc4;
    11'b01101001100: data <= 32'h39f7b537;
    11'b01101001101: data <= 32'hb972b5b4;
    11'b01101001110: data <= 32'hbc67ae23;
    11'b01101001111: data <= 32'hb7ca3d17;
    11'b01101010000: data <= 32'hb5c640f3;
    11'b01101010001: data <= 32'hbc333eb9;
    11'b01101010010: data <= 32'hbd05b812;
    11'b01101010011: data <= 32'hb57dbdec;
    11'b01101010100: data <= 32'h3962b277;
    11'b01101010101: data <= 32'h3baf3d7e;
    11'b01101010110: data <= 32'h3c8a3ce9;
    11'b01101010111: data <= 32'h3efb2bf4;
    11'b01101011000: data <= 32'h3f46b1a1;
    11'b01101011001: data <= 32'h362838a4;
    11'b01101011010: data <= 32'hbd883913;
    11'b01101011011: data <= 32'hbd61b8f3;
    11'b01101011100: data <= 32'h3725bf37;
    11'b01101011101: data <= 32'h3e49bf38;
    11'b01101011110: data <= 32'h392dbce7;
    11'b01101011111: data <= 32'hba42bb2f;
    11'b01101100000: data <= 32'hb9f0b625;
    11'b01101100001: data <= 32'h323b3a84;
    11'b01101100010: data <= 32'h228b3ea2;
    11'b01101100011: data <= 32'hbdeb3ab1;
    11'b01101100100: data <= 32'hc0b8bad4;
    11'b01101100101: data <= 32'hbe0bbcc8;
    11'b01101100110: data <= 32'haa37343c;
    11'b01101100111: data <= 32'h395e3ddf;
    11'b01101101000: data <= 32'h3afa3b55;
    11'b01101101001: data <= 32'h3cefae69;
    11'b01101101010: data <= 32'h3d0835f4;
    11'b01101101011: data <= 32'h340b3f35;
    11'b01101101100: data <= 32'hbb073fa5;
    11'b01101101101: data <= 32'hb86b2f21;
    11'b01101101110: data <= 32'h3b8dbebc;
    11'b01101101111: data <= 32'h3e51bf81;
    11'b01101110000: data <= 32'h38c1bc7a;
    11'b01101110001: data <= 32'hb4b4b998;
    11'b01101110010: data <= 32'h362cb815;
    11'b01101110011: data <= 32'h3d9d2f85;
    11'b01101110100: data <= 32'h38f5393a;
    11'b01101110101: data <= 32'hbe8c2daf;
    11'b01101110110: data <= 32'hc1b5bc2e;
    11'b01101110111: data <= 32'hbf65bc82;
    11'b01101111000: data <= 32'hb20f95c7;
    11'b01101111001: data <= 32'h35a1390e;
    11'b01101111010: data <= 32'h2d78ab24;
    11'b01101111011: data <= 32'h3171b808;
    11'b01101111100: data <= 32'h37463a88;
    11'b01101111101: data <= 32'h2bc94167;
    11'b01101111110: data <= 32'hb9484151;
    11'b01101111111: data <= 32'hb7d0380a;
    11'b01110000000: data <= 32'h3824bd46;
    11'b01110000001: data <= 32'h3b96bcb2;
    11'b01110000010: data <= 32'h36b2b17d;
    11'b01110000011: data <= 32'h35bba114;
    11'b01110000100: data <= 32'h3e41b798;
    11'b01110000101: data <= 32'h40dfb5c6;
    11'b01110000110: data <= 32'h3c9332d1;
    11'b01110000111: data <= 32'hbd8c2e23;
    11'b01110001000: data <= 32'hc0dcba02;
    11'b01110001001: data <= 32'hbcc4bc8a;
    11'b01110001010: data <= 32'h3442b9dc;
    11'b01110001011: data <= 32'h3124b8ff;
    11'b01110001100: data <= 32'hb97bbcbb;
    11'b01110001101: data <= 32'hb906bc10;
    11'b01110001110: data <= 32'h2f963a6b;
    11'b01110001111: data <= 32'h30114165;
    11'b01110010000: data <= 32'hb9d240d9;
    11'b01110010001: data <= 32'hbc95358e;
    11'b01110010010: data <= 32'hb8f9bb69;
    11'b01110010011: data <= 32'hac7db21c;
    11'b01110010100: data <= 32'h2b9d3b14;
    11'b01110010101: data <= 32'h3927385b;
    11'b01110010110: data <= 32'h4006b790;
    11'b01110010111: data <= 32'h4154b681;
    11'b01110011000: data <= 32'h3d223915;
    11'b01110011001: data <= 32'hbb163bc0;
    11'b01110011010: data <= 32'hbd9d25a5;
    11'b01110011011: data <= 32'hab4ebc14;
    11'b01110011100: data <= 32'h3b16bd4d;
    11'b01110011101: data <= 32'h2d8cbdda;
    11'b01110011110: data <= 32'hbbfcbf28;
    11'b01110011111: data <= 32'hb8a5bd7b;
    11'b01110100000: data <= 32'h39133514;
    11'b01110100001: data <= 32'h38f23f4a;
    11'b01110100010: data <= 32'hbac93db8;
    11'b01110100011: data <= 32'hbfedb188;
    11'b01110100100: data <= 32'hbee3b973;
    11'b01110100101: data <= 32'hbb223756;
    11'b01110100110: data <= 32'hb5ad3d1d;
    11'b01110100111: data <= 32'h350e369c;
    11'b01110101000: data <= 32'h3dccb9d9;
    11'b01110101001: data <= 32'h3ff5b142;
    11'b01110101010: data <= 32'h3c013e49;
    11'b01110101011: data <= 32'hb6d54056;
    11'b01110101100: data <= 32'hb73f3b09;
    11'b01110101101: data <= 32'h39cfb9c2;
    11'b01110101110: data <= 32'h3c5abd29;
    11'b01110101111: data <= 32'ha88ebd3e;
    11'b01110110000: data <= 32'hba6fbe12;
    11'b01110110001: data <= 32'h3406bd8a;
    11'b01110110010: data <= 32'h3f06b568;
    11'b01110110011: data <= 32'h3d7a3974;
    11'b01110110100: data <= 32'hba403695;
    11'b01110110101: data <= 32'hc0a9b891;
    11'b01110110110: data <= 32'hc008b893;
    11'b01110110111: data <= 32'hbc063785;
    11'b01110111000: data <= 32'hb8e639f5;
    11'b01110111001: data <= 32'hb71ab756;
    11'b01110111010: data <= 32'h344fbd25;
    11'b01110111011: data <= 32'h3b7a25e4;
    11'b01110111100: data <= 32'h38c44096;
    11'b01110111101: data <= 32'hb24341c1;
    11'b01110111110: data <= 32'hb0313d2c;
    11'b01110111111: data <= 32'h38dfb5c1;
    11'b01111000000: data <= 32'h389bb8b9;
    11'b01111000001: data <= 32'hb5c2b437;
    11'b01111000010: data <= 32'hb6e5b8d9;
    11'b01111000011: data <= 32'h3ce8bc8f;
    11'b01111000100: data <= 32'h4182ba73;
    11'b01111000101: data <= 32'h3fd41cf9;
    11'b01111000110: data <= 32'hb7a92eb0;
    11'b01111000111: data <= 32'hbf85b6ba;
    11'b01111001000: data <= 32'hbd19b71d;
    11'b01111001001: data <= 32'hb5d327bc;
    11'b01111001010: data <= 32'hb8e5b49a;
    11'b01111001011: data <= 32'hbcc3be35;
    11'b01111001100: data <= 32'hb9f3bf9a;
    11'b01111001101: data <= 32'h3486ae3e;
    11'b01111001110: data <= 32'h37df4077;
    11'b01111001111: data <= 32'hb0de4125;
    11'b01111010000: data <= 32'hb7e53bed;
    11'b01111010001: data <= 32'hb491b020;
    11'b01111010010: data <= 32'hb67d35e0;
    11'b01111010011: data <= 32'hbad33be8;
    11'b01111010100: data <= 32'hb4cc3427;
    11'b01111010101: data <= 32'h3e5dbb8e;
    11'b01111010110: data <= 32'h41dbbb7a;
    11'b01111010111: data <= 32'h4000305b;
    11'b01111011000: data <= 32'hae5939b2;
    11'b01111011001: data <= 32'hbafb34d4;
    11'b01111011010: data <= 32'h28d7b1a1;
    11'b01111011011: data <= 32'h3874b5d7;
    11'b01111011100: data <= 32'hb7a2bc10;
    11'b01111011101: data <= 32'hbe3dc040;
    11'b01111011110: data <= 32'hbbd4c06c;
    11'b01111011111: data <= 32'h381eb811;
    11'b01111100000: data <= 32'h3b483d75;
    11'b01111100001: data <= 32'haf403dad;
    11'b01111100010: data <= 32'hbc6531fc;
    11'b01111100011: data <= 32'hbd00ae44;
    11'b01111100100: data <= 32'hbcd73c34;
    11'b01111100101: data <= 32'hbd1c3e9d;
    11'b01111100110: data <= 32'hb8da36dd;
    11'b01111100111: data <= 32'h3c15bc69;
    11'b01111101000: data <= 32'h403bbac2;
    11'b01111101001: data <= 32'h3dd93a8d;
    11'b01111101010: data <= 32'h30ce3f02;
    11'b01111101011: data <= 32'h2e493c9c;
    11'b01111101100: data <= 32'h3c5731e5;
    11'b01111101101: data <= 32'h3c4cb4c5;
    11'b01111101110: data <= 32'hb786bab7;
    11'b01111101111: data <= 32'hbe03befa;
    11'b01111110000: data <= 32'hb69bc004;
    11'b01111110001: data <= 32'h3dcfbbc3;
    11'b01111110010: data <= 32'h3ea032d2;
    11'b01111110011: data <= 32'h2ac930ac;
    11'b01111110100: data <= 32'hbd76b850;
    11'b01111110101: data <= 32'hbe04b0ac;
    11'b01111110110: data <= 32'hbcfa3cba;
    11'b01111110111: data <= 32'hbd783d96;
    11'b01111111000: data <= 32'hbcceb380;
    11'b01111111001: data <= 32'hb14dbe95;
    11'b01111111010: data <= 32'h3a91ba46;
    11'b01111111011: data <= 32'h39c73daa;
    11'b01111111100: data <= 32'h325e40cd;
    11'b01111111101: data <= 32'h382a3e0f;
    11'b01111111110: data <= 32'h3d0236ea;
    11'b01111111111: data <= 32'h3a61346d;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    