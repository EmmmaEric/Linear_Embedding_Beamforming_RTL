
module memory_rom_41(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hba743d71;
    11'b00000000001: data <= 32'hb6923a78;
    11'b00000000010: data <= 32'h37eeba32;
    11'b00000000011: data <= 32'h3e4cbc0e;
    11'b00000000100: data <= 32'h3e4139d1;
    11'b00000000101: data <= 32'h3737409d;
    11'b00000000110: data <= 32'hb0ee3f66;
    11'b00000000111: data <= 32'h38243187;
    11'b00000001000: data <= 32'h3c43baaa;
    11'b00000001001: data <= 32'h318ebb69;
    11'b00000001010: data <= 32'hbc16bc97;
    11'b00000001011: data <= 32'hb7bdbe53;
    11'b00000001100: data <= 32'h3db9bd0f;
    11'b00000001101: data <= 32'h4051b27b;
    11'b00000001110: data <= 32'h383b3512;
    11'b00000001111: data <= 32'hbe6ab12e;
    11'b00000010000: data <= 32'hc02ab68f;
    11'b00000010001: data <= 32'hbcff35d3;
    11'b00000010010: data <= 32'hba643b71;
    11'b00000010011: data <= 32'hbbe9aa4d;
    11'b00000010100: data <= 32'hb97abdf9;
    11'b00000010101: data <= 32'h351bbc68;
    11'b00000010110: data <= 32'h3add3cbd;
    11'b00000010111: data <= 32'h3727419f;
    11'b00000011000: data <= 32'h2e58402e;
    11'b00000011001: data <= 32'h37363607;
    11'b00000011010: data <= 32'h3886b2af;
    11'b00000011011: data <= 32'hb4ae330c;
    11'b00000011100: data <= 32'hbb4a2ab4;
    11'b00000011101: data <= 32'h33bcbbb8;
    11'b00000011110: data <= 32'h4093bdc6;
    11'b00000011111: data <= 32'h4163ba2f;
    11'b00000100000: data <= 32'h3a84a7c1;
    11'b00000100001: data <= 32'hbc77ab65;
    11'b00000100010: data <= 32'hbcacb2bd;
    11'b00000100011: data <= 32'hb4482f66;
    11'b00000100100: data <= 32'hb6432db1;
    11'b00000100101: data <= 32'hbdbebc48;
    11'b00000100110: data <= 32'hbe72c054;
    11'b00000100111: data <= 32'hb6babd5b;
    11'b00000101000: data <= 32'h39153be0;
    11'b00000101001: data <= 32'h37854098;
    11'b00000101010: data <= 32'hb1733dd5;
    11'b00000101011: data <= 32'hb55c3325;
    11'b00000101100: data <= 32'hb68a37ac;
    11'b00000101101: data <= 32'hbb533dc6;
    11'b00000101110: data <= 32'hbbe13c63;
    11'b00000101111: data <= 32'h3663b85e;
    11'b00000110000: data <= 32'h4080bdcf;
    11'b00000110001: data <= 32'h40f1b92f;
    11'b00000110010: data <= 32'h3b31384d;
    11'b00000110011: data <= 32'hb4d239a3;
    11'b00000110100: data <= 32'h321c32f9;
    11'b00000110101: data <= 32'h3b6faa8e;
    11'b00000110110: data <= 32'h2d1cb6bc;
    11'b00000110111: data <= 32'hbe5bbddb;
    11'b00000111000: data <= 32'hbf31c09d;
    11'b00000111001: data <= 32'hb29cbe58;
    11'b00000111010: data <= 32'h3c643238;
    11'b00000111011: data <= 32'h39413c12;
    11'b00000111100: data <= 32'hb89c34f7;
    11'b00000111101: data <= 32'hbc83b12b;
    11'b00000111110: data <= 32'hbc6b3b0a;
    11'b00000111111: data <= 32'hbd1c4015;
    11'b00001000000: data <= 32'hbd0b3d47;
    11'b00001000001: data <= 32'hb2dfb984;
    11'b00001000010: data <= 32'h3cf6bdd1;
    11'b00001000011: data <= 32'h3e3faed4;
    11'b00001000100: data <= 32'h39ba3ded;
    11'b00001000101: data <= 32'h35ed3e2a;
    11'b00001000110: data <= 32'h3cbf38f7;
    11'b00001000111: data <= 32'h3e4a2dc2;
    11'b00001001000: data <= 32'h32b3af61;
    11'b00001001001: data <= 32'hbe1cbac1;
    11'b00001001010: data <= 32'hbd36befd;
    11'b00001001011: data <= 32'h399abea6;
    11'b00001001100: data <= 32'h3fa5b9ab;
    11'b00001001101: data <= 32'h3ba0b424;
    11'b00001001110: data <= 32'hb99eb909;
    11'b00001001111: data <= 32'hbce4b74a;
    11'b00001010000: data <= 32'hbb4f3b19;
    11'b00001010001: data <= 32'hbc433f22;
    11'b00001010010: data <= 32'hbe3d393a;
    11'b00001010011: data <= 32'hbd00bd54;
    11'b00001010100: data <= 32'hb0bbbe46;
    11'b00001010101: data <= 32'h382b3529;
    11'b00001010110: data <= 32'h36b33ff8;
    11'b00001010111: data <= 32'h38913efe;
    11'b00001011000: data <= 32'h3d2f3951;
    11'b00001011001: data <= 32'h3d2f379f;
    11'b00001011010: data <= 32'hb0fb3b2d;
    11'b00001011011: data <= 32'hbdce37a8;
    11'b00001011100: data <= 32'hb925ba5f;
    11'b00001011101: data <= 32'h3e21be1b;
    11'b00001011110: data <= 32'h40d7bcce;
    11'b00001011111: data <= 32'h3c7fba4b;
    11'b00001100000: data <= 32'hb67eba43;
    11'b00001100001: data <= 32'hb6cfb640;
    11'b00001100010: data <= 32'h31b23961;
    11'b00001100011: data <= 32'hb5633c28;
    11'b00001100100: data <= 32'hbeb9b509;
    11'b00001100101: data <= 32'hc029bff0;
    11'b00001100110: data <= 32'hbc47beef;
    11'b00001100111: data <= 32'h2023343a;
    11'b00001101000: data <= 32'h34463e4e;
    11'b00001101001: data <= 32'h35313c15;
    11'b00001101010: data <= 32'h391132d4;
    11'b00001101011: data <= 32'h36823ac2;
    11'b00001101100: data <= 32'hba124006;
    11'b00001101101: data <= 32'hbdf83ed1;
    11'b00001101110: data <= 32'hb641ab78;
    11'b00001101111: data <= 32'h3e4bbd45;
    11'b00001110000: data <= 32'h403ebc53;
    11'b00001110001: data <= 32'h3b8bb5cc;
    11'b00001110010: data <= 32'h2ee0b083;
    11'b00001110011: data <= 32'h3a94203c;
    11'b00001110100: data <= 32'h3e373807;
    11'b00001110101: data <= 32'h379737a9;
    11'b00001110110: data <= 32'hbe54ba26;
    11'b00001110111: data <= 32'hc080c024;
    11'b00001111000: data <= 32'hbc11bf06;
    11'b00001111001: data <= 32'h34f2b402;
    11'b00001111010: data <= 32'h3670367d;
    11'b00001111011: data <= 32'hac1ab4d4;
    11'b00001111100: data <= 32'hb164b82f;
    11'b00001111101: data <= 32'hb5463bb7;
    11'b00001111110: data <= 32'hbc5c4127;
    11'b00001111111: data <= 32'hbe5c4034;
    11'b00010000000: data <= 32'hba190ed6;
    11'b00010000001: data <= 32'h395cbcf2;
    11'b00010000010: data <= 32'h3c31b884;
    11'b00010000011: data <= 32'h3684386d;
    11'b00010000100: data <= 32'h37ae39b0;
    11'b00010000101: data <= 32'h3f14365c;
    11'b00010000110: data <= 32'h40c7381e;
    11'b00010000111: data <= 32'h3ac938a5;
    11'b00010001000: data <= 32'hbd98b405;
    11'b00010001001: data <= 32'hbf1dbd78;
    11'b00010001010: data <= 32'hb16abdf7;
    11'b00010001011: data <= 32'h3c6fbac4;
    11'b00010001100: data <= 32'h398cba82;
    11'b00010001101: data <= 32'hb46abdca;
    11'b00010001110: data <= 32'hb6d2bc68;
    11'b00010001111: data <= 32'hb38a3a7f;
    11'b00010010000: data <= 32'hba1440ab;
    11'b00010010001: data <= 32'hbe4b3e19;
    11'b00010010010: data <= 32'hbdf9b8c1;
    11'b00010010011: data <= 32'hb939bd5f;
    11'b00010010100: data <= 32'hb2adad5b;
    11'b00010010101: data <= 32'hb2c23cc0;
    11'b00010010110: data <= 32'h37bb3c08;
    11'b00010010111: data <= 32'h3f8e35a8;
    11'b00010011000: data <= 32'h407638fb;
    11'b00010011001: data <= 32'h388f3d35;
    11'b00010011010: data <= 32'hbd373bfe;
    11'b00010011011: data <= 32'hbc5eb25f;
    11'b00010011100: data <= 32'h3a01bc07;
    11'b00010011101: data <= 32'h3eccbc6d;
    11'b00010011110: data <= 32'h3a70bd5f;
    11'b00010011111: data <= 32'hb2e6bf01;
    11'b00010100000: data <= 32'h2e96bcad;
    11'b00010100001: data <= 32'h3a3b3872;
    11'b00010100010: data <= 32'h31b33e51;
    11'b00010100011: data <= 32'hbd563806;
    11'b00010100100: data <= 32'hc021bd42;
    11'b00010100101: data <= 32'hbe46bde5;
    11'b00010100110: data <= 32'hbb3a2a87;
    11'b00010100111: data <= 32'hb85f3c0e;
    11'b00010101000: data <= 32'h314a35cd;
    11'b00010101001: data <= 32'h3ceab4a1;
    11'b00010101010: data <= 32'h3d4a3910;
    11'b00010101011: data <= 32'had544049;
    11'b00010101100: data <= 32'hbd50406c;
    11'b00010101101: data <= 32'hb97d39fb;
    11'b00010101110: data <= 32'h3c07b882;
    11'b00010101111: data <= 32'h3df3bb09;
    11'b00010110000: data <= 32'h374fbb6f;
    11'b00010110001: data <= 32'ha9ccbc84;
    11'b00010110010: data <= 32'h3c49b9fd;
    11'b00010110011: data <= 32'h4045361d;
    11'b00010110100: data <= 32'h3cdf3b38;
    11'b00010110101: data <= 32'hbba3b07f;
    11'b00010110110: data <= 32'hc02ebdfd;
    11'b00010110111: data <= 32'hbe1fbd70;
    11'b00010111000: data <= 32'hb94eb0a1;
    11'b00010111001: data <= 32'hb6da2f9e;
    11'b00010111010: data <= 32'hb357bb7d;
    11'b00010111011: data <= 32'h3579bd10;
    11'b00010111100: data <= 32'h36c636ff;
    11'b00010111101: data <= 32'hb821410e;
    11'b00010111110: data <= 32'hbd4c4141;
    11'b00010111111: data <= 32'hba273b46;
    11'b00011000000: data <= 32'h35f9b6b0;
    11'b00011000001: data <= 32'h3723b57d;
    11'b00011000010: data <= 32'hb52629db;
    11'b00011000011: data <= 32'ha1cdb0ac;
    11'b00011000100: data <= 32'h3f44b41c;
    11'b00011000101: data <= 32'h41fb3530;
    11'b00011000110: data <= 32'h3ef13a02;
    11'b00011000111: data <= 32'hb93d2f67;
    11'b00011001000: data <= 32'hbe4dbab4;
    11'b00011001001: data <= 32'hb926bae3;
    11'b00011001010: data <= 32'h3370b63a;
    11'b00011001011: data <= 32'ha9bbbb07;
    11'b00011001100: data <= 32'hb7bbc037;
    11'b00011001101: data <= 32'hb03dc00e;
    11'b00011001110: data <= 32'h34482f6b;
    11'b00011001111: data <= 32'hb3fb406f;
    11'b00011010000: data <= 32'hbc5f400d;
    11'b00011010001: data <= 32'hbc98341e;
    11'b00011010010: data <= 32'hb9b8b8c4;
    11'b00011010011: data <= 32'hbab6313c;
    11'b00011010100: data <= 32'hbca33ae5;
    11'b00011010101: data <= 32'hb341362d;
    11'b00011010110: data <= 32'h3f5bb2fe;
    11'b00011010111: data <= 32'h41a733f5;
    11'b00011011000: data <= 32'h3dc63c88;
    11'b00011011001: data <= 32'hb8cc3c7c;
    11'b00011011010: data <= 32'hbaf235ac;
    11'b00011011011: data <= 32'h36ddb032;
    11'b00011011100: data <= 32'h3c29b635;
    11'b00011011101: data <= 32'h3145bd26;
    11'b00011011110: data <= 32'hb893c0d8;
    11'b00011011111: data <= 32'h2cf5c043;
    11'b00011100000: data <= 32'h3c20b078;
    11'b00011100001: data <= 32'h399f3dc2;
    11'b00011100010: data <= 32'hb8c43b05;
    11'b00011100011: data <= 32'hbdb0b947;
    11'b00011100100: data <= 32'hbdf1baac;
    11'b00011100101: data <= 32'hbe4236a3;
    11'b00011100110: data <= 32'hbe543bdc;
    11'b00011100111: data <= 32'hb8bb9e72;
    11'b00011101000: data <= 32'h3c96bade;
    11'b00011101001: data <= 32'h3f43189b;
    11'b00011101010: data <= 32'h38f33e9d;
    11'b00011101011: data <= 32'hb9e04056;
    11'b00011101100: data <= 32'hb5f93d64;
    11'b00011101101: data <= 32'h3ba5373d;
    11'b00011101110: data <= 32'h3c55abbd;
    11'b00011101111: data <= 32'hb11cba9e;
    11'b00011110000: data <= 32'hb929bee7;
    11'b00011110001: data <= 32'h39babe4b;
    11'b00011110010: data <= 32'h406ab2c0;
    11'b00011110011: data <= 32'h3f31398f;
    11'b00011110100: data <= 32'ha7cda30b;
    11'b00011110101: data <= 32'hbd2ebc64;
    11'b00011110110: data <= 32'hbd89ba23;
    11'b00011110111: data <= 32'hbd1e3711;
    11'b00011111000: data <= 32'hbd7d36b4;
    11'b00011111001: data <= 32'hbb3abc71;
    11'b00011111010: data <= 32'h32a3bf94;
    11'b00011111011: data <= 32'h398cb6a1;
    11'b00011111100: data <= 32'hac6d3f5c;
    11'b00011111101: data <= 32'hba6a4101;
    11'b00011111110: data <= 32'hb4283dfa;
    11'b00011111111: data <= 32'h3930387c;
    11'b00100000000: data <= 32'h33f436d1;
    11'b00100000001: data <= 32'hbbf43227;
    11'b00100000010: data <= 32'hbad8b85c;
    11'b00100000011: data <= 32'h3ce6baac;
    11'b00100000100: data <= 32'h41eeb197;
    11'b00100000101: data <= 32'h40a83602;
    11'b00100000110: data <= 32'h349facef;
    11'b00100000111: data <= 32'hba4eb949;
    11'b00100001000: data <= 32'hb741b330;
    11'b00100001001: data <= 32'hb2dc3742;
    11'b00100001010: data <= 32'hba14b509;
    11'b00100001011: data <= 32'hbc32c058;
    11'b00100001100: data <= 32'hb683c165;
    11'b00100001101: data <= 32'h334bba7d;
    11'b00100001110: data <= 32'ha95c3df6;
    11'b00100001111: data <= 32'hb8653f6a;
    11'b00100010000: data <= 32'hb61d39a2;
    11'b00100010001: data <= 32'hb0ef31dd;
    11'b00100010010: data <= 32'hbb533a97;
    11'b00100010011: data <= 32'hbf953c80;
    11'b00100010100: data <= 32'hbccb3488;
    11'b00100010101: data <= 32'h3ca8b851;
    11'b00100010110: data <= 32'h417eb3c9;
    11'b00100010111: data <= 32'h3fbb3814;
    11'b00100011000: data <= 32'h31e03905;
    11'b00100011001: data <= 32'hb1b13654;
    11'b00100011010: data <= 32'h39c138af;
    11'b00100011011: data <= 32'h3afd3908;
    11'b00100011100: data <= 32'hb489b8c8;
    11'b00100011101: data <= 32'hbc67c0dd;
    11'b00100011110: data <= 32'hb6d2c178;
    11'b00100011111: data <= 32'h3971bba2;
    11'b00100100000: data <= 32'h3a083a4d;
    11'b00100100001: data <= 32'h283638ec;
    11'b00100100010: data <= 32'hb71eb79c;
    11'b00100100011: data <= 32'hba16b533;
    11'b00100100100: data <= 32'hbe543c0d;
    11'b00100100101: data <= 32'hc0973dd0;
    11'b00100100110: data <= 32'hbe0532a8;
    11'b00100100111: data <= 32'h3824bc00;
    11'b00100101000: data <= 32'h3e9fb887;
    11'b00100101001: data <= 32'h3af23a5e;
    11'b00100101010: data <= 32'hb2e63de8;
    11'b00100101011: data <= 32'h33933d4d;
    11'b00100101100: data <= 32'h3dbc3cbf;
    11'b00100101101: data <= 32'h3cf23ba9;
    11'b00100101110: data <= 32'hb677b0d0;
    11'b00100101111: data <= 32'hbcedbea6;
    11'b00100110000: data <= 32'ha81fbfdd;
    11'b00100110001: data <= 32'h3e84ba37;
    11'b00100110010: data <= 32'h3f1d303d;
    11'b00100110011: data <= 32'h3934b72b;
    11'b00100110100: data <= 32'hb422bcf2;
    11'b00100110101: data <= 32'hb914b7c8;
    11'b00100110110: data <= 32'hbcf03c4b;
    11'b00100110111: data <= 32'hbfa73c8a;
    11'b00100111000: data <= 32'hbe64b92e;
    11'b00100111001: data <= 32'hb54cbfcf;
    11'b00100111010: data <= 32'h3601bc3c;
    11'b00100111011: data <= 32'hb0973af9;
    11'b00100111100: data <= 32'hb8473efe;
    11'b00100111101: data <= 32'h35bb3dad;
    11'b00100111110: data <= 32'h3d793cad;
    11'b00100111111: data <= 32'h395e3d11;
    11'b00101000000: data <= 32'hbc8d3a4e;
    11'b00101000001: data <= 32'hbe20b56b;
    11'b00101000010: data <= 32'h3530bb46;
    11'b00101000011: data <= 32'h4095b787;
    11'b00101000100: data <= 32'h4087b169;
    11'b00101000101: data <= 32'h3b23b9fa;
    11'b00101000110: data <= 32'h2fedbc5b;
    11'b00101000111: data <= 32'h3376ac58;
    11'b00101001000: data <= 32'ha9643cb6;
    11'b00101001001: data <= 32'hbbfe38ac;
    11'b00101001010: data <= 32'hbdddbe56;
    11'b00101001011: data <= 32'hbb3cc16f;
    11'b00101001100: data <= 32'hb518bdb3;
    11'b00101001101: data <= 32'hb6d338bc;
    11'b00101001110: data <= 32'hb6fb3c8d;
    11'b00101001111: data <= 32'h35223821;
    11'b00101010000: data <= 32'h3a2d3823;
    11'b00101010001: data <= 32'hb5723d92;
    11'b00101010010: data <= 32'hc0023ea7;
    11'b00101010011: data <= 32'hbf8c39ab;
    11'b00101010100: data <= 32'h347bb492;
    11'b00101010101: data <= 32'h402cb59d;
    11'b00101010110: data <= 32'h3f16aea0;
    11'b00101010111: data <= 32'h3864b440;
    11'b00101011000: data <= 32'h37b6b2d1;
    11'b00101011001: data <= 32'h3d5e39a2;
    11'b00101011010: data <= 32'h3d043d9a;
    11'b00101011011: data <= 32'hb1ce355b;
    11'b00101011100: data <= 32'hbd2fbf54;
    11'b00101011101: data <= 32'hbbc2c15a;
    11'b00101011110: data <= 32'hae69bd7e;
    11'b00101011111: data <= 32'h310f2f06;
    11'b00101100000: data <= 32'h2e1da915;
    11'b00101100001: data <= 32'h3553bae3;
    11'b00101100010: data <= 32'h33cab565;
    11'b00101100011: data <= 32'hbbcb3d56;
    11'b00101100100: data <= 32'hc0b24007;
    11'b00101100101: data <= 32'hc0183afd;
    11'b00101100110: data <= 32'hb1e9b805;
    11'b00101100111: data <= 32'h3c31b8cc;
    11'b00101101000: data <= 32'h382c2e11;
    11'b00101101001: data <= 32'hb2223775;
    11'b00101101010: data <= 32'h39113949;
    11'b00101101011: data <= 32'h401f3d16;
    11'b00101101100: data <= 32'h3f733e8c;
    11'b00101101101: data <= 32'ha6cb3928;
    11'b00101101110: data <= 32'hbd49bc6e;
    11'b00101101111: data <= 32'hb951bef6;
    11'b00101110000: data <= 32'h3998baf5;
    11'b00101110001: data <= 32'h3c65b46f;
    11'b00101110010: data <= 32'h398ebc5f;
    11'b00101110011: data <= 32'h37a3bf7c;
    11'b00101110100: data <= 32'h347cba6d;
    11'b00101110101: data <= 32'hb94a3d05;
    11'b00101110110: data <= 32'hbf4c3f1c;
    11'b00101110111: data <= 32'hbf5e322e;
    11'b00101111000: data <= 32'hba2bbd5f;
    11'b00101111001: data <= 32'hb2d9bc50;
    11'b00101111010: data <= 32'hb9ef3167;
    11'b00101111011: data <= 32'hbabf3a3c;
    11'b00101111100: data <= 32'h38a63a37;
    11'b00101111101: data <= 32'h40213c91;
    11'b00101111110: data <= 32'h3df93ebf;
    11'b00101111111: data <= 32'hb8ed3d5a;
    11'b00110000000: data <= 32'hbe673229;
    11'b00110000001: data <= 32'hb57ab6f0;
    11'b00110000010: data <= 32'h3d70b2b8;
    11'b00110000011: data <= 32'h3e61b5fc;
    11'b00110000100: data <= 32'h3ad7bdcd;
    11'b00110000101: data <= 32'h3931bfc4;
    11'b00110000110: data <= 32'h3b72b884;
    11'b00110000111: data <= 32'h38083d4b;
    11'b00110001000: data <= 32'hb95b3d21;
    11'b00110001001: data <= 32'hbd62b9a1;
    11'b00110001010: data <= 32'hbc75c034;
    11'b00110001011: data <= 32'hbba3bd91;
    11'b00110001100: data <= 32'hbd0f2a0a;
    11'b00110001101: data <= 32'hbbb7359f;
    11'b00110001110: data <= 32'h37c3ae36;
    11'b00110001111: data <= 32'h3e26344c;
    11'b00110010000: data <= 32'h38713dd1;
    11'b00110010001: data <= 32'hbdd83fdf;
    11'b00110010010: data <= 32'hbfb53d1b;
    11'b00110010011: data <= 32'hb46f3734;
    11'b00110010100: data <= 32'h3d333185;
    11'b00110010101: data <= 32'h3c86b303;
    11'b00110010110: data <= 32'h3510bc2e;
    11'b00110010111: data <= 32'h3959bcb0;
    11'b00110011000: data <= 32'h3f2a3142;
    11'b00110011001: data <= 32'h3f503e23;
    11'b00110011010: data <= 32'h36c53bbd;
    11'b00110011011: data <= 32'hbafcbc3f;
    11'b00110011100: data <= 32'hbc38c02e;
    11'b00110011101: data <= 32'hba85bcb4;
    11'b00110011110: data <= 32'hba94b012;
    11'b00110011111: data <= 32'hb80cb8af;
    11'b00110100000: data <= 32'h37dabdfc;
    11'b00110100001: data <= 32'h3bdbbaf0;
    11'b00110100010: data <= 32'hb0f23c3e;
    11'b00110100011: data <= 32'hbf594052;
    11'b00110100100: data <= 32'hbfd63e12;
    11'b00110100101: data <= 32'hb7913691;
    11'b00110100110: data <= 32'h37ca28be;
    11'b00110100111: data <= 32'hb056a0b4;
    11'b00110101000: data <= 32'hb9a4b519;
    11'b00110101001: data <= 32'h3774b41c;
    11'b00110101010: data <= 32'h40a63a1c;
    11'b00110101011: data <= 32'h41053eb6;
    11'b00110101100: data <= 32'h3a503c34;
    11'b00110101101: data <= 32'hb9ebb859;
    11'b00110101110: data <= 32'hb9c5bc95;
    11'b00110101111: data <= 32'ha9bab66c;
    11'b00110110000: data <= 32'h2ff7b0e4;
    11'b00110110001: data <= 32'h2f8ebdbf;
    11'b00110110010: data <= 32'h38a0c128;
    11'b00110110011: data <= 32'h3ab6be4e;
    11'b00110110100: data <= 32'ha7033a34;
    11'b00110110101: data <= 32'hbd423f7a;
    11'b00110110110: data <= 32'hbe023b11;
    11'b00110110111: data <= 32'hb99fb65c;
    11'b00110111000: data <= 32'hb883b736;
    11'b00110111001: data <= 32'hbde32e27;
    11'b00110111010: data <= 32'hbe833026;
    11'b00110111011: data <= 32'h313725b2;
    11'b00110111100: data <= 32'h407e3935;
    11'b00110111101: data <= 32'h40663e0a;
    11'b00110111110: data <= 32'h34553d9e;
    11'b00110111111: data <= 32'hbc023855;
    11'b00111000000: data <= 32'hb61a3376;
    11'b00111000001: data <= 32'h39af386b;
    11'b00111000010: data <= 32'h3a0f2937;
    11'b00111000011: data <= 32'h34f9bebf;
    11'b00111000100: data <= 32'h3890c170;
    11'b00111000101: data <= 32'h3cb5bdcd;
    11'b00111000110: data <= 32'h3b643a57;
    11'b00111000111: data <= 32'hae193d6f;
    11'b00111001000: data <= 32'hb99aacd1;
    11'b00111001001: data <= 32'hb9c9bd11;
    11'b00111001010: data <= 32'hbcb2ba72;
    11'b00111001011: data <= 32'hc0292f4e;
    11'b00111001100: data <= 32'hbfa0a59c;
    11'b00111001101: data <= 32'ha69eb925;
    11'b00111001110: data <= 32'h3ecbb463;
    11'b00111001111: data <= 32'h3ce83bc6;
    11'b00111010000: data <= 32'hb93e3ec3;
    11'b00111010001: data <= 32'hbd7d3de7;
    11'b00111010010: data <= 32'hb2cc3cdb;
    11'b00111010011: data <= 32'h3b1e3c8e;
    11'b00111010100: data <= 32'h37e3355e;
    11'b00111010101: data <= 32'hb432bcfe;
    11'b00111010110: data <= 32'h34cebfc5;
    11'b00111010111: data <= 32'h3ebfb961;
    11'b00111011000: data <= 32'h402a3c2d;
    11'b00111011001: data <= 32'h3c6a3bc1;
    11'b00111011010: data <= 32'h252db918;
    11'b00111011011: data <= 32'hb799bdc8;
    11'b00111011100: data <= 32'hbbe2b89b;
    11'b00111011101: data <= 32'hbea03280;
    11'b00111011110: data <= 32'hbdc2b8eb;
    11'b00111011111: data <= 32'h1e96bf79;
    11'b00111100000: data <= 32'h3c5cbe14;
    11'b00111100001: data <= 32'h358c34c0;
    11'b00111100010: data <= 32'hbcd83e97;
    11'b00111100011: data <= 32'hbda63e99;
    11'b00111100100: data <= 32'hb1a73ce2;
    11'b00111100101: data <= 32'h367c3c2c;
    11'b00111100110: data <= 32'hb8c2385c;
    11'b00111100111: data <= 32'hbd90b7be;
    11'b00111101000: data <= 32'hb297bb1c;
    11'b00111101001: data <= 32'h3fca2e00;
    11'b00111101010: data <= 32'h415b3cde;
    11'b00111101011: data <= 32'h3e2b3adb;
    11'b00111101100: data <= 32'h33e4b6d8;
    11'b00111101101: data <= 32'haea0b976;
    11'b00111101110: data <= 32'hb1d934c3;
    11'b00111101111: data <= 32'hb8d337da;
    11'b00111110000: data <= 32'hb956bcab;
    11'b00111110001: data <= 32'h3076c1b3;
    11'b00111110010: data <= 32'h3a4cc0a6;
    11'b00111110011: data <= 32'h31fab051;
    11'b00111110100: data <= 32'hbb063d19;
    11'b00111110101: data <= 32'hbafc3bd6;
    11'b00111110110: data <= 32'hae1a3570;
    11'b00111110111: data <= 32'hb54a36f9;
    11'b00111111000: data <= 32'hbf4938c8;
    11'b00111111001: data <= 32'hc0dc2dd6;
    11'b00111111010: data <= 32'hb9a5b58c;
    11'b00111111011: data <= 32'h3ef831aa;
    11'b00111111100: data <= 32'h40a73bec;
    11'b00111111101: data <= 32'h3bdf3b4d;
    11'b00111111110: data <= 32'hae2f3559;
    11'b00111111111: data <= 32'h3217389d;
    11'b01000000000: data <= 32'h39613d8a;
    11'b01000000001: data <= 32'h34413b67;
    11'b01000000010: data <= 32'hb462bcfd;
    11'b01000000011: data <= 32'h2ea0c1e3;
    11'b01000000100: data <= 32'h3acfc063;
    11'b01000000101: data <= 32'h3a83ad4e;
    11'b01000000110: data <= 32'h32c13a55;
    11'b01000000111: data <= 32'h2c81abc1;
    11'b01000001000: data <= 32'h3124b9e8;
    11'b01000001001: data <= 32'hb9deaf8d;
    11'b01000001010: data <= 32'hc0c138ec;
    11'b01000001011: data <= 32'hc17c31dd;
    11'b01000001100: data <= 32'hbb4ab98c;
    11'b01000001101: data <= 32'h3cc6b8d2;
    11'b01000001110: data <= 32'h3d233509;
    11'b01000001111: data <= 32'hafe63b2f;
    11'b01000010000: data <= 32'hb9413c1d;
    11'b01000010001: data <= 32'h35613e02;
    11'b01000010010: data <= 32'h3c414016;
    11'b01000010011: data <= 32'h34f93d2c;
    11'b01000010100: data <= 32'hb97cba35;
    11'b01000010101: data <= 32'hb49ec035;
    11'b01000010110: data <= 32'h3c34bd10;
    11'b01000010111: data <= 32'h3ed53571;
    11'b01000011000: data <= 32'h3d653704;
    11'b01000011001: data <= 32'h3b31ba74;
    11'b01000011010: data <= 32'h3853bcdc;
    11'b01000011011: data <= 32'hb798ac2e;
    11'b01000011100: data <= 32'hbf993a6c;
    11'b01000011101: data <= 32'hc053ae9b;
    11'b01000011110: data <= 32'hb9e0be8b;
    11'b01000011111: data <= 32'h3902bf1e;
    11'b01000100000: data <= 32'h33bfb7ef;
    11'b01000100001: data <= 32'hbbb8395c;
    11'b01000100010: data <= 32'hbb1d3c60;
    11'b01000100011: data <= 32'h37173dda;
    11'b01000100100: data <= 32'h3afc3f83;
    11'b01000100101: data <= 32'hb7c03d97;
    11'b01000100110: data <= 32'hbeefa9ec;
    11'b01000100111: data <= 32'hbb93bb47;
    11'b01000101000: data <= 32'h3c54b347;
    11'b01000101001: data <= 32'h405139be;
    11'b01000101010: data <= 32'h3eff3488;
    11'b01000101011: data <= 32'h3c6bbaff;
    11'b01000101100: data <= 32'h3adbba04;
    11'b01000101101: data <= 32'h34ed39b2;
    11'b01000101110: data <= 32'hb9cc3cfc;
    11'b01000101111: data <= 32'hbc8db655;
    11'b01000110000: data <= 32'hb63fc0e3;
    11'b01000110001: data <= 32'h34e5c11a;
    11'b01000110010: data <= 32'hb1a7bba5;
    11'b01000110011: data <= 32'hbb8234b5;
    11'b01000110100: data <= 32'hb77336bc;
    11'b01000110101: data <= 32'h396837aa;
    11'b01000110110: data <= 32'h36ab3c31;
    11'b01000110111: data <= 32'hbe0b3cfa;
    11'b01000111000: data <= 32'hc17d3831;
    11'b01000111001: data <= 32'hbe13b019;
    11'b01000111010: data <= 32'h3a8a316b;
    11'b01000111011: data <= 32'h3f19390f;
    11'b01000111100: data <= 32'h3c6b3277;
    11'b01000111101: data <= 32'h389db673;
    11'b01000111110: data <= 32'h3bb63498;
    11'b01000111111: data <= 32'h3c953f17;
    11'b01001000000: data <= 32'h35d43f2a;
    11'b01001000001: data <= 32'hb6d8b5cf;
    11'b01001000010: data <= 32'hb421c0f3;
    11'b01001000011: data <= 32'h341ac0b4;
    11'b01001000100: data <= 32'h30fcba1b;
    11'b01001000101: data <= 32'hadc8a859;
    11'b01001000110: data <= 32'h3726b8cd;
    11'b01001000111: data <= 32'h3c49ba66;
    11'b01001001000: data <= 32'h318a31cc;
    11'b01001001001: data <= 32'hbfec3c47;
    11'b01001001010: data <= 32'hc203399d;
    11'b01001001011: data <= 32'hbe89b1d7;
    11'b01001001100: data <= 32'h361ab592;
    11'b01001001101: data <= 32'h39f318cb;
    11'b01001001110: data <= 32'hb1ea2799;
    11'b01001001111: data <= 32'hb4922dea;
    11'b01001010000: data <= 32'h3b383c6a;
    11'b01001010001: data <= 32'h3e6340cd;
    11'b01001010010: data <= 32'h398d403e;
    11'b01001010011: data <= 32'hb8732980;
    11'b01001010100: data <= 32'hb8a6be8c;
    11'b01001010101: data <= 32'h34b2bd0a;
    11'b01001010110: data <= 32'h3a8fab5f;
    11'b01001010111: data <= 32'h3b54b1a3;
    11'b01001011000: data <= 32'h3d0ebd8a;
    11'b01001011001: data <= 32'h3ddfbe35;
    11'b01001011010: data <= 32'h36aeac5b;
    11'b01001011011: data <= 32'hbdf63ca2;
    11'b01001011100: data <= 32'hc092388f;
    11'b01001011101: data <= 32'hbcd0bafb;
    11'b01001011110: data <= 32'h247ebd79;
    11'b01001011111: data <= 32'hb52fba77;
    11'b01001100000: data <= 32'hbd2db43a;
    11'b01001100001: data <= 32'hbaaf2fba;
    11'b01001100010: data <= 32'h3b0c3c27;
    11'b01001100011: data <= 32'h3e2e4040;
    11'b01001100100: data <= 32'h31504006;
    11'b01001100101: data <= 32'hbdb138b2;
    11'b01001100110: data <= 32'hbcf5b6c2;
    11'b01001100111: data <= 32'h330928cc;
    11'b01001101000: data <= 32'h3cbd3932;
    11'b01001101001: data <= 32'h3d18b19c;
    11'b01001101010: data <= 32'h3d91be4c;
    11'b01001101011: data <= 32'h3e7dbd77;
    11'b01001101100: data <= 32'h3c2d3804;
    11'b01001101101: data <= 32'hb4cf3e60;
    11'b01001101110: data <= 32'hbc10368b;
    11'b01001101111: data <= 32'hb833be35;
    11'b01001110000: data <= 32'hafe3c02a;
    11'b01001110001: data <= 32'hbac7bce2;
    11'b01001110010: data <= 32'hbe38b846;
    11'b01001110011: data <= 32'hb92db6f6;
    11'b01001110100: data <= 32'h3c592907;
    11'b01001110101: data <= 32'h3cf03c48;
    11'b01001110110: data <= 32'hb9973e21;
    11'b01001110111: data <= 32'hc0b83bb3;
    11'b01001111000: data <= 32'hbf2a3729;
    11'b01001111001: data <= 32'h1c8439d7;
    11'b01001111010: data <= 32'h3afd3aa5;
    11'b01001111011: data <= 32'h38e7b298;
    11'b01001111100: data <= 32'h3954bd05;
    11'b01001111101: data <= 32'h3db1b824;
    11'b01001111110: data <= 32'h3eba3de1;
    11'b01001111111: data <= 32'h3ae74047;
    11'b01010000000: data <= 32'h9c163718;
    11'b01010000001: data <= 32'hae13be74;
    11'b01010000010: data <= 32'haddfbf73;
    11'b01010000011: data <= 32'hb953baea;
    11'b01010000100: data <= 32'hbb62b8bc;
    11'b01010000101: data <= 32'h30d7bd0f;
    11'b01010000110: data <= 32'h3dfcbd36;
    11'b01010000111: data <= 32'h3c25ae53;
    11'b01010001000: data <= 32'hbca23c22;
    11'b01010001001: data <= 32'hc1323c1b;
    11'b01010001010: data <= 32'hbf1d384d;
    11'b01010001011: data <= 32'hb2943749;
    11'b01010001100: data <= 32'h2364357d;
    11'b01010001101: data <= 32'hb9ddb64e;
    11'b01010001110: data <= 32'hb7dcbaba;
    11'b01010001111: data <= 32'h3c163407;
    11'b01010010000: data <= 32'h3ff74026;
    11'b01010010001: data <= 32'h3d5040c2;
    11'b01010010010: data <= 32'h30543962;
    11'b01010010011: data <= 32'hb3a7bb5c;
    11'b01010010100: data <= 32'habbeb9c2;
    11'b01010010101: data <= 32'haf142fdb;
    11'b01010010110: data <= 32'h10deb644;
    11'b01010010111: data <= 32'h3b87bf8e;
    11'b01010011000: data <= 32'h3f5ec05d;
    11'b01010011001: data <= 32'h3ca0b919;
    11'b01010011010: data <= 32'hba463b3c;
    11'b01010011011: data <= 32'hbf563b0b;
    11'b01010011100: data <= 32'hbc5ba662;
    11'b01010011101: data <= 32'hb38eb728;
    11'b01010011110: data <= 32'hbb12b6df;
    11'b01010011111: data <= 32'hbfd9b95c;
    11'b01010100000: data <= 32'hbd65b9ec;
    11'b01010100001: data <= 32'h39f3345c;
    11'b01010100010: data <= 32'h3f973f10;
    11'b01010100011: data <= 32'h3b7f4016;
    11'b01010100100: data <= 32'hb8a33b3d;
    11'b01010100101: data <= 32'hbab92fe8;
    11'b01010100110: data <= 32'hb074398b;
    11'b01010100111: data <= 32'h34723c9c;
    11'b01010101000: data <= 32'h369fae6a;
    11'b01010101001: data <= 32'h3c30c005;
    11'b01010101010: data <= 32'h3f3dc047;
    11'b01010101011: data <= 32'h3e03b40c;
    11'b01010101100: data <= 32'h33b53d04;
    11'b01010101101: data <= 32'hb74639df;
    11'b01010101110: data <= 32'had28b97e;
    11'b01010101111: data <= 32'hab98bcbd;
    11'b01010110000: data <= 32'hbd41baa6;
    11'b01010110001: data <= 32'hc0bdba65;
    11'b01010110010: data <= 32'hbd86bc3c;
    11'b01010110011: data <= 32'h3aa6b894;
    11'b01010110100: data <= 32'h3e6638e6;
    11'b01010110101: data <= 32'h2fc23cf2;
    11'b01010110110: data <= 32'hbe073b8f;
    11'b01010110111: data <= 32'hbd8b3b0c;
    11'b01010111000: data <= 32'hb41f3e28;
    11'b01010111001: data <= 32'h31013e5b;
    11'b01010111010: data <= 32'haf0326f9;
    11'b01010111011: data <= 32'h33a6bec5;
    11'b01010111100: data <= 32'h3d33bd75;
    11'b01010111101: data <= 32'h3f343967;
    11'b01010111110: data <= 32'h3d1b3f2b;
    11'b01010111111: data <= 32'h39ba39ab;
    11'b01011000000: data <= 32'h3921bb21;
    11'b01011000001: data <= 32'h3188bc55;
    11'b01011000010: data <= 32'hbc7cb691;
    11'b01011000011: data <= 32'hbf58b89c;
    11'b01011000100: data <= 32'hb940be3c;
    11'b01011000101: data <= 32'h3ce5bf1d;
    11'b01011000110: data <= 32'h3d7cb9bb;
    11'b01011000111: data <= 32'hb70036a6;
    11'b01011001000: data <= 32'hbf623a22;
    11'b01011001001: data <= 32'hbd513b88;
    11'b01011001010: data <= 32'hb3313d89;
    11'b01011001011: data <= 32'hb6553cdd;
    11'b01011001100: data <= 32'hbd45b010;
    11'b01011001101: data <= 32'hbc4bbd14;
    11'b01011001110: data <= 32'h3878b844;
    11'b01011001111: data <= 32'h3f533d72;
    11'b01011010000: data <= 32'h3ec54005;
    11'b01011010001: data <= 32'h3bf639e5;
    11'b01011010010: data <= 32'h3940b796;
    11'b01011010011: data <= 32'h3446acd0;
    11'b01011010100: data <= 32'hb88b39c8;
    11'b01011010101: data <= 32'hbb18a77a;
    11'b01011010110: data <= 32'h3237bf84;
    11'b01011010111: data <= 32'h3e41c12e;
    11'b01011011000: data <= 32'h3d55bda7;
    11'b01011011001: data <= 32'hb4e92d13;
    11'b01011011010: data <= 32'hbcd93824;
    11'b01011011011: data <= 32'hb80e361f;
    11'b01011011100: data <= 32'h2d7537d7;
    11'b01011011101: data <= 32'hbbd13689;
    11'b01011011110: data <= 32'hc0efb68e;
    11'b01011011111: data <= 32'hc035bc35;
    11'b01011100000: data <= 32'h2737b4dc;
    11'b01011100001: data <= 32'h3e5e3cb8;
    11'b01011100010: data <= 32'h3d323e3f;
    11'b01011100011: data <= 32'h3526392b;
    11'b01011100100: data <= 32'h2b053405;
    11'b01011100101: data <= 32'h31c83d01;
    11'b01011100110: data <= 32'hae5d3fc1;
    11'b01011100111: data <= 32'hb4cf386e;
    11'b01011101000: data <= 32'h36d2bf3f;
    11'b01011101001: data <= 32'h3dcac112;
    11'b01011101010: data <= 32'h3d8abc67;
    11'b01011101011: data <= 32'h36833636;
    11'b01011101100: data <= 32'h2cce35e0;
    11'b01011101101: data <= 32'h398eb54d;
    11'b01011101110: data <= 32'h38aeb626;
    11'b01011101111: data <= 32'hbcbcaf44;
    11'b01011110000: data <= 32'hc1b6b7c8;
    11'b01011110001: data <= 32'hc07bbc73;
    11'b01011110010: data <= 32'h26febad0;
    11'b01011110011: data <= 32'h3d123005;
    11'b01011110100: data <= 32'h372f387f;
    11'b01011110101: data <= 32'hb9aa3578;
    11'b01011110110: data <= 32'hb8cc3a0d;
    11'b01011110111: data <= 32'h2d984024;
    11'b01011111000: data <= 32'h9c524106;
    11'b01011111001: data <= 32'hb8603a8f;
    11'b01011111010: data <= 32'hb462bdc0;
    11'b01011111011: data <= 32'h3a13bef2;
    11'b01011111100: data <= 32'h3d52aeae;
    11'b01011111101: data <= 32'h3cac3c11;
    11'b01011111110: data <= 32'h3cdc3560;
    11'b01011111111: data <= 32'h3e57b9b3;
    11'b01100000000: data <= 32'h3c08b849;
    11'b01100000001: data <= 32'hbb323215;
    11'b01100000010: data <= 32'hc09baed9;
    11'b01100000011: data <= 32'hbdeebd12;
    11'b01100000100: data <= 32'h37c4bf14;
    11'b01100000101: data <= 32'h3c2bbcaa;
    11'b01100000110: data <= 32'hb409b743;
    11'b01100000111: data <= 32'hbd1aad08;
    11'b01100001000: data <= 32'hb9573981;
    11'b01100001001: data <= 32'h33e93f9f;
    11'b01100001010: data <= 32'hb3644049;
    11'b01100001011: data <= 32'hbdda3914;
    11'b01100001100: data <= 32'hbe2bbc11;
    11'b01100001101: data <= 32'hb23bba55;
    11'b01100001110: data <= 32'h3c4c3a4b;
    11'b01100001111: data <= 32'h3dad3d75;
    11'b01100010000: data <= 32'h3df4344c;
    11'b01100010001: data <= 32'h3e99b8c0;
    11'b01100010010: data <= 32'h3c7731de;
    11'b01100010011: data <= 32'hb56d3d13;
    11'b01100010100: data <= 32'hbd0e3944;
    11'b01100010101: data <= 32'hb73ebd15;
    11'b01100010110: data <= 32'h3bacc0c5;
    11'b01100010111: data <= 32'h3b81bf72;
    11'b01100011000: data <= 32'hb63ebb17;
    11'b01100011001: data <= 32'hbb63b652;
    11'b01100011010: data <= 32'h2d942e91;
    11'b01100011011: data <= 32'h3a283b89;
    11'b01100011100: data <= 32'hb7a83cc0;
    11'b01100011101: data <= 32'hc0c9331d;
    11'b01100011110: data <= 32'hc126ba17;
    11'b01100011111: data <= 32'hbaeab52d;
    11'b01100100000: data <= 32'h39b13b0b;
    11'b01100100001: data <= 32'h3bc73c00;
    11'b01100100010: data <= 32'h3a1ea522;
    11'b01100100011: data <= 32'h3b80b2a0;
    11'b01100100100: data <= 32'h3b533d18;
    11'b01100100101: data <= 32'h30c140f9;
    11'b01100100110: data <= 32'hb7823daa;
    11'b01100100111: data <= 32'h2a15bc1a;
    11'b01100101000: data <= 32'h3b92c07e;
    11'b01100101001: data <= 32'h3a86be10;
    11'b01100101010: data <= 32'ha19db815;
    11'b01100101011: data <= 32'h2f6db75b;
    11'b01100101100: data <= 32'h3d2ab8f8;
    11'b01100101101: data <= 32'h3de5af2b;
    11'b01100101110: data <= 32'hb75e368b;
    11'b01100101111: data <= 32'hc15625b4;
    11'b01100110000: data <= 32'hc162b96c;
    11'b01100110001: data <= 32'hbac6b862;
    11'b01100110010: data <= 32'h36ea2d5a;
    11'b01100110011: data <= 32'h2f081cd3;
    11'b01100110100: data <= 32'hb6b3b863;
    11'b01100110101: data <= 32'h29962871;
    11'b01100110110: data <= 32'h39783fd4;
    11'b01100110111: data <= 32'h35ac421e;
    11'b01100111000: data <= 32'hb68e3edd;
    11'b01100111001: data <= 32'hb62ab932;
    11'b01100111010: data <= 32'h346fbdb2;
    11'b01100111011: data <= 32'h383db63a;
    11'b01100111100: data <= 32'h37553553;
    11'b01100111101: data <= 32'h3c65b590;
    11'b01100111110: data <= 32'h4065bc56;
    11'b01100111111: data <= 32'h3feeb862;
    11'b01101000000: data <= 32'hafda36fe;
    11'b01101000001: data <= 32'hc02835be;
    11'b01101000010: data <= 32'hbf4fb8dc;
    11'b01101000011: data <= 32'hb28fbc9e;
    11'b01101000100: data <= 32'h357fbc21;
    11'b01101000101: data <= 32'hb937bc2b;
    11'b01101000110: data <= 32'hbcfebc6a;
    11'b01101000111: data <= 32'hb4dfb06a;
    11'b01101001000: data <= 32'h3a333ef2;
    11'b01101001001: data <= 32'h355a4139;
    11'b01101001010: data <= 32'hbc053d8b;
    11'b01101001011: data <= 32'hbdd6b590;
    11'b01101001100: data <= 32'hb9b7b6e6;
    11'b01101001101: data <= 32'h2e3239f5;
    11'b01101001110: data <= 32'h386f3bb4;
    11'b01101001111: data <= 32'h3d36b522;
    11'b01101010000: data <= 32'h406dbc97;
    11'b01101010001: data <= 32'h3ffbb0c4;
    11'b01101010010: data <= 32'h35883d37;
    11'b01101010011: data <= 32'hbbfa3ca2;
    11'b01101010100: data <= 32'hb897b675;
    11'b01101010101: data <= 32'h3861be49;
    11'b01101010110: data <= 32'h35afbe90;
    11'b01101010111: data <= 32'hbb92bdd4;
    11'b01101011000: data <= 32'hbcdabd86;
    11'b01101011001: data <= 32'h3312b95b;
    11'b01101011010: data <= 32'h3d4639e1;
    11'b01101011011: data <= 32'h34f43dd2;
    11'b01101011100: data <= 32'hbece39a4;
    11'b01101011101: data <= 32'hc0c6b324;
    11'b01101011110: data <= 32'hbd943173;
    11'b01101011111: data <= 32'hb4983c99;
    11'b01101100000: data <= 32'h2f623ac4;
    11'b01101100001: data <= 32'h384fb8e4;
    11'b01101100010: data <= 32'h3d52bbe6;
    11'b01101100011: data <= 32'h3e303975;
    11'b01101100100: data <= 32'h399040ce;
    11'b01101100101: data <= 32'hadbf3fcd;
    11'b01101100110: data <= 32'h336cad49;
    11'b01101100111: data <= 32'h3a6abd91;
    11'b01101101000: data <= 32'h3418bd00;
    11'b01101101001: data <= 32'hba50bb8e;
    11'b01101101010: data <= 32'hb733bcf0;
    11'b01101101011: data <= 32'h3d2abd0b;
    11'b01101101100: data <= 32'h4025b6a0;
    11'b01101101101: data <= 32'h37383611;
    11'b01101101110: data <= 32'hbf913304;
    11'b01101101111: data <= 32'hc0e8b227;
    11'b01101110000: data <= 32'hbd1c3103;
    11'b01101110001: data <= 32'hb66c3929;
    11'b01101110010: data <= 32'hb90f1907;
    11'b01101110011: data <= 32'hb9d1bccb;
    11'b01101110100: data <= 32'h30e7bb41;
    11'b01101110101: data <= 32'h3c123cf7;
    11'b01101110110: data <= 32'h3a8e41d7;
    11'b01101110111: data <= 32'h31454060;
    11'b01101111000: data <= 32'h2eb731d4;
    11'b01101111001: data <= 32'h34f5b93e;
    11'b01101111010: data <= 32'had6caa3c;
    11'b01101111011: data <= 32'hb8153132;
    11'b01101111100: data <= 32'h35fbba9a;
    11'b01101111101: data <= 32'h4047be7a;
    11'b01101111110: data <= 32'h411ebc1b;
    11'b01101111111: data <= 32'h39de2dce;
    11'b01110000000: data <= 32'hbd6a3598;
    11'b01110000001: data <= 32'hbe15ad3f;
    11'b01110000010: data <= 32'hb65fb3ba;
    11'b01110000011: data <= 32'hb297b47d;
    11'b01110000100: data <= 32'hbd1cbbd6;
    11'b01110000101: data <= 32'hbedfbf12;
    11'b01110000110: data <= 32'hb826bc52;
    11'b01110000111: data <= 32'h3afa3c26;
    11'b01110001000: data <= 32'h3a8640d1;
    11'b01110001001: data <= 32'hb2e03e9d;
    11'b01110001010: data <= 32'hb9ff332a;
    11'b01110001011: data <= 32'hb8d63306;
    11'b01110001100: data <= 32'hb87f3cef;
    11'b01110001101: data <= 32'hb7803c7a;
    11'b01110001110: data <= 32'h3879b846;
    11'b01110001111: data <= 32'h4034beae;
    11'b01110010000: data <= 32'h40d0babf;
    11'b01110010001: data <= 32'h3bd239b2;
    11'b01110010010: data <= 32'hb6203c35;
    11'b01110010011: data <= 32'hb02131e3;
    11'b01110010100: data <= 32'h3972b873;
    11'b01110010101: data <= 32'h2dd4bab0;
    11'b01110010110: data <= 32'hbe22bd67;
    11'b01110010111: data <= 32'hbf92bfb6;
    11'b01110011000: data <= 32'hb431bdbb;
    11'b01110011001: data <= 32'h3d2c303b;
    11'b01110011010: data <= 32'h3ada3c81;
    11'b01110011011: data <= 32'hba2f393b;
    11'b01110011100: data <= 32'hbe5e2a6b;
    11'b01110011101: data <= 32'hbcff3a15;
    11'b01110011110: data <= 32'hbb043f61;
    11'b01110011111: data <= 32'hba3f3d2d;
    11'b01110100000: data <= 32'hb018b95e;
    11'b01110100001: data <= 32'h3c6cbe46;
    11'b01110100010: data <= 32'h3ea2b19d;
    11'b01110100011: data <= 32'h3c1a3ec7;
    11'b01110100100: data <= 32'h372b3f3e;
    11'b01110100101: data <= 32'h3b0b37b1;
    11'b01110100110: data <= 32'h3d00b72e;
    11'b01110100111: data <= 32'h31beb7f7;
    11'b01110101000: data <= 32'hbdafb9f4;
    11'b01110101001: data <= 32'hbd3fbe0c;
    11'b01110101010: data <= 32'h394abef0;
    11'b01110101011: data <= 32'h4005bb71;
    11'b01110101100: data <= 32'h3c09b0c3;
    11'b01110101101: data <= 32'hbbddb165;
    11'b01110101110: data <= 32'hbebeb08b;
    11'b01110101111: data <= 32'hbc3a3a2f;
    11'b01110110000: data <= 32'hba1c3e25;
    11'b01110110001: data <= 32'hbd0f3907;
    11'b01110110010: data <= 32'hbd38bcd5;
    11'b01110110011: data <= 32'hb433be1b;
    11'b01110110100: data <= 32'h3a3d35bd;
    11'b01110110101: data <= 32'h3b28406d;
    11'b01110110110: data <= 32'h39a93ff8;
    11'b01110110111: data <= 32'h3bb23884;
    11'b01110111000: data <= 32'h3bc32bcc;
    11'b01110111001: data <= 32'hade838f4;
    11'b01110111010: data <= 32'hbcc93855;
    11'b01110111011: data <= 32'hb869ba00;
    11'b01110111100: data <= 32'h3df5bf40;
    11'b01110111101: data <= 32'h40eabe1c;
    11'b01110111110: data <= 32'h3ca4b940;
    11'b01110111111: data <= 32'hb907b49b;
    11'b01111000000: data <= 32'hba9bb02d;
    11'b01111000001: data <= 32'ha31e36f8;
    11'b01111000010: data <= 32'hb33c39aa;
    11'b01111000011: data <= 32'hbe7ab4f5;
    11'b01111000100: data <= 32'hc086bf07;
    11'b01111000101: data <= 32'hbca4be76;
    11'b01111000110: data <= 32'h358b34b8;
    11'b01111000111: data <= 32'h3a093f10;
    11'b01111001000: data <= 32'h362a3d41;
    11'b01111001001: data <= 32'h338f3495;
    11'b01111001010: data <= 32'h3018392d;
    11'b01111001011: data <= 32'hb8733f6f;
    11'b01111001100: data <= 32'hbc753eeb;
    11'b01111001101: data <= 32'hb44fb077;
    11'b01111001110: data <= 32'h3e05bec1;
    11'b01111001111: data <= 32'h4060bd8f;
    11'b01111010000: data <= 32'h3c77b21c;
    11'b01111010001: data <= 32'h2c3e34ea;
    11'b01111010010: data <= 32'h38262fa2;
    11'b01111010011: data <= 32'h3d312f79;
    11'b01111010100: data <= 32'h36a32e50;
    11'b01111010101: data <= 32'hbea8b9cf;
    11'b01111010110: data <= 32'hc0f1bf50;
    11'b01111010111: data <= 32'hbc56bee2;
    11'b01111011000: data <= 32'h38f6b5b4;
    11'b01111011001: data <= 32'h3a1c3841;
    11'b01111011010: data <= 32'hb0d82d58;
    11'b01111011011: data <= 32'hb8f5b3e7;
    11'b01111011100: data <= 32'hb8643b9b;
    11'b01111011101: data <= 32'hba8340fc;
    11'b01111011110: data <= 32'hbce94037;
    11'b01111011111: data <= 32'hb9d7ad8e;
    11'b01111100000: data <= 32'h387ebe1e;
    11'b01111100001: data <= 32'h3ce1ba10;
    11'b01111100010: data <= 32'h3a673a24;
    11'b01111100011: data <= 32'h391f3c52;
    11'b01111100100: data <= 32'h3e2b3626;
    11'b01111100101: data <= 32'h40302cde;
    11'b01111100110: data <= 32'h39e533ca;
    11'b01111100111: data <= 32'hbddbb197;
    11'b01111101000: data <= 32'hbfbabcdc;
    11'b01111101001: data <= 32'hb2f8beab;
    11'b01111101010: data <= 32'h3d50bc9b;
    11'b01111101011: data <= 32'h3b35ba01;
    11'b01111101100: data <= 32'hb76cbbe3;
    11'b01111101101: data <= 32'hbaf8b9ba;
    11'b01111101110: data <= 32'hb6a53aba;
    11'b01111101111: data <= 32'hb8464075;
    11'b01111110000: data <= 32'hbd863e21;
    11'b01111110001: data <= 32'hbe8fb8b0;
    11'b01111110010: data <= 32'hba75bde8;
    11'b01111110011: data <= 32'h2d12b111;
    11'b01111110100: data <= 32'h35a53da5;
    11'b01111110101: data <= 32'h39f33d4a;
    11'b01111110110: data <= 32'h3eaf3562;
    11'b01111110111: data <= 32'h3fc334a3;
    11'b01111111000: data <= 32'h38523c6a;
    11'b01111111001: data <= 32'hbce63c6a;
    11'b01111111010: data <= 32'hbc8bb1fd;
    11'b01111111011: data <= 32'h399dbd9a;
    11'b01111111100: data <= 32'h3f58be3f;
    11'b01111111101: data <= 32'h3ba1bd3a;
    11'b01111111110: data <= 32'hb5d8bd15;
    11'b01111111111: data <= 32'hb408ba99;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    