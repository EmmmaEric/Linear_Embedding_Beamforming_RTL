
    module interp_rom_3(
    CLK, rst,
    Addr, CEB, Q
    );

    input CLK, rst;
    input [9:0] Addr;
    input CEB;		
    output [20:0] Q;

    (*rom_style = "block" *) reg [20:0] data;

    always @(posedge CLK) begin
    if (rst) begin
        data <= 20'd0;
    end else begin
    if (CEB)
    case(Addr)
            10'b00000000: data <= 20'b10010100010001000100;
        10'b00000001: data <= 20'b10011101011001010000;
        10'b00000010: data <= 20'b10010011101001100000;
        10'b00000011: data <= 20'b10010100100000111010;
        10'b00000100: data <= 20'b00001111010001001110;
        10'b00000101: data <= 20'b00010001000000101111;
        10'b00000110: data <= 20'b00010101010000011100;
        10'b00000111: data <= 20'b10001011111001101110;
        10'b00001000: data <= 20'b10010010001001010110;
        10'b00001001: data <= 20'b00010110011001101000;
        10'b00001010: data <= 20'b00001111101000100001;
        10'b00001011: data <= 20'b10001001001001010010;
        10'b00001100: data <= 20'b10011000011000010110;
        10'b00001101: data <= 20'b10010111110001000010;
        10'b00001110: data <= 20'b10010100001001000110;
        10'b00001111: data <= 20'b10001010100000111011;
        10'b00010000: data <= 20'b00010011101001001100;
        10'b00010001: data <= 20'b10010110111001010000;
        10'b00010010: data <= 20'b10010100100001100000;
        10'b00010011: data <= 20'b00001000110001001100;
        10'b00010100: data <= 20'b00010101000001010010;
        10'b00010101: data <= 20'b00011000011001001101;
        10'b00010110: data <= 20'b10010111001001000101;
        10'b00010111: data <= 20'b10001001000001000011;
        10'b00011000: data <= 20'b00000011001000010001;
        10'b00011001: data <= 20'b10000100111001110000;
        10'b00011010: data <= 20'b10011001101001111011;
        10'b00011011: data <= 20'b10010101100001001110;
        10'b00011100: data <= 20'b00010000010001000111;
        10'b00011101: data <= 20'b00011000101001100101;
        10'b00011110: data <= 20'b00001111000001010010;
        10'b00011111: data <= 20'b00010111001001011111;
        10'b00100000: data <= 20'b00001000100001001101;
        10'b00100001: data <= 20'b00010010000001101011;
        10'b00100010: data <= 20'b00010100001001010000;
        10'b00100011: data <= 20'b10001011000001010001;
        10'b00100100: data <= 20'b00001010110001001011;
        10'b00100101: data <= 20'b00010001110001000000;
        10'b00100110: data <= 20'b10011001111001100010;
        10'b00100111: data <= 20'b10010110001000101000;
        10'b00101000: data <= 20'b00010110101000000101;
        10'b00101001: data <= 20'b00001000111001011111;
        10'b00101010: data <= 20'b00001100000001011101;
        10'b00101011: data <= 20'b00010011001001011011;
        10'b00101100: data <= 20'b10001100000001001111;
        10'b00101101: data <= 20'b00010101001001111100;
        10'b00101110: data <= 20'b10001100111001001000;
        10'b00101111: data <= 20'b00100001010010000111;
        10'b00110000: data <= 20'b00001001011000100100;
        10'b00110001: data <= 20'b10001111001000000010;
        10'b00110010: data <= 20'b10000111110001000111;
        10'b00110011: data <= 20'b10011001001001011100;
        10'b00110100: data <= 20'b00011001011001110101;
        10'b00110101: data <= 20'b10000110000000001000;
        10'b00110110: data <= 20'b00000110110001010101;
        10'b00110111: data <= 20'b10011000101001100000;
        10'b00111000: data <= 20'b00001000111001010011;
        10'b00111001: data <= 20'b00010101101001011111;
        10'b00111010: data <= 20'b10001001011001011001;
        10'b00111011: data <= 20'b10010110101000111000;
        10'b00111100: data <= 20'b10010000100000110001;
        10'b00111101: data <= 20'b10011001100001011010;
        10'b00111110: data <= 20'b00011000001001001101;
        10'b00111111: data <= 20'b10010100001001001000;
        10'b01000000: data <= 20'b10011000001001000010;
        10'b01000001: data <= 20'b10010001010001001010;
        10'b01000010: data <= 20'b00010100000001010100;
        10'b01000011: data <= 20'b00010111010001010010;
        10'b01000100: data <= 20'b10010000011001010101;
        10'b01000101: data <= 20'b10010100111000001111;
        10'b01000110: data <= 20'b10010011010001000000;
        10'b01000111: data <= 20'b10001100101001000110;
        10'b01001000: data <= 20'b10001011011001001110;
        10'b01001001: data <= 20'b00010000111001011010;
        10'b01001010: data <= 20'b10010010100000010011;
        10'b01001011: data <= 20'b00001101010001100001;
        10'b01001100: data <= 20'b00011011101010000001;
        10'b01001101: data <= 20'b00011000110001110101;
        10'b01001110: data <= 20'b00010010010001001010;
        10'b01001111: data <= 20'b00010101111001000001;
        10'b01010000: data <= 20'b00010101100000111110;
        10'b01010001: data <= 20'b00001011101001000110;
        10'b01010010: data <= 20'b00010101011000111111;
        10'b01010011: data <= 20'b10010001100001000001;
        10'b01010100: data <= 20'b10001000001001100010;
        10'b01010101: data <= 20'b10010010001001011010;
        10'b01010110: data <= 20'b00011001010000110000;
        10'b01010111: data <= 20'b00010110000000001101;
        10'b01011000: data <= 20'b00010010010000100110;
        10'b01011001: data <= 20'b10011010111001100010;
        10'b01011010: data <= 20'b10010100101000111001;
        10'b01011011: data <= 20'b00010100011001000101;
        10'b01011100: data <= 20'b10010000000000000111;
        10'b01011101: data <= 20'b00000110110001000111;
        10'b01011110: data <= 20'b10010101011000001100;
        10'b01011111: data <= 20'b00010111111001010011;
        10'b01100000: data <= 20'b10010001010000011101;
        10'b01100001: data <= 20'b00001110001000000100;
        10'b01100010: data <= 20'b00010010101001000100;
        10'b01100011: data <= 20'b10011000010000111100;
        10'b01100100: data <= 20'b10010101011001100001;
        10'b01100101: data <= 20'b00001110101000110100;
        10'b01100110: data <= 20'b10100000110001110100;
        10'b01100111: data <= 20'b10011010100010000001;
        10'b01101000: data <= 20'b00011100011001111110;
        10'b01101001: data <= 20'b00010010111000110111;
        10'b01101010: data <= 20'b00001110100000100011;
        10'b01101011: data <= 20'b10001000001001101010;
        10'b01101100: data <= 20'b10010101110001000100;
        10'b01101101: data <= 20'b10010011001001001101;
        10'b01101110: data <= 20'b00001100101001000111;
        10'b01101111: data <= 20'b10010000100000010001;
        10'b01110000: data <= 20'b00001101001000110011;
        10'b01110001: data <= 20'b10001101111001010111;
        10'b01110010: data <= 20'b10010100110000001011;
        10'b01110011: data <= 20'b10010111011000110101;
        10'b01110100: data <= 20'b00011001010001100111;
        10'b01110101: data <= 20'b00000010000001110010;
        10'b01110110: data <= 20'b00000011000001010011;
        10'b01110111: data <= 20'b00010100111001000111;
        10'b01111000: data <= 20'b10011001100001110001;
        10'b01111001: data <= 20'b00001110001001001110;
        10'b01111010: data <= 20'b10011000010001100111;
        10'b01111011: data <= 20'b00010001111000100101;
        10'b01111100: data <= 20'b10010000100000011000;
        10'b01111101: data <= 20'b10011000010001100011;
        10'b01111110: data <= 20'b00001100001000110101;
        10'b01111111: data <= 20'b10010011011001100110;
        10'b10000000: data <= 20'b10001111111000111011;
        10'b10000001: data <= 20'b10010010110001000000;
        10'b10000010: data <= 20'b00001011110001001001;
        10'b10000011: data <= 20'b10010111010001011001;
        10'b10000100: data <= 20'b00100011010001101011;
        10'b10000101: data <= 20'b10010110100001000100;
        10'b10000110: data <= 20'b00010011100001011000;
        10'b10000111: data <= 20'b00010000001001010001;
        10'b10001000: data <= 20'b00010010010000110111;
        10'b10001001: data <= 20'b00010001000000111110;
        10'b10001010: data <= 20'b10010100011000110100;
        10'b10001011: data <= 20'b10010110011001001010;
        10'b10001100: data <= 20'b10100001011001110110;
        10'b10001101: data <= 20'b00010110001001001010;
        10'b10001110: data <= 20'b00010001001001100000;
        10'b10001111: data <= 20'b10000000101000110100;
        10'b10010000: data <= 20'b10001000111000100101;
        10'b10010001: data <= 20'b00010001110000110100;
        10'b10010010: data <= 20'b10010010011001000010;
        10'b10010011: data <= 20'b00010101101001111001;
        10'b10010100: data <= 20'b10011010110001000001;
        10'b10010101: data <= 20'b00010011011000111011;
        10'b10010110: data <= 20'b00001100101000010110;
        10'b10010111: data <= 20'b10001101101000110100;
        10'b10011000: data <= 20'b10000010000000101010;
        10'b10011001: data <= 20'b00010111000000111000;
        10'b10011010: data <= 20'b00010101101000111010;
        10'b10011011: data <= 20'b10010001001000111010;
        10'b10011100: data <= 20'b10001111100000100110;
        10'b10011101: data <= 20'b00000101100000001111;
        10'b10011110: data <= 20'b00010110001001110000;
        10'b10011111: data <= 20'b10010100100001001001;
        10'b10100000: data <= 20'b00001000001000111101;
        10'b10100001: data <= 20'b10010000010001001111;
        10'b10100010: data <= 20'b00000110110000001011;
        10'b10100011: data <= 20'b10001000101000110010;
        10'b10100100: data <= 20'b10010001111001000010;
        10'b10100101: data <= 20'b10010101010001010011;
        10'b10100110: data <= 20'b10010111101001101011;
        10'b10100111: data <= 20'b00010101100001000001;
        10'b10101000: data <= 20'b10000101001001001000;
        10'b10101001: data <= 20'b00010101011000111011;
        10'b10101010: data <= 20'b10001011111001000000;
        10'b10101011: data <= 20'b00011000001001011000;
        10'b10101100: data <= 20'b10010100001001000001;
        10'b10101101: data <= 20'b00001101111001001000;
        10'b10101110: data <= 20'b10010100111001010010;
        10'b10101111: data <= 20'b00010011111000110101;
        10'b10110000: data <= 20'b00100001011001000110;
        10'b10110001: data <= 20'b00011010010001011001;
        10'b10110010: data <= 20'b10011000100001010010;
        10'b10110011: data <= 20'b00011000001000000110;
        10'b10110100: data <= 20'b00010111100001011011;
        10'b10110101: data <= 20'b10010100010001100111;
        10'b10110110: data <= 20'b00010100111000110101;
        10'b10110111: data <= 20'b00000101101001000011;
        10'b10111000: data <= 20'b10010001000001101100;
        10'b10111001: data <= 20'b10010001010001001001;
        10'b10111010: data <= 20'b10011010011010010100;
        10'b10111011: data <= 20'b00010111100001010010;
        10'b10111100: data <= 20'b10010100000001000100;
        10'b10111101: data <= 20'b00000010100001010001;
        10'b10111110: data <= 20'b00010110011000101011;
        10'b10111111: data <= 20'b10011101010001010000;
        10'b11000000: data <= 20'b00010010101001010100;
        10'b11000001: data <= 20'b00010110110001011111;
        10'b11000010: data <= 20'b10000010100001100100;
        10'b11000011: data <= 20'b00001101100000001010;
        10'b11000100: data <= 20'b00010000001001010101;
        10'b11000101: data <= 20'b00001101001000100010;
        10'b11000110: data <= 20'b10001110001001000000;
        10'b11000111: data <= 20'b10010000010001011010;
        10'b11001000: data <= 20'b10010100001001100111;
        10'b11001001: data <= 20'b00011100001000100010;
        10'b11001010: data <= 20'b10001001010001010101;
        10'b11001011: data <= 20'b00010101111000111100;
        10'b11001100: data <= 20'b10010011011001000110;
        10'b11001101: data <= 20'b00010001011001011000;
        10'b11001110: data <= 20'b10010010010001010010;
        10'b11001111: data <= 20'b10001110000001010110;
        10'b11010000: data <= 20'b10010110101000011111;
        10'b11010001: data <= 20'b00010111010010000100;
        10'b11010010: data <= 20'b00010101111000111101;
        10'b11010011: data <= 20'b00011000010001101010;
        10'b11010100: data <= 20'b10001110110001010100;
        10'b11010101: data <= 20'b00010011011000111011;
        10'b11010110: data <= 20'b00000100001001001101;
        10'b11010111: data <= 20'b00001000110000111111;
        10'b11011000: data <= 20'b00001111101000111101;
        10'b11011001: data <= 20'b00001011100000010000;
        10'b11011010: data <= 20'b10010010001001010110;
        10'b11011011: data <= 20'b10000101111001011111;
        10'b11011100: data <= 20'b10010111100001100011;
        10'b11011101: data <= 20'b00010111010000101111;
        10'b11011110: data <= 20'b00010000101001011101;
        10'b11011111: data <= 20'b00010100110001000010;
        10'b11100000: data <= 20'b00010100111000111010;
        10'b11100001: data <= 20'b00010011010001000100;
        10'b11100010: data <= 20'b10011101000001001001;
        10'b11100011: data <= 20'b10011100011000111001;
        10'b11100100: data <= 20'b00010000100001010111;
        10'b11100101: data <= 20'b00001101000001010011;
        10'b11100110: data <= 20'b00010101001001100100;
        10'b11100111: data <= 20'b10011000000001101010;
        10'b11101000: data <= 20'b00010000001000011010;
        10'b11101001: data <= 20'b10000011101000110001;
        10'b11101010: data <= 20'b10001110000001000001;
        10'b11101011: data <= 20'b00000010100000010001;
        10'b11101100: data <= 20'b10001111011000001010;
        10'b11101101: data <= 20'b10000001111000011111;
        10'b11101110: data <= 20'b00011010001010000011;
        10'b11101111: data <= 20'b10011001111001100011;
        10'b11110000: data <= 20'b10010000111001001010;
        10'b11110001: data <= 20'b10010101100000100101;
        10'b11110010: data <= 20'b00011000011001000111;
        10'b11110011: data <= 20'b10010100111000100010;
        10'b11110100: data <= 20'b10010101110001001110;
        10'b11110101: data <= 20'b00010001000000101001;
        10'b11110110: data <= 20'b10010110001000100100;
        10'b11110111: data <= 20'b00010101000001000000;
        10'b11111000: data <= 20'b00100100111001111110;
        10'b11111001: data <= 20'b00010001100001011010;
        10'b11111010: data <= 20'b00010010001001011111;
        10'b11111011: data <= 20'b00010101100000110100;
        10'b11111100: data <= 20'b10001110100001010001;
        10'b11111101: data <= 20'b00010100101000011010;
        10'b11111110: data <= 20'b10001010111001010011;
        10'b11111111: data <= 20'b10010011110001000000;
        10'b100000000: data <= 20'b10010001010001011010;
        10'b100000001: data <= 20'b10001101000000111000;
        10'b100000010: data <= 20'b10001101101001010110;
        10'b100000011: data <= 20'b10010011101000110011;
        10'b100000100: data <= 20'b10001010100001011000;
        10'b100000101: data <= 20'b10001111110000100010;
        10'b100000110: data <= 20'b00001110100000100010;
        10'b100000111: data <= 20'b00010111010001101010;
        10'b100001000: data <= 20'b10010010011001010000;
        10'b100001001: data <= 20'b10010100101001000111;
        10'b100001010: data <= 20'b00010010001000010100;
        10'b100001011: data <= 20'b10011000000001011111;
        10'b100001100: data <= 20'b00010000101001011011;
        10'b100001101: data <= 20'b00010111101001000010;
        10'b100001110: data <= 20'b00010011001000111010;
        10'b100001111: data <= 20'b00011010000001000001;
        10'b100010000: data <= 20'b00011000111001011010;
        10'b100010001: data <= 20'b10011100001001100001;
        10'b100010010: data <= 20'b00010000000000111000;
        10'b100010011: data <= 20'b00010111011001110000;
        10'b100010100: data <= 20'b10100000100001111101;
        10'b100010101: data <= 20'b10010110000001100000;
        10'b100010110: data <= 20'b00001110100001001110;
        10'b100010111: data <= 20'b00010111110001010001;
        10'b100011000: data <= 20'b00010111100000100000;
        10'b100011001: data <= 20'b00011010110001000000;
        10'b100011010: data <= 20'b00010010011000100100;
        10'b100011011: data <= 20'b10010001101001010101;
        10'b100011100: data <= 20'b10010100101000110101;
        10'b100011101: data <= 20'b10010001011000110010;
        10'b100011110: data <= 20'b10010010110000101110;
        10'b100011111: data <= 20'b00010011101001000001;
        10'b100100000: data <= 20'b00001001001001100000;
        10'b100100001: data <= 20'b10011000100000111101;
        10'b100100010: data <= 20'b00011110101001011100;
        10'b100100011: data <= 20'b00010110111001010001;
        10'b100100100: data <= 20'b00010111101001001110;
        10'b100100101: data <= 20'b10100000100010000011;
        10'b100100110: data <= 20'b00001110011000110111;
        10'b100100111: data <= 20'b00001011011001000101;
        10'b100101000: data <= 20'b10010010011001100011;
        10'b100101001: data <= 20'b10011000000001100101;
        10'b100101010: data <= 20'b00010111011000111001;
        10'b100101011: data <= 20'b10010110011001001011;
        10'b100101100: data <= 20'b00010101111001010000;
        10'b100101101: data <= 20'b00001110011001010000;
        10'b100101110: data <= 20'b10010010011000101111;
        10'b100101111: data <= 20'b10001100101001000010;
        10'b100110000: data <= 20'b10010001011000111010;
        10'b100110001: data <= 20'b00010001000001000001;
        10'b100110010: data <= 20'b00010001101001110001;
        10'b100110011: data <= 20'b00011110011001101000;
        10'b100110100: data <= 20'b10001001110001000010;
        10'b100110101: data <= 20'b10000101011001001100;
        10'b100110110: data <= 20'b10010111011001110101;
        10'b100110111: data <= 20'b10010100100000000101;
        10'b100111000: data <= 20'b00010101100001010101;
        10'b100111001: data <= 20'b00011000000001000001;
        10'b100111010: data <= 20'b00011000101001101001;
        10'b100111011: data <= 20'b00011100010001010101;
        10'b100111100: data <= 20'b10010000000001010101;
        10'b100111101: data <= 20'b00010010010001001000;
        10'b100111110: data <= 20'b00000001000001011000;
        10'b100111111: data <= 20'b00010001000001010010;
        10'b101000000: data <= 20'b10010000001001000101;
        10'b101000001: data <= 20'b10010110011001100001;
        10'b101000010: data <= 20'b10010001001001010010;
        10'b101000011: data <= 20'b10011000011000110010;
        10'b101000100: data <= 20'b00011010110001101000;
        10'b101000101: data <= 20'b10011000101001101000;
        10'b101000110: data <= 20'b00010001111001010011;
        10'b101000111: data <= 20'b00010001111001010111;
        10'b101001000: data <= 20'b00010110010001000100;
        10'b101001001: data <= 20'b00011010010001100010;
        10'b101001010: data <= 20'b00011000101001010101;
        10'b101001011: data <= 20'b00001011101001001000;
        10'b101001100: data <= 20'b10010000100001000011;
        10'b101001101: data <= 20'b10011110001010000000;
        10'b101001110: data <= 20'b10011001000001001000;
        10'b101001111: data <= 20'b00011000010000111000;
        10'b101010000: data <= 20'b00010001110001000111;
        10'b101010001: data <= 20'b10001011000001001001;
        10'b101010010: data <= 20'b10010101100000100000;
        10'b101010011: data <= 20'b00010011011001100111;
        10'b101010100: data <= 20'b10010110011001010001;
        10'b101010101: data <= 20'b10011010101001010111;
        10'b101010110: data <= 20'b10010000010000011000;
        10'b101010111: data <= 20'b10010110110001100000;
        10'b101011000: data <= 20'b10011000001000011110;
        10'b101011001: data <= 20'b00000011011001011001;
        10'b101011010: data <= 20'b00010010010000011101;
        10'b101011011: data <= 20'b10011000111001010010;
        10'b101011100: data <= 20'b10000011110001010001;
        10'b101011101: data <= 20'b10011011100001100100;
        10'b101011110: data <= 20'b10011100111001101100;
        10'b101011111: data <= 20'b00100000101001101011;
        10'b101100000: data <= 20'b00010001000000001001;
        10'b101100001: data <= 20'b00011100001001000111;
        10'b101100010: data <= 20'b00011001101001101010;
        10'b101100011: data <= 20'b10011001101001001101;
        10'b101100100: data <= 20'b00001110110000000010;
        10'b101100101: data <= 20'b10001000111001000001;
        10'b101100110: data <= 20'b00010011101001010111;
        10'b101100111: data <= 20'b10010110001001010000;
        10'b101101000: data <= 20'b10001101111000101000;
        10'b101101001: data <= 20'b10010010100001000111;
        10'b101101010: data <= 20'b00010101110001011011;
        10'b101101011: data <= 20'b00010010101001000000;
        10'b101101100: data <= 20'b10001110101000111011;
        10'b101101101: data <= 20'b10010011011010000110;
        10'b101101110: data <= 20'b10010101011001011000;
        10'b101101111: data <= 20'b10011101111001110101;
        10'b101110000: data <= 20'b00011000101000110010;
        10'b101110001: data <= 20'b00010110010001001001;
        10'b101110010: data <= 20'b00001111010001011001;
        10'b101110011: data <= 20'b00001111111001000101;
        10'b101110100: data <= 20'b00010100011001011010;
        10'b101110101: data <= 20'b00011010101001100100;
        10'b101110110: data <= 20'b10010101000001010100;
        10'b101110111: data <= 20'b10000010110001010000;
        10'b101111000: data <= 20'b10010000000000110010;
        10'b101111001: data <= 20'b00010100010001000001;
        10'b101111010: data <= 20'b10000100101000110001;
        10'b101111011: data <= 20'b00001001000000110110;
        10'b101111100: data <= 20'b00001001111000101010;
        10'b101111101: data <= 20'b10010100110000101010;
        10'b101111110: data <= 20'b00001000010000111111;
        10'b101111111: data <= 20'b00001110001001010101;
        10'b110000000: data <= 20'b10001101110001000000;
        10'b110000001: data <= 20'b10001010010001001010;
        10'b110000010: data <= 20'b10010010100000110001;
        10'b110000011: data <= 20'b10010001100001010001;
        10'b110000100: data <= 20'b10001111001000110001;
        10'b110000101: data <= 20'b10010010001001010011;
        10'b110000110: data <= 20'b00010010000001010110;
        10'b110000111: data <= 20'b10010101111001001111;
        10'b110001000: data <= 20'b10001000011001100010;
        10'b110001001: data <= 20'b10011000001001011110;
        10'b110001010: data <= 20'b00001101110000111100;
        10'b110001011: data <= 20'b10010010000001000110;
        10'b110001100: data <= 20'b00010011000001011010;
        10'b110001101: data <= 20'b10011001001001011000;
        10'b110001110: data <= 20'b10010010001001110011;
        10'b110001111: data <= 20'b00011000010001011101;
        10'b110010000: data <= 20'b00010101011000000100;
        10'b110010001: data <= 20'b00010000110001000101;
        10'b110010010: data <= 20'b00010001000001001011;
        10'b110010011: data <= 20'b10011000000001000100;
        10'b110010100: data <= 20'b00011100011001101010;
        10'b110010101: data <= 20'b00010110111000111100;
        10'b110010110: data <= 20'b00010011010001101010;
        10'b110010111: data <= 20'b00001010010001010001;
        10'b110011000: data <= 20'b10001100111001001101;
        10'b110011001: data <= 20'b00001110010000100101;
        10'b110011010: data <= 20'b10001001010001000011;
        10'b110011011: data <= 20'b00000001001000100110;
        10'b110011100: data <= 20'b00010101101010000001;
        10'b110011101: data <= 20'b00000101011001011001;
        10'b110011110: data <= 20'b10011100001001011011;
        10'b110011111: data <= 20'b10000010110000101010;
        10'b110100000: data <= 20'b00001011111001000000;
        10'b110100001: data <= 20'b10010110110001001101;
        10'b110100010: data <= 20'b00000001011001000010;
        10'b110100011: data <= 20'b00010100000001011011;
        10'b110100100: data <= 20'b10011101001001010010;
        10'b110100101: data <= 20'b00001100011001100110;
        10'b110100110: data <= 20'b10010100111001010101;
        10'b110100111: data <= 20'b00000000101001010011;
        10'b110101000: data <= 20'b00010000111000011110;
        10'b110101001: data <= 20'b10000010010001010010;
        10'b110101010: data <= 20'b00011000100001100001;
        10'b110101011: data <= 20'b10011011101000111101;
        10'b110101100: data <= 20'b10011110001001110001;
        10'b110101101: data <= 20'b00001111011001001001;
        10'b110101110: data <= 20'b00011000111001010101;
        10'b110101111: data <= 20'b00001011000001100000;
        10'b110110000: data <= 20'b00001011100001011010;
        10'b110110001: data <= 20'b00001100111001000011;
        10'b110110010: data <= 20'b10011110001001110101;
        10'b110110011: data <= 20'b10010010111000100110;
        10'b110110100: data <= 20'b00010001100001101011;
        10'b110110101: data <= 20'b10010100110000110101;
        10'b110110110: data <= 20'b00010100111001100100;
        10'b110110111: data <= 20'b00001111010001011110;
        10'b110111000: data <= 20'b10010110000001010101;
        10'b110111001: data <= 20'b00010000010000101010;
        10'b110111010: data <= 20'b00010010011001000111;
        10'b110111011: data <= 20'b10010100100001000010;
        10'b110111100: data <= 20'b10010111010001011111;
        10'b110111101: data <= 20'b00001110001000110110;
        10'b110111110: data <= 20'b10010100100001101101;
        10'b110111111: data <= 20'b00001100111001000110;
        10'b111000000: data <= 20'b00001101110000110100;
        10'b111000001: data <= 20'b00010000000001000101;
        10'b111000010: data <= 20'b10010100111001010101;
        10'b111000011: data <= 20'b10001101100001001101;
        10'b111000100: data <= 20'b00001101010001010110;
        10'b111000101: data <= 20'b10001111100001010000;
        10'b111000110: data <= 20'b10011101001001100011;
        10'b111000111: data <= 20'b10010010111001100001;
        10'b111001000: data <= 20'b00010110011000010110;
        10'b111001001: data <= 20'b00001000110001001100;
        10'b111001010: data <= 20'b00001010010000101110;
        10'b111001011: data <= 20'b00010010000001100001;
        10'b111001100: data <= 20'b10011000010010001001;
        10'b111001101: data <= 20'b10010110101001010100;
        10'b111001110: data <= 20'b00010100101000100111;
        10'b111001111: data <= 20'b00010000001000110011;
        10'b111010000: data <= 20'b00010001001001001011;
        10'b111010001: data <= 20'b10001001111001110110;
        10'b111010010: data <= 20'b10010000000001010100;
        10'b111010011: data <= 20'b00010101010001001100;
        10'b111010100: data <= 20'b10010010100000100101;
        10'b111010101: data <= 20'b00011010001001110010;
        10'b111010110: data <= 20'b00010001011000110001;
        10'b111010111: data <= 20'b10001001100001000011;
        10'b111011000: data <= 20'b10010100111001011001;
        10'b111011001: data <= 20'b10001100011001000111;
        10'b111011010: data <= 20'b10001010100000010011;
        10'b111011011: data <= 20'b00010100010001000101;
        10'b111011100: data <= 20'b10010100001001000101;
        10'b111011101: data <= 20'b00010100100001011010;
        10'b111011110: data <= 20'b00001111000000001001;
        10'b111011111: data <= 20'b10010100000001011110;
        10'b111100000: data <= 20'b00001100011000101011;
        10'b111100001: data <= 20'b10101001011001001111;
        10'b111100010: data <= 20'b10001110011001001010;
        10'b111100011: data <= 20'b10010000011000011110;
        10'b111100100: data <= 20'b10010111010000111000;
        10'b111100101: data <= 20'b10010001001001000010;
        10'b111100110: data <= 20'b10010100110001100001;
        10'b111100111: data <= 20'b00010111100000101000;
        10'b111101000: data <= 20'b00001100011000110100;
        10'b111101001: data <= 20'b00001110011001000101;
        10'b111101010: data <= 20'b10010010011001110110;
        10'b111101011: data <= 20'b10010000010000001010;
        10'b111101100: data <= 20'b00001100001000110000;
        10'b111101101: data <= 20'b10011000111001100110;
        10'b111101110: data <= 20'b00010011001000101100;
        10'b111101111: data <= 20'b10001100000001000110;
        10'b111110000: data <= 20'b00000110011000110111;
        10'b111110001: data <= 20'b10001110111000100011;
        10'b111110010: data <= 20'b00010010100001111110;
        10'b111110011: data <= 20'b10010010011000111010;
        10'b111110100: data <= 20'b00010010010001001011;
        10'b111110101: data <= 20'b10000011100001011101;
        10'b111110110: data <= 20'b10001101101001011010;
        10'b111110111: data <= 20'b00010101001001100011;
        10'b111111000: data <= 20'b00010111100001011100;
        10'b111111001: data <= 20'b10011010100000110011;
        10'b111111010: data <= 20'b00001100010001000110;
        10'b111111011: data <= 20'b10000100000000101000;
        10'b111111100: data <= 20'b00001100100001001000;
        10'b111111101: data <= 20'b00001000010001011001;
        10'b111111110: data <= 20'b10010111101001001000;
        10'b111111111: data <= 20'b10010111000001001100;
        10'b1000000000: data <= 20'b00001010100001100110;
        10'b1000000001: data <= 20'b00010001000000111011;
        10'b1000000010: data <= 20'b00011000011001010100;
        10'b1000000011: data <= 20'b10000010111001101001;
        10'b1000000100: data <= 20'b10011111011001100000;
        10'b1000000101: data <= 20'b00010000100001100110;
        10'b1000000110: data <= 20'b00010001000001011010;
        10'b1000000111: data <= 20'b10100101000001011111;
        10'b1000001000: data <= 20'b10010011000001100001;
        10'b1000001001: data <= 20'b00010101001001111011;
        10'b1000001010: data <= 20'b10001000001001011010;
        10'b1000001011: data <= 20'b00010010100000010101;
        10'b1000001100: data <= 20'b10001100100001001110;
        10'b1000001101: data <= 20'b10010101000000111101;
        10'b1000001110: data <= 20'b00011010101001010100;
        10'b1000001111: data <= 20'b10001011001001001111;
        10'b1000010000: data <= 20'b00011010001001000110;
        10'b1000010001: data <= 20'b10001111011001100110;
        10'b1000010010: data <= 20'b00000000010001011010;
        10'b1000010011: data <= 20'b10001001010001011100;
        10'b1000010100: data <= 20'b10010010100001101001;
        10'b1000010101: data <= 20'b00011000110001000011;
        10'b1000010110: data <= 20'b00010011110001011100;
        10'b1000010111: data <= 20'b00011101110001100100;
        10'b1000011000: data <= 20'b00010010111000000110;
        10'b1000011001: data <= 20'b00001101010000101110;
        10'b1000011010: data <= 20'b00010010000001110001;
        10'b1000011011: data <= 20'b10011101101001100001;
        10'b1000011100: data <= 20'b10100011001010000000;
        10'b1000011101: data <= 20'b00011000000000100000;
        10'b1000011110: data <= 20'b10010011110001001010;
        10'b1000011111: data <= 20'b00010001000000101111;
        10'b1000100000: data <= 20'b00011010101001011111;
        10'b1000100001: data <= 20'b10000011101001011101;
        10'b1000100010: data <= 20'b00011100010001001100;
        10'b1000100011: data <= 20'b00100010111010000110;
        10'b1000100100: data <= 20'b00001111110001000010;
        10'b1000100101: data <= 20'b10001110001001010010;
        10'b1000100110: data <= 20'b00011100011001011011;
        10'b1000100111: data <= 20'b10001000001001011110;
        10'b1000101000: data <= 20'b10010100001001000101;
        10'b1000101001: data <= 20'b10010100101001011010;
        10'b1000101010: data <= 20'b00001101000001001001;
        10'b1000101011: data <= 20'b00011100101001101001;
        10'b1000101100: data <= 20'b00001100011001000000;
        10'b1000101101: data <= 20'b10010110000001011011;
        10'b1000101110: data <= 20'b00010111010001000001;
        10'b1000101111: data <= 20'b10011011111001010011;
        10'b1000110000: data <= 20'b00011101101001010001;
        10'b1000110001: data <= 20'b00010101110000110111;
        10'b1000110010: data <= 20'b00011000010000100101;
        10'b1000110011: data <= 20'b00011001010001010101;
        10'b1000110100: data <= 20'b00010111010001010011;
        10'b1000110101: data <= 20'b00010100100000001110;
        10'b1000110110: data <= 20'b00010000001000111110;
        10'b1000110111: data <= 20'b10010100011000001101;
        10'b1000111000: data <= 20'b10001000100001000101;
        10'b1000111001: data <= 20'b00010101101001101100;
        10'b1000111010: data <= 20'b10010001111001001010;
        10'b1000111011: data <= 20'b10001011110001000100;
        10'b1000111100: data <= 20'b00010111100001011100;
        10'b1000111101: data <= 20'b00001100011000011111;
        10'b1000111110: data <= 20'b00011001110001101110;
        10'b1000111111: data <= 20'b00010000001000100000;
        10'b1001000000: data <= 20'b10010000001001000111;
        10'b1001000001: data <= 20'b00010010100000001110;
        10'b1001000010: data <= 20'b00010000011001001111;
        10'b1001000011: data <= 20'b00010110001000000000;
        10'b1001000100: data <= 20'b10011000000000010110;
        10'b1001000101: data <= 20'b10001100101001001011;
        10'b1001000110: data <= 20'b00010011010000110000;
        10'b1001000111: data <= 20'b10010110110000111100;
        10'b1001001000: data <= 20'b00010000110001101010;
        10'b1001001001: data <= 20'b10001010011001100000;
        10'b1001001010: data <= 20'b10011001010001100010;
        10'b1001001011: data <= 20'b00010100101001001111;
        10'b1001001100: data <= 20'b00011000101001001111;
        10'b1001001101: data <= 20'b10011111100000010101;
        10'b1001001110: data <= 20'b00010100000000111010;
        10'b1001001111: data <= 20'b00010100110001001010;
        10'b1001010000: data <= 20'b00011000000001000001;
        10'b1001010001: data <= 20'b00001011000001011100;
        10'b1001010010: data <= 20'b00010001001001100111;
        10'b1001010011: data <= 20'b00010111001001101101;
        10'b1001010100: data <= 20'b10010001000000000110;
        10'b1001010101: data <= 20'b10001101100000101010;
        10'b1001010110: data <= 20'b10010100101001010000;
        10'b1001010111: data <= 20'b00011001011000000011;
        10'b1001011000: data <= 20'b10010111110001000011;
        10'b1001011001: data <= 20'b10010011011000000000;
        10'b1001011010: data <= 20'b00000100101000100011;
        10'b1001011011: data <= 20'b10001101100001010001;
        10'b1001011100: data <= 20'b00001001011001010110;
        10'b1001011101: data <= 20'b10000110011000101110;
        10'b1001011110: data <= 20'b00001100100001000100;
        10'b1001011111: data <= 20'b10010000101001010011;
        10'b1001100000: data <= 20'b00010000101001010000;
        10'b1001100001: data <= 20'b10010000001001000111;
        10'b1001100010: data <= 20'b10010101000000101011;
        10'b1001100011: data <= 20'b10010000110001000101;
        10'b1001100100: data <= 20'b00001111100000101100;
        10'b1001100101: data <= 20'b00011001100001010000;
        10'b1001100110: data <= 20'b00010001010000110110;
        10'b1001100111: data <= 20'b00001010110001011000;
        10'b1001101000: data <= 20'b10010001011001000001;
        10'b1001101001: data <= 20'b10010100101001000011;
        10'b1001101010: data <= 20'b10010100100001001110;
        10'b1001101011: data <= 20'b00010100001001000001;
        10'b1001101100: data <= 20'b10010000010001000001;
        10'b1001101101: data <= 20'b10000111101000000000;
        10'b1001101110: data <= 20'b00010110101001011011;
        10'b1001101111: data <= 20'b10000100100001010000;
        10'b1001110000: data <= 20'b10011000111001100000;
        10'b1001110001: data <= 20'b10001100100001011001;
        10'b1001110010: data <= 20'b10001010000001011010;
        10'b1001110011: data <= 20'b00001110100000111011;
        10'b1001110100: data <= 20'b10001110011001000001;
        10'b1001110101: data <= 20'b00010110010001001101;
        10'b1001110110: data <= 20'b10011011011001010110;
        10'b1001110111: data <= 20'b10010101110001001100;
        10'b1001111000: data <= 20'b10001011110001100000;
        10'b1001111001: data <= 20'b00010000100001011011;
        10'b1001111010: data <= 20'b10000011010001000000;
        10'b1001111011: data <= 20'b00011000000001100000;
        10'b1001111100: data <= 20'b10010111001001011100;
        10'b1001111101: data <= 20'b00011100010001100101;
        10'b1001111110: data <= 20'b10001000100001010010;
        10'b1001111111: data <= 20'b00010010010001010111;
        10'b1010000000: data <= 20'b10001110110001011100;
        10'b1010000001: data <= 20'b10001001001001000010;
        10'b1010000010: data <= 20'b10010111111001000001;
        10'b1010000011: data <= 20'b10010011011001001101;
        10'b1010000100: data <= 20'b10001110000001001010;
        10'b1010000101: data <= 20'b10010100100001000010;
        10'b1010000110: data <= 20'b00011111011001110100;
        10'b1010000111: data <= 20'b10010010011001101100;
        10'b1010001000: data <= 20'b00010010101001001101;
        10'b1010001001: data <= 20'b10000011000000111101;
        10'b1010001010: data <= 20'b00000100100000111100;
        10'b1010001011: data <= 20'b10010011011001010111;
        10'b1010001100: data <= 20'b10011100011001110011;
        10'b1010001101: data <= 20'b10000100011001110110;
        10'b1010001110: data <= 20'b10010000100001001100;
        10'b1010001111: data <= 20'b00000000000001000101;
        10'b1010010000: data <= 20'b10001110001001010010;
        10'b1010010001: data <= 20'b10010100000001011011;
        10'b1010010010: data <= 20'b00010100110000110101;
        10'b1010010011: data <= 20'b10001111110001010010;
        10'b1010010100: data <= 20'b10010000110001011010;
        10'b1010010101: data <= 20'b10100111010010010010;
        10'b1010010110: data <= 20'b00010111111001001010;
        10'b1010010111: data <= 20'b10010001010001001011;
        10'b1010011000: data <= 20'b00010001010001000010;
        10'b1010011001: data <= 20'b00011001111001011111;
        10'b1010011010: data <= 20'b00100000111001111011;
        10'b1010011011: data <= 20'b00010001010000111000;
        10'b1010011100: data <= 20'b10001010111001000111;
        10'b1010011101: data <= 20'b10000110000000100101;
        10'b1010011110: data <= 20'b00000011011001100010;
        10'b1010011111: data <= 20'b10010010000001000000;
        10'b1010100000: data <= 20'b10001010001000111101;
        10'b1010100001: data <= 20'b00001101101001010000;
        10'b1010100010: data <= 20'b10010000100001010100;
        10'b1010100011: data <= 20'b10001001101001010001;
        10'b1010100100: data <= 20'b00000010000001011011;
        10'b1010100101: data <= 20'b00001110000000101010;
        10'b1010100110: data <= 20'b10011010000001010101;
        10'b1010100111: data <= 20'b00011110101001011111;
        10'b1010101000: data <= 20'b10010101000000110001;
        10'b1010101001: data <= 20'b10010000100000010000;
        10'b1010101010: data <= 20'b10010101110001100010;
        10'b1010101011: data <= 20'b10100010010001011000;
        10'b1010101100: data <= 20'b00010110101000101100;
        10'b1010101101: data <= 20'b00011010001000100101;
        10'b1010101110: data <= 20'b00001001011000110110;
        10'b1010101111: data <= 20'b10010101100000001000;
        10'b1010110000: data <= 20'b10010000011000001101;
        10'b1010110001: data <= 20'b10001111101000111101;
        10'b1010110010: data <= 20'b10010100101000111111;
        10'b1010110011: data <= 20'b00010000101001000100;
        10'b1010110100: data <= 20'b00010111101001010110;
        10'b1010110101: data <= 20'b10010101001001100000;
        10'b1010110110: data <= 20'b10011100011001101011;
        10'b1010110111: data <= 20'b00010101111000111110;
        10'b1010111000: data <= 20'b00010000010001010001;
        10'b1010111001: data <= 20'b00001011100001001110;
        10'b1010111010: data <= 20'b10011010111000101100;
        10'b1010111011: data <= 20'b00010011101001001101;
        10'b1010111100: data <= 20'b10001110101001100110;
        10'b1010111101: data <= 20'b00010101010001010010;
        10'b1010111110: data <= 20'b10010111100001010001;
        10'b1010111111: data <= 20'b00011000010001101100;
        10'b1011000000: data <= 20'b00010100010001101000;
        10'b1011000001: data <= 20'b00010001111001000010;
        10'b1011000010: data <= 20'b00001101101001000011;
        10'b1011000011: data <= 20'b10010000100000111010;
        10'b1011000100: data <= 20'b00000000011001001010;
        10'b1011000101: data <= 20'b00001010001000111100;
        10'b1011000110: data <= 20'b00010000101001000110;
        10'b1011000111: data <= 20'b10011011100000101111;
        10'b1011001000: data <= 20'b10010100001000001010;
        10'b1011001001: data <= 20'b00010000111001010110;
        10'b1011001010: data <= 20'b00011000000000010100;
        10'b1011001011: data <= 20'b10010001010000000110;
        10'b1011001100: data <= 20'b00001110000001000110;
        10'b1011001101: data <= 20'b00010001001000101000;
        10'b1011001110: data <= 20'b00001100111001100110;
        10'b1011001111: data <= 20'b10011010100001011100;
        10'b1011010000: data <= 20'b10001001111001010111;
        10'b1011010001: data <= 20'b00001100001001010100;
        10'b1011010010: data <= 20'b10001111011001001001;
        10'b1011010011: data <= 20'b00011000110001010001;
        10'b1011010100: data <= 20'b10010100011000011010;
        10'b1011010101: data <= 20'b00010010001001101011;
        10'b1011010110: data <= 20'b00010111010001000000;
        10'b1011010111: data <= 20'b00001100101001011001;
        10'b1011011000: data <= 20'b10001111110001011100;
        10'b1011011001: data <= 20'b00011000101000111010;
        10'b1011011010: data <= 20'b10010011101001011100;
        10'b1011011011: data <= 20'b00000111101000100000;
        10'b1011011100: data <= 20'b10010001001001010001;
        10'b1011011101: data <= 20'b00010000110001010100;
        10'b1011011110: data <= 20'b00001000100000100101;
        10'b1011011111: data <= 20'b10001110001000001010;
        10'b1011100000: data <= 20'b10010101101000110010;
        10'b1011100001: data <= 20'b00000000011001010110;
        10'b1011100010: data <= 20'b10010101111001101101;
        10'b1011100011: data <= 20'b00011110110001010001;
        10'b1011100100: data <= 20'b00011001001001011111;
        10'b1011100101: data <= 20'b10001101000001100100;
        10'b1011100110: data <= 20'b00010011010000111010;
        10'b1011100111: data <= 20'b00010110111000110010;
        10'b1011101000: data <= 20'b10001100111001011010;
        10'b1011101001: data <= 20'b10011111001001101111;
        10'b1011101010: data <= 20'b00010101011001011101;
        10'b1011101011: data <= 20'b00010000000001010100;
        10'b1011101100: data <= 20'b00010001111000011010;
        10'b1011101101: data <= 20'b00010101110000110010;
        10'b1011101110: data <= 20'b00001100100001010110;
        10'b1011101111: data <= 20'b10010110010000110110;
        10'b1011110000: data <= 20'b00010101000001101100;
        10'b1011110001: data <= 20'b10001000010001001000;
        10'b1011110010: data <= 20'b10100000101000100100;
        10'b1011110011: data <= 20'b00011001101001100010;
        10'b1011110100: data <= 20'b10010010001001010011;
        10'b1011110101: data <= 20'b00001110101000100000;
        10'b1011110110: data <= 20'b00010100100001010111;
        10'b1011110111: data <= 20'b00011010001001100001;
        10'b1011111000: data <= 20'b10011011100001100101;
        10'b1011111001: data <= 20'b00010000110001001111;
        10'b1011111010: data <= 20'b10001101100001000101;
        10'b1011111011: data <= 20'b00000011000000011010;
        10'b1011111100: data <= 20'b10001101111000101000;
        10'b1011111101: data <= 20'b00000100100001010000;
        10'b1011111110: data <= 20'b00010100000001101100;
        10'b1011111111: data <= 20'b10010101000000110100;
        10'b1100000000: data <= 20'b10001100010000110010;
        10'b1100000001: data <= 20'b10001100111001001100;
        10'b1100000010: data <= 20'b00010100000000111010;
        10'b1100000011: data <= 20'b10010001011001000110;
        10'b1100000100: data <= 20'b10010111000001100011;
        10'b1100000101: data <= 20'b10010101000000000110;
        10'b1100000110: data <= 20'b00000010011001100001;
        10'b1100000111: data <= 20'b00010011011001010010;
        10'b1100001000: data <= 20'b00010100000001101010;
        10'b1100001001: data <= 20'b10011100100000110110;
        10'b1100001010: data <= 20'b00010101011001101111;
        10'b1100001011: data <= 20'b00001100110000111011;
        10'b1100001100: data <= 20'b00010111001001011001;
        10'b1100001101: data <= 20'b00010011010000000100;
        10'b1100001110: data <= 20'b10001011001000110001;
        10'b1100001111: data <= 20'b00000011001001001110;
        10'b1100010000: data <= 20'b10011000110001100111;
        10'b1100010001: data <= 20'b10011001111001001010;
        10'b1100010010: data <= 20'b00010010010001010000;
        10'b1100010011: data <= 20'b00010100100001000111;
        10'b1100010100: data <= 20'b10010001011001110100;
        10'b1100010101: data <= 20'b00011110001001101001;
        10'b1100010110: data <= 20'b10001100110001001001;
        10'b1100010111: data <= 20'b10010100001000110111;
        10'b1100011000: data <= 20'b10001010011001010001;
        10'b1100011001: data <= 20'b00001111001000000011;
        10'b1100011010: data <= 20'b00011001011001101010;
        10'b1100011011: data <= 20'b10010100011001011011;
        10'b1100011100: data <= 20'b00010010000001110011;
        10'b1100011101: data <= 20'b00011000010000011000;
        10'b1100011110: data <= 20'b00010011110001000010;
        10'b1100011111: data <= 20'b00010101111001011011;
        10'b1100100000: data <= 20'b10010110100001001101;
        10'b1100100001: data <= 20'b10011100110001010001;
        10'b1100100010: data <= 20'b10010101101001010000;
        10'b1100100011: data <= 20'b00010100011001001001;
        10'b1100100100: data <= 20'b00010100001000111110;
        10'b1100100101: data <= 20'b00010100010001001000;
        10'b1100100110: data <= 20'b00001010110000011010;
        10'b1100100111: data <= 20'b00001000010000111000;
        10'b1100101000: data <= 20'b10001110100000100001;
        10'b1100101001: data <= 20'b00010110001001010011;
        10'b1100101010: data <= 20'b00001111110001000000;
        10'b1100101011: data <= 20'b10010100100000000000;
        10'b1100101100: data <= 20'b10010000001000100110;
        10'b1100101101: data <= 20'b10010100011000100010;
        10'b1100101110: data <= 20'b10010001001001010001;
        10'b1100101111: data <= 20'b10010001100001100101;
        10'b1100110000: data <= 20'b00001100111001000010;
        10'b1100110001: data <= 20'b10010101110001000100;
        10'b1100110010: data <= 20'b10011111110001110000;
        10'b1100110011: data <= 20'b10010011111000101101;
        10'b1100110100: data <= 20'b00010101001000111101;
        10'b1100110101: data <= 20'b00001110111000101010;
        10'b1100110110: data <= 20'b10001100010000111001;
        10'b1100110111: data <= 20'b10000110011000011100;
        10'b1100111000: data <= 20'b00010000001000001011;
        10'b1100111001: data <= 20'b10011000111001101000;
        10'b1100111010: data <= 20'b00000011011001011011;
        10'b1100111011: data <= 20'b10010111011001000111;
        10'b1100111100: data <= 20'b00000100001001000010;
        10'b1100111101: data <= 20'b00010111111001101100;
        10'b1100111110: data <= 20'b10001100110001000101;
        10'b1100111111: data <= 20'b00001000101001010010;
        10'b1101000000: data <= 20'b00001011100001010010;
        10'b1101000001: data <= 20'b00000001001001011101;
        10'b1101000010: data <= 20'b00010111011001010110;
        10'b1101000011: data <= 20'b00010000001000111100;
        10'b1101000100: data <= 20'b00010000011000101010;
        10'b1101000101: data <= 20'b10001001011001000011;
        10'b1101000110: data <= 20'b00010011011000111101;
        10'b1101000111: data <= 20'b10010000001001010100;
        10'b1101001000: data <= 20'b10001100011001000001;
        10'b1101001001: data <= 20'b00010111010001011100;
        10'b1101001010: data <= 20'b10010000011001010000;
        10'b1101001011: data <= 20'b00000001000001001110;
        10'b1101001100: data <= 20'b10000110011000110100;
        10'b1101001101: data <= 20'b10011000110001010001;
        10'b1101001110: data <= 20'b10010100001000110111;
        10'b1101001111: data <= 20'b10010111111001000000;
        10'b1101010000: data <= 20'b10001111100001010110;
        10'b1101010001: data <= 20'b00001101111001000010;
        10'b1101010010: data <= 20'b00010010011000100111;
        10'b1101010011: data <= 20'b10010100000000001001;
        10'b1101010100: data <= 20'b10001000011000001001;
        10'b1101010101: data <= 20'b00010011010001001000;
        10'b1101010110: data <= 20'b10010011011001001110;
        10'b1101010111: data <= 20'b10010000001001010111;
        10'b1101011000: data <= 20'b00011111010001001011;
        10'b1101011001: data <= 20'b00001110001001100110;
        10'b1101011010: data <= 20'b10011111111001110101;
        10'b1101011011: data <= 20'b10010000011001110101;
        10'b1101011100: data <= 20'b00000010001000011111;
        10'b1101011101: data <= 20'b00011001010001101010;
        10'b1101011110: data <= 20'b10001101111001110111;
        10'b1101011111: data <= 20'b10010101001000110110;
        10'b1101100000: data <= 20'b00001011010001100001;
        10'b1101100001: data <= 20'b00000000010000111100;
        10'b1101100010: data <= 20'b00001111011001001010;
        10'b1101100011: data <= 20'b00001011011001101111;
        10'b1101100100: data <= 20'b00001100000001101010;
        10'b1101100101: data <= 20'b00010011101001010010;
        10'b1101100110: data <= 20'b00010100100001000000;
        10'b1101100111: data <= 20'b10010101000001101011;
        10'b1101101000: data <= 20'b00100000001001100011;
        10'b1101101001: data <= 20'b10000101000001010011;
        10'b1101101010: data <= 20'b00001110010001011001;
        10'b1101101011: data <= 20'b10001110100000111000;
        10'b1101101100: data <= 20'b00000111001000011100;
        10'b1101101101: data <= 20'b00001100101001001111;
        10'b1101101110: data <= 20'b10001110101000100001;
        10'b1101101111: data <= 20'b10010100011000101001;
        10'b1101110000: data <= 20'b10001011111000111011;
        10'b1101110001: data <= 20'b00010001110001010000;
        10'b1101110010: data <= 20'b00001100101001001011;
        10'b1101110011: data <= 20'b10010010110001010010;
        10'b1101110100: data <= 20'b10010001000001100111;
        10'b1101110101: data <= 20'b10010110011001101010;
        10'b1101110110: data <= 20'b10010000001000001110;
        10'b1101110111: data <= 20'b10001111010000111111;
        10'b1101111000: data <= 20'b10010100010001001000;
        10'b1101111001: data <= 20'b00010010001001000011;
        10'b1101111010: data <= 20'b00100000101010001010;
        10'b1101111011: data <= 20'b00010010001001010101;
        10'b1101111100: data <= 20'b10010101111001010111;
        10'b1101111101: data <= 20'b00010100100000111011;
        10'b1101111110: data <= 20'b00011000000001100110;
        10'b1101111111: data <= 20'b00001010010001010100;
        10'b1110000000: data <= 20'b10010101101001110101;
        10'b1110000001: data <= 20'b00011011011001110001;
        10'b1110000010: data <= 20'b10001111100001100001;
        10'b1110000011: data <= 20'b00001001010001100000;
        10'b1110000100: data <= 20'b00010100101001100111;
        10'b1110000101: data <= 20'b00010100101000000101;
        10'b1110000110: data <= 20'b00010101111001000101;
        10'b1110000111: data <= 20'b10001110000001011101;
        10'b1110001000: data <= 20'b00001101111001000011;
        10'b1110001001: data <= 20'b00001100011001010000;
        10'b1110001010: data <= 20'b00001000011000100100;
        10'b1110001011: data <= 20'b00001011001001010000;
        10'b1110001100: data <= 20'b10010101101000101001;
        10'b1110001101: data <= 20'b10010110111000101111;
        10'b1110001110: data <= 20'b00001001111001001000;
        10'b1110001111: data <= 20'b10011011000001001100;
        10'b1110010000: data <= 20'b00010001000001100101;
        10'b1110010001: data <= 20'b00011000111001110000;
        10'b1110010010: data <= 20'b00001100100001100001;
        10'b1110010011: data <= 20'b00010111010001000100;
        10'b1110010100: data <= 20'b00010100001001010001;
        10'b1110010101: data <= 20'b00001110101001001101;
        10'b1110010110: data <= 20'b00010000111001010100;
        10'b1110010111: data <= 20'b10010001110000110101;
        10'b1110011000: data <= 20'b00010110011000111010;
        10'b1110011001: data <= 20'b10010101010001000010;
        10'b1110011010: data <= 20'b00000001001001001000;
        10'b1110011011: data <= 20'b00010010001001000101;
        10'b1110011100: data <= 20'b00010101000001010000;
        10'b1110011101: data <= 20'b00010100001001100001;
        10'b1110011110: data <= 20'b10011000110001000001;
        10'b1110011111: data <= 20'b10010110000001110001;
        10'b1110100000: data <= 20'b00010100111000011101;
        10'b1110100001: data <= 20'b00011100010001100110;
        10'b1110100010: data <= 20'b10011111000001110010;
        10'b1110100011: data <= 20'b00011100011001001111;
        10'b1110100100: data <= 20'b00011001010001000101;
        10'b1110100101: data <= 20'b10010101101000111010;
        10'b1110100110: data <= 20'b10010011110001010001;
        10'b1110100111: data <= 20'b10011000011001100001;
        10'b1110101000: data <= 20'b10010001101000110111;
        10'b1110101001: data <= 20'b00010110111001001110;
        10'b1110101010: data <= 20'b10010011101001101000;
        10'b1110101011: data <= 20'b00010001010000110100;
        10'b1110101100: data <= 20'b00010011110001000001;
        10'b1110101101: data <= 20'b10011000000001001000;
        10'b1110101110: data <= 20'b10010111100001001000;
        10'b1110101111: data <= 20'b10001010000001001101;
        10'b1110110000: data <= 20'b00010001000000010100;
        10'b1110110001: data <= 20'b00011101011000111010;
        10'b1110110010: data <= 20'b00010011010001111111;
        10'b1110110011: data <= 20'b10011101110001100001;
        10'b1110110100: data <= 20'b10001110100001001110;
        10'b1110110101: data <= 20'b00010100010000110000;
        10'b1110110110: data <= 20'b00010100001001000001;
        10'b1110110111: data <= 20'b10011000001001011010;
        10'b1110111000: data <= 20'b10010001000001001100;
        10'b1110111001: data <= 20'b10000011100000101111;
        10'b1110111010: data <= 20'b10011010111001100011;
        10'b1110111011: data <= 20'b00011001100001001011;
        10'b1110111100: data <= 20'b10001101111001000100;
        10'b1110111101: data <= 20'b10010000111001000000;
        10'b1110111110: data <= 20'b10010100011001001110;
        10'b1110111111: data <= 20'b00011000110000001111;
        10'b1111000000: data <= 20'b10000000101001011001;
        10'b1111000001: data <= 20'b00011001010001100000;
        10'b1111000010: data <= 20'b00010100011000101101;
        10'b1111000011: data <= 20'b10001110101001010110;
        10'b1111000100: data <= 20'b10001100010000001110;
        10'b1111000101: data <= 20'b00010010011000111101;
        10'b1111000110: data <= 20'b10010010011000000111;
        10'b1111000111: data <= 20'b10000011001001011110;
        10'b1111001000: data <= 20'b10011010001001100111;
        10'b1111001001: data <= 20'b00011000101000010000;
        10'b1111001010: data <= 20'b10000010110001100001;
        10'b1111001011: data <= 20'b00001111111000000000;
        10'b1111001100: data <= 20'b00010000011000110010;
        10'b1111001101: data <= 20'b00011011001001101001;
        10'b1111001110: data <= 20'b10010110001000110001;
        10'b1111001111: data <= 20'b00010000110001011001;
        10'b1111010000: data <= 20'b00010000101000010010;
        10'b1111010001: data <= 20'b00010110101001010111;
        10'b1111010010: data <= 20'b10010011100000111010;
        10'b1111010011: data <= 20'b10010101110001011010;
        10'b1111010100: data <= 20'b10010100001000100111;
        10'b1111010101: data <= 20'b00010100000001000111;
        10'b1111010110: data <= 20'b10010100000001101010;
        10'b1111010111: data <= 20'b10010100011000100000;
        10'b1111011000: data <= 20'b10100100100001100011;
        10'b1111011001: data <= 20'b00010110111001000000;
        10'b1111011010: data <= 20'b00010111111001000110;
        10'b1111011011: data <= 20'b00001111010001001010;
        10'b1111011100: data <= 20'b00011001001000001011;
        10'b1111011101: data <= 20'b00001000101001011001;
        10'b1111011110: data <= 20'b10011010110000101001;
        10'b1111011111: data <= 20'b00001111010001001000;
        10'b1111100000: data <= 20'b10011000001000011011;
        10'b1111100001: data <= 20'b00010111000000101001;
        10'b1111100010: data <= 20'b10011110110000110111;
        10'b1111100011: data <= 20'b00011100110001010111;
        10'b1111100100: data <= 20'b10001101000001101010;
        10'b1111100101: data <= 20'b00010101111000110010;
        10'b1111100110: data <= 20'b10011011100001001010;
        10'b1111100111: data <= 20'b00011000000001000110;
        10'b1111101000: data <= 20'b10100000001000111010;
        10'b1111101001: data <= 20'b00010001001001000010;
        10'b1111101010: data <= 20'b00011000110000101001;
        10'b1111101011: data <= 20'b00010011100000110001;
        10'b1111101100: data <= 20'b10011110000001110000;
        10'b1111101101: data <= 20'b10001000011001001101;
        10'b1111101110: data <= 20'b00001111001000111110;
        10'b1111101111: data <= 20'b00000100111001000101;
        10'b1111110000: data <= 20'b00010110000001001010;
        10'b1111110001: data <= 20'b10010000011001011111;
        10'b1111110010: data <= 20'b10010001111001011011;
        10'b1111110011: data <= 20'b00011010101001110000;
        10'b1111110100: data <= 20'b00001011011001101010;
        10'b1111110101: data <= 20'b10010011001000101010;
        10'b1111110110: data <= 20'b00000010110001010001;
        10'b1111110111: data <= 20'b00010101100001000000;
        10'b1111111000: data <= 20'b10010000111001000111;
        10'b1111111001: data <= 20'b10000100100001010111;
        10'b1111111010: data <= 20'b10010111101001110110;
        10'b1111111011: data <= 20'b10010000000001011000;
        10'b1111111100: data <= 20'b10001101001001011000;
    
    endcase
    end
    end

    assign Q = data;

    endmodule

        