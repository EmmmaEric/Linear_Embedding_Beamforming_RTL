
module memory_rom_3(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbafbbd50;
    11'b00000000001: data <= 32'hb788b94e;
    11'b00000000010: data <= 32'h37f23b23;
    11'b00000000011: data <= 32'h2f273f7d;
    11'b00000000100: data <= 32'hbdcf3bad;
    11'b00000000101: data <= 32'hc084b9d3;
    11'b00000000110: data <= 32'hbe02bb76;
    11'b00000000111: data <= 32'hb554379c;
    11'b00000001000: data <= 32'h347f3d50;
    11'b00000001001: data <= 32'h3a483800;
    11'b00000001010: data <= 32'h3e1ab661;
    11'b00000001011: data <= 32'h3e5f361c;
    11'b00000001100: data <= 32'h360e3fad;
    11'b00000001101: data <= 32'hbab93fcf;
    11'b00000001110: data <= 32'hb73c3279;
    11'b00000001111: data <= 32'h3b96bda7;
    11'b00000010000: data <= 32'h3d21be99;
    11'b00000010001: data <= 32'h316abd0a;
    11'b00000010010: data <= 32'hb73abc86;
    11'b00000010011: data <= 32'h38aeba8c;
    11'b00000010100: data <= 32'h3ea33059;
    11'b00000010101: data <= 32'h39be3a56;
    11'b00000010110: data <= 32'hbe4c30ed;
    11'b00000010111: data <= 32'hc16cbb6b;
    11'b00000011000: data <= 32'hbf46ba87;
    11'b00000011001: data <= 32'hb7b734a5;
    11'b00000011010: data <= 32'hac84388e;
    11'b00000011011: data <= 32'haa95b6d8;
    11'b00000011100: data <= 32'h367aba6a;
    11'b00000011101: data <= 32'h39f73a53;
    11'b00000011110: data <= 32'h3204418b;
    11'b00000011111: data <= 32'hb8834157;
    11'b00000100000: data <= 32'hb4bf38cf;
    11'b00000100001: data <= 32'h38d5bc0f;
    11'b00000100010: data <= 32'h3987bb39;
    11'b00000100011: data <= 32'ha427b452;
    11'b00000100100: data <= 32'h310cb6ae;
    11'b00000100101: data <= 32'h3ed8ba5b;
    11'b00000100110: data <= 32'h4150b66f;
    11'b00000100111: data <= 32'h3cf43426;
    11'b00000101000: data <= 32'hbd2f2d02;
    11'b00000101001: data <= 32'hc07eb955;
    11'b00000101010: data <= 32'hbc83ba65;
    11'b00000101011: data <= 32'ha453b61f;
    11'b00000101100: data <= 32'hb48cb904;
    11'b00000101101: data <= 32'hbb0bbe0f;
    11'b00000101110: data <= 32'hb79fbd39;
    11'b00000101111: data <= 32'h355d3a0a;
    11'b00000110000: data <= 32'h334a4176;
    11'b00000110001: data <= 32'hb8c340cf;
    11'b00000110010: data <= 32'hbb073703;
    11'b00000110011: data <= 32'hb767b8c1;
    11'b00000110100: data <= 32'hb4943069;
    11'b00000110101: data <= 32'hb5ea3ada;
    11'b00000110110: data <= 32'h36c53237;
    11'b00000110111: data <= 32'h4040ba3a;
    11'b00000111000: data <= 32'h41b5b7e1;
    11'b00000111001: data <= 32'h3d7a38c3;
    11'b00000111010: data <= 32'hba283aee;
    11'b00000111011: data <= 32'hbca92be0;
    11'b00000111100: data <= 32'h2c38b975;
    11'b00000111101: data <= 32'h3923bb8e;
    11'b00000111110: data <= 32'hb5c4bdb6;
    11'b00000111111: data <= 32'hbcfbc02e;
    11'b00001000000: data <= 32'hb824be97;
    11'b00001000001: data <= 32'h3a1b340c;
    11'b00001000010: data <= 32'h39623f3e;
    11'b00001000011: data <= 32'hb9a53d70;
    11'b00001000100: data <= 32'hbeacaf06;
    11'b00001000101: data <= 32'hbe0db553;
    11'b00001000110: data <= 32'hbc4b3ac8;
    11'b00001000111: data <= 32'hba2c3d57;
    11'b00001001000: data <= 32'h2d5c308f;
    11'b00001001001: data <= 32'h3e1dbbfa;
    11'b00001001010: data <= 32'h4045b44b;
    11'b00001001011: data <= 32'h3c423de2;
    11'b00001001100: data <= 32'hb4a44000;
    11'b00001001101: data <= 32'hb0ce3b04;
    11'b00001001110: data <= 32'h3b75b648;
    11'b00001001111: data <= 32'h3b49bb2d;
    11'b00001010000: data <= 32'hb758bcfe;
    11'b00001010001: data <= 32'hbc53bf25;
    11'b00001010010: data <= 32'h33d4be91;
    11'b00001010011: data <= 32'h3f3ab6b2;
    11'b00001010100: data <= 32'h3d7e38e1;
    11'b00001010101: data <= 32'hb9323436;
    11'b00001010110: data <= 32'hbffdb882;
    11'b00001010111: data <= 32'hbf1bb359;
    11'b00001011000: data <= 32'hbca23b3c;
    11'b00001011001: data <= 32'hbc0c3b0b;
    11'b00001011010: data <= 32'hb97db92f;
    11'b00001011011: data <= 32'h34d6bdff;
    11'b00001011100: data <= 32'h3c0fac9c;
    11'b00001011101: data <= 32'h38e44054;
    11'b00001011110: data <= 32'haae14154;
    11'b00001011111: data <= 32'h33663d05;
    11'b00001100000: data <= 32'h3b37aa34;
    11'b00001100001: data <= 32'h37a4b20e;
    11'b00001100010: data <= 32'hb9e8b150;
    11'b00001100011: data <= 32'hb9a8ba96;
    11'b00001100100: data <= 32'h3cbabd6f;
    11'b00001100101: data <= 32'h417fbb2a;
    11'b00001100110: data <= 32'h3fa8b033;
    11'b00001100111: data <= 32'hb5deb056;
    11'b00001101000: data <= 32'hbe26b7d2;
    11'b00001101001: data <= 32'hbc04b047;
    11'b00001101010: data <= 32'hb7a337b2;
    11'b00001101011: data <= 32'hbbdfae8b;
    11'b00001101100: data <= 32'hbdc5beb7;
    11'b00001101101: data <= 32'hba28c01e;
    11'b00001101110: data <= 32'h3468b154;
    11'b00001101111: data <= 32'h36fc4030;
    11'b00001110000: data <= 32'ha77440a8;
    11'b00001110001: data <= 32'hae1c3b54;
    11'b00001110010: data <= 32'h2cb53126;
    11'b00001110011: data <= 32'hb6f23a3b;
    11'b00001110100: data <= 32'hbcb53c8a;
    11'b00001110101: data <= 32'hb8662f78;
    11'b00001110110: data <= 32'h3e26bc68;
    11'b00001110111: data <= 32'h41c6bc0e;
    11'b00001111000: data <= 32'h3fa8aa54;
    11'b00001111001: data <= 32'ha18d363c;
    11'b00001111010: data <= 32'hb8283104;
    11'b00001111011: data <= 32'h359f2d88;
    11'b00001111100: data <= 32'h38052c7b;
    11'b00001111101: data <= 32'hba6aba85;
    11'b00001111110: data <= 32'hbf3dc06c;
    11'b00001111111: data <= 32'hbc3cc0a3;
    11'b00010000000: data <= 32'h36aeb85c;
    11'b00010000001: data <= 32'h3a2f3ce3;
    11'b00010000010: data <= 32'ha82a3c8a;
    11'b00010000011: data <= 32'hb9992be1;
    11'b00010000100: data <= 32'hbae13111;
    11'b00010000101: data <= 32'hbcc33de1;
    11'b00010000110: data <= 32'hbe323f6c;
    11'b00010000111: data <= 32'hba8c35f4;
    11'b00010001000: data <= 32'h3bc3bcb9;
    11'b00010001001: data <= 32'h4014bb1b;
    11'b00010001010: data <= 32'h3d4f38ed;
    11'b00010001011: data <= 32'h32b33d83;
    11'b00010001100: data <= 32'h376b3b93;
    11'b00010001101: data <= 32'h3dd03648;
    11'b00010001110: data <= 32'h3c632e6b;
    11'b00010001111: data <= 32'hb9d4b929;
    11'b00010010000: data <= 32'hbee9bf32;
    11'b00010010001: data <= 32'hb82ec022;
    11'b00010010010: data <= 32'h3d26bbca;
    11'b00010010011: data <= 32'h3dc72bab;
    11'b00010010100: data <= 32'h2cffb21b;
    11'b00010010101: data <= 32'hbbf4b9df;
    11'b00010010110: data <= 32'hbc732b85;
    11'b00010010111: data <= 32'hbcc73e5d;
    11'b00010011000: data <= 32'hbe5b3e8d;
    11'b00010011001: data <= 32'hbd7eb2eb;
    11'b00010011010: data <= 32'hb2eabe91;
    11'b00010011011: data <= 32'h3998ba2b;
    11'b00010011100: data <= 32'h38303ced;
    11'b00010011101: data <= 32'h32ed4005;
    11'b00010011110: data <= 32'h3b203d13;
    11'b00010011111: data <= 32'h3eaf38b9;
    11'b00010100000: data <= 32'h3b2e390f;
    11'b00010100001: data <= 32'hbb943664;
    11'b00010100010: data <= 32'hbdc8b90e;
    11'b00010100011: data <= 32'h34cebdbe;
    11'b00010100100: data <= 32'h405abccf;
    11'b00010100101: data <= 32'h3fceb9ad;
    11'b00010100110: data <= 32'h3447bac8;
    11'b00010100111: data <= 32'hb952bb6a;
    11'b00010101000: data <= 32'hb5ee2c47;
    11'b00010101001: data <= 32'hb54c3d0f;
    11'b00010101010: data <= 32'hbceb3a66;
    11'b00010101011: data <= 32'hbf80bcaf;
    11'b00010101100: data <= 32'hbd35c05e;
    11'b00010101101: data <= 32'hb4e5ba91;
    11'b00010101110: data <= 32'h29d73cfc;
    11'b00010101111: data <= 32'h2fa53ec8;
    11'b00010110000: data <= 32'h39473a32;
    11'b00010110001: data <= 32'h3c1037fc;
    11'b00010110010: data <= 32'h2d903d68;
    11'b00010110011: data <= 32'hbd823ed1;
    11'b00010110100: data <= 32'hbd26389d;
    11'b00010110101: data <= 32'h3997bac6;
    11'b00010110110: data <= 32'h40a8bca6;
    11'b00010110111: data <= 32'h3f4db9ba;
    11'b00010111000: data <= 32'h35ccb830;
    11'b00010111001: data <= 32'h2fd4b6a3;
    11'b00010111010: data <= 32'h3bde346e;
    11'b00010111011: data <= 32'h3b513b19;
    11'b00010111100: data <= 32'hb9912d60;
    11'b00010111101: data <= 32'hc01abed7;
    11'b00010111110: data <= 32'hbeabc0b4;
    11'b00010111111: data <= 32'hb63dbbe1;
    11'b00011000000: data <= 32'h32b238a0;
    11'b00011000001: data <= 32'h2dec380a;
    11'b00011000010: data <= 32'h2f62b562;
    11'b00011000011: data <= 32'h2f80305b;
    11'b00011000100: data <= 32'hb9583f52;
    11'b00011000101: data <= 32'hbec340fb;
    11'b00011000110: data <= 32'hbd903c52;
    11'b00011000111: data <= 32'h34e5b9ae;
    11'b00011001000: data <= 32'h3df2bbea;
    11'b00011001001: data <= 32'h3bfeb009;
    11'b00011001010: data <= 32'h3340364b;
    11'b00011001011: data <= 32'h3b0c35be;
    11'b00011001100: data <= 32'h4049386d;
    11'b00011001101: data <= 32'h3f1d3a6e;
    11'b00011001110: data <= 32'hb5d82f19;
    11'b00011001111: data <= 32'hbf90bd3e;
    11'b00011010000: data <= 32'hbcdbbf8c;
    11'b00011010001: data <= 32'h35f5bc4b;
    11'b00011010010: data <= 32'h3abbb5b1;
    11'b00011010011: data <= 32'h3224bb00;
    11'b00011010100: data <= 32'hb3debdac;
    11'b00011010101: data <= 32'hb3d4b423;
    11'b00011010110: data <= 32'hb9893f5e;
    11'b00011010111: data <= 32'hbe3540b8;
    11'b00011011000: data <= 32'hbe893912;
    11'b00011011001: data <= 32'hb940bc68;
    11'b00011011010: data <= 32'h2e27baef;
    11'b00011011011: data <= 32'hae943823;
    11'b00011011100: data <= 32'hadff3c66;
    11'b00011011101: data <= 32'h3cae39a6;
    11'b00011011110: data <= 32'h40e738e7;
    11'b00011011111: data <= 32'h3f053c41;
    11'b00011100000: data <= 32'hb7a13b8a;
    11'b00011100001: data <= 32'hbe65ae97;
    11'b00011100010: data <= 32'hb64ebba6;
    11'b00011100011: data <= 32'h3d36bb9d;
    11'b00011100100: data <= 32'h3d7ebbb4;
    11'b00011100101: data <= 32'h3484be81;
    11'b00011100110: data <= 32'hb09bbf4d;
    11'b00011100111: data <= 32'h34d3b668;
    11'b00011101000: data <= 32'h326b3df8;
    11'b00011101001: data <= 32'hbb3f3e30;
    11'b00011101010: data <= 32'hbf1ab548;
    11'b00011101011: data <= 32'hbe3ebea8;
    11'b00011101100: data <= 32'hbc06bacf;
    11'b00011101101: data <= 32'hbaa739b5;
    11'b00011101110: data <= 32'hb6333bb0;
    11'b00011101111: data <= 32'h3b2c3249;
    11'b00011110000: data <= 32'h3f5f3423;
    11'b00011110001: data <= 32'h3bc33db7;
    11'b00011110010: data <= 32'hbb52401c;
    11'b00011110011: data <= 32'hbd9a3ccf;
    11'b00011110100: data <= 32'h30a2ad51;
    11'b00011110101: data <= 32'h3e70b958;
    11'b00011110110: data <= 32'h3cfebb38;
    11'b00011110111: data <= 32'h30b1bd78;
    11'b00011111000: data <= 32'h34eebd85;
    11'b00011111001: data <= 32'h3dd6b280;
    11'b00011111010: data <= 32'h3e293c5e;
    11'b00011111011: data <= 32'hac4139d3;
    11'b00011111100: data <= 32'hbeaabc04;
    11'b00011111101: data <= 32'hbf56bf65;
    11'b00011111110: data <= 32'hbcb1ba92;
    11'b00011111111: data <= 32'hba4035a9;
    11'b00100000000: data <= 32'hb75ea89b;
    11'b00100000001: data <= 32'h3563bc02;
    11'b00100000010: data <= 32'h3b00b6b8;
    11'b00100000011: data <= 32'h2e913e5e;
    11'b00100000100: data <= 32'hbd094174;
    11'b00100000101: data <= 32'hbd653f39;
    11'b00100000110: data <= 32'h27a232e3;
    11'b00100000111: data <= 32'h3ba9b67d;
    11'b00100001000: data <= 32'h3583b4b8;
    11'b00100001001: data <= 32'hb4ddb69e;
    11'b00100001010: data <= 32'h39deb82b;
    11'b00100001011: data <= 32'h40fa2f3d;
    11'b00100001100: data <= 32'h41083b21;
    11'b00100001101: data <= 32'h37903815;
    11'b00100001110: data <= 32'hbd7aba52;
    11'b00100001111: data <= 32'hbd68bd4b;
    11'b00100010000: data <= 32'hb675b8db;
    11'b00100010001: data <= 32'hae5fb3ae;
    11'b00100010010: data <= 32'hb52cbd1a;
    11'b00100010011: data <= 32'haee4c06a;
    11'b00100010100: data <= 32'h34dbbc42;
    11'b00100010101: data <= 32'hae943dad;
    11'b00100010110: data <= 32'hbc58411a;
    11'b00100010111: data <= 32'hbd413d84;
    11'b00100011000: data <= 32'hb8c2b1e1;
    11'b00100011001: data <= 32'hb48cb4e4;
    11'b00100011010: data <= 32'hbb1e3685;
    11'b00100011011: data <= 32'hbb48377e;
    11'b00100011100: data <= 32'h3a6210b1;
    11'b00100011101: data <= 32'h417a3146;
    11'b00100011110: data <= 32'h41153b3f;
    11'b00100011111: data <= 32'h36683c10;
    11'b00100100000: data <= 32'hbc4b342c;
    11'b00100100001: data <= 32'hb7c9b429;
    11'b00100100010: data <= 32'h395bb193;
    11'b00100100011: data <= 32'h38c2b8b2;
    11'b00100100100: data <= 32'hb2f2bfd4;
    11'b00100100101: data <= 32'hb2d6c163;
    11'b00100100110: data <= 32'h3854bd31;
    11'b00100100111: data <= 32'h38fd3c21;
    11'b00100101000: data <= 32'hb5173ecd;
    11'b00100101001: data <= 32'hbc8534db;
    11'b00100101010: data <= 32'hbcd8bb1d;
    11'b00100101011: data <= 32'hbd3bb526;
    11'b00100101100: data <= 32'hbee93a34;
    11'b00100101101: data <= 32'hbd6538eb;
    11'b00100101110: data <= 32'h3726b55c;
    11'b00100101111: data <= 32'h402fb4a9;
    11'b00100110000: data <= 32'h3eb53b99;
    11'b00100110001: data <= 32'hb0f83f49;
    11'b00100110010: data <= 32'hbb4f3de9;
    11'b00100110011: data <= 32'h322d39fa;
    11'b00100110100: data <= 32'h3cf434f1;
    11'b00100110101: data <= 32'h3933b682;
    11'b00100110110: data <= 32'hb6dbbea5;
    11'b00100110111: data <= 32'hac4dc069;
    11'b00100111000: data <= 32'h3d8abc12;
    11'b00100111001: data <= 32'h3f753957;
    11'b00100111010: data <= 32'h39633a1e;
    11'b00100111011: data <= 32'hba34b8e3;
    11'b00100111100: data <= 32'hbd4abd0a;
    11'b00100111101: data <= 32'hbdbfb3cf;
    11'b00100111110: data <= 32'hbeb33995;
    11'b00100111111: data <= 32'hbd8aac56;
    11'b00101000000: data <= 32'hadccbdb1;
    11'b00101000001: data <= 32'h3c1ebc83;
    11'b00101000010: data <= 32'h38bc3aa6;
    11'b00101000011: data <= 32'hb9814096;
    11'b00101000100: data <= 32'hbabb4014;
    11'b00101000101: data <= 32'h35573c58;
    11'b00101000110: data <= 32'h3b2d38b7;
    11'b00101000111: data <= 32'hb02e327a;
    11'b00101001000: data <= 32'hbc23b908;
    11'b00101001001: data <= 32'h2b1bbca0;
    11'b00101001010: data <= 32'h405fb822;
    11'b00101001011: data <= 32'h4198378a;
    11'b00101001100: data <= 32'h3d2c3518;
    11'b00101001101: data <= 32'hb66db9a0;
    11'b00101001110: data <= 32'hba73baff;
    11'b00101001111: data <= 32'hb8d02f37;
    11'b00101010000: data <= 32'hbab436a9;
    11'b00101010001: data <= 32'hbc50bc3a;
    11'b00101010010: data <= 32'hb81bc12b;
    11'b00101010011: data <= 32'h341bbf8f;
    11'b00101010100: data <= 32'h2d8c3835;
    11'b00101010101: data <= 32'hb9664018;
    11'b00101010110: data <= 32'hb97b3e3c;
    11'b00101010111: data <= 32'h25723895;
    11'b00101011000: data <= 32'had013864;
    11'b00101011001: data <= 32'hbd443b03;
    11'b00101011010: data <= 32'hbf2536da;
    11'b00101011011: data <= 32'hac10b584;
    11'b00101011100: data <= 32'h40a9b491;
    11'b00101011101: data <= 32'h418d3649;
    11'b00101011110: data <= 32'h3c9b3828;
    11'b00101011111: data <= 32'hb2942c57;
    11'b00101100000: data <= 32'h28b83039;
    11'b00101100001: data <= 32'h38ff39b2;
    11'b00101100010: data <= 32'h303234b8;
    11'b00101100011: data <= 32'hba3abe6a;
    11'b00101100100: data <= 32'hb972c212;
    11'b00101100101: data <= 32'h3296c033;
    11'b00101100110: data <= 32'h382a3212;
    11'b00101100111: data <= 32'h25143cd0;
    11'b00101101000: data <= 32'hb53c3591;
    11'b00101101001: data <= 32'hb55db630;
    11'b00101101010: data <= 32'hbb863556;
    11'b00101101011: data <= 32'hc0443d1d;
    11'b00101101100: data <= 32'hc0823ac2;
    11'b00101101101: data <= 32'hb6a9b60e;
    11'b00101101110: data <= 32'h3eb0b928;
    11'b00101101111: data <= 32'h3f2f3447;
    11'b00101110000: data <= 32'h35e83c2c;
    11'b00101110001: data <= 32'hb3a23c65;
    11'b00101110010: data <= 32'h39da3c82;
    11'b00101110011: data <= 32'h3dc73d17;
    11'b00101110100: data <= 32'h37eb3842;
    11'b00101110101: data <= 32'hbaedbd18;
    11'b00101110110: data <= 32'hb97fc0e7;
    11'b00101110111: data <= 32'h3a0abe86;
    11'b00101111000: data <= 32'h3e3516db;
    11'b00101111001: data <= 32'h3c023438;
    11'b00101111010: data <= 32'h30bbba68;
    11'b00101111011: data <= 32'hb560bc47;
    11'b00101111100: data <= 32'hbc0d3430;
    11'b00101111101: data <= 32'hc0043d53;
    11'b00101111110: data <= 32'hc04a3759;
    11'b00101111111: data <= 32'hba71bcf2;
    11'b00110000000: data <= 32'h38debddd;
    11'b00110000001: data <= 32'h37de963e;
    11'b00110000010: data <= 32'hb79f3d6c;
    11'b00110000011: data <= 32'hb56b3e53;
    11'b00110000100: data <= 32'h3bd33dae;
    11'b00110000101: data <= 32'h3d983dd9;
    11'b00110000110: data <= 32'ha89f3c20;
    11'b00110000111: data <= 32'hbdc5b3a9;
    11'b00110001000: data <= 32'hb9d9bccf;
    11'b00110001001: data <= 32'h3d6eba97;
    11'b00110001010: data <= 32'h40c49d5f;
    11'b00110001011: data <= 32'h3e65b440;
    11'b00110001100: data <= 32'h37cebcbe;
    11'b00110001101: data <= 32'h2f9ebba3;
    11'b00110001110: data <= 32'hb163388d;
    11'b00110001111: data <= 32'hbbf73ce2;
    11'b00110010000: data <= 32'hbe34b4da;
    11'b00110010001: data <= 32'hbc1fc08d;
    11'b00110010010: data <= 32'hb34cc072;
    11'b00110010011: data <= 32'hb4dcb53a;
    11'b00110010100: data <= 32'hba0c3c7b;
    11'b00110010101: data <= 32'hb4233c50;
    11'b00110010110: data <= 32'h3aac3a12;
    11'b00110010111: data <= 32'h39603caa;
    11'b00110011000: data <= 32'hbc513e0e;
    11'b00110011001: data <= 32'hc0683aec;
    11'b00110011010: data <= 32'hbb57aed6;
    11'b00110011011: data <= 32'h3ddbb475;
    11'b00110011100: data <= 32'h40a82613;
    11'b00110011101: data <= 32'h3d5bb31c;
    11'b00110011110: data <= 32'h378bb974;
    11'b00110011111: data <= 32'h3a50af40;
    11'b00110100000: data <= 32'h3c623cba;
    11'b00110100001: data <= 32'h33e93cd3;
    11'b00110100010: data <= 32'hbb61ba26;
    11'b00110100011: data <= 32'hbc3dc15d;
    11'b00110100100: data <= 32'hb6bbc0b3;
    11'b00110100101: data <= 32'hb0dbb802;
    11'b00110100110: data <= 32'hb41136b6;
    11'b00110100111: data <= 32'h2ee8b14a;
    11'b00110101000: data <= 32'h38e8b758;
    11'b00110101001: data <= 32'hac7538f5;
    11'b00110101010: data <= 32'hbf5f3f03;
    11'b00110101011: data <= 32'hc13d3d9f;
    11'b00110101100: data <= 32'hbca630ef;
    11'b00110101101: data <= 32'h3b4eb697;
    11'b00110101110: data <= 32'h3d42adfd;
    11'b00110101111: data <= 32'h351b30ab;
    11'b00110110000: data <= 32'h2f673230;
    11'b00110110001: data <= 32'h3d3a3a8c;
    11'b00110110010: data <= 32'h400c3ee7;
    11'b00110110011: data <= 32'h3b513d91;
    11'b00110110100: data <= 32'hba03b811;
    11'b00110110101: data <= 32'hbc20c021;
    11'b00110110110: data <= 32'ha85bbeab;
    11'b00110110111: data <= 32'h3989b62f;
    11'b00110111000: data <= 32'h392db577;
    11'b00110111001: data <= 32'h38bbbda5;
    11'b00110111010: data <= 32'h38e9bdcf;
    11'b00110111011: data <= 32'hb1883424;
    11'b00110111100: data <= 32'hbec23ef6;
    11'b00110111101: data <= 32'hc0ab3cba;
    11'b00110111110: data <= 32'hbd1fb7cf;
    11'b00110111111: data <= 32'h2574bc84;
    11'b00111000000: data <= 32'had04b629;
    11'b00111000001: data <= 32'hbab83691;
    11'b00111000010: data <= 32'hb4c53956;
    11'b00111000011: data <= 32'h3dd73c58;
    11'b00111000100: data <= 32'h40453f1e;
    11'b00111000101: data <= 32'h39003ea6;
    11'b00111000110: data <= 32'hbcc735e9;
    11'b00111000111: data <= 32'hbc65b9e3;
    11'b00111001000: data <= 32'h37bfb866;
    11'b00111001001: data <= 32'h3de8abf9;
    11'b00111001010: data <= 32'h3ce1ba06;
    11'b00111001011: data <= 32'h3ab7bfcc;
    11'b00111001100: data <= 32'h3b22be6a;
    11'b00111001101: data <= 32'h384a3661;
    11'b00111001110: data <= 32'hb8d83e95;
    11'b00111001111: data <= 32'hbdc6383c;
    11'b00111010000: data <= 32'hbcabbdc9;
    11'b00111010001: data <= 32'hb96cbf70;
    11'b00111010010: data <= 32'hbc17b944;
    11'b00111010011: data <= 32'hbda634c5;
    11'b00111010100: data <= 32'hb6c4345f;
    11'b00111010101: data <= 32'h3d4135d9;
    11'b00111010110: data <= 32'h3e253cd9;
    11'b00111010111: data <= 32'hb4e53f41;
    11'b00111011000: data <= 32'hbfad3d4d;
    11'b00111011001: data <= 32'hbd10380a;
    11'b00111011010: data <= 32'h394b34fc;
    11'b00111011011: data <= 32'h3e0232c0;
    11'b00111011100: data <= 32'h3b52b97d;
    11'b00111011101: data <= 32'h38b3be59;
    11'b00111011110: data <= 32'h3d03bb42;
    11'b00111011111: data <= 32'h3e983bb2;
    11'b00111100000: data <= 32'h3a353e8a;
    11'b00111100001: data <= 32'hb7b228cc;
    11'b00111100010: data <= 32'hbb53bf9e;
    11'b00111100011: data <= 32'hba94bfd0;
    11'b00111100100: data <= 32'hbc1ab91c;
    11'b00111100101: data <= 32'hbc5eb020;
    11'b00111100110: data <= 32'hb02aba99;
    11'b00111100111: data <= 32'h3c72bbdc;
    11'b00111101000: data <= 32'h3a743532;
    11'b00111101001: data <= 32'hbc603ef9;
    11'b00111101010: data <= 32'hc0a23f2b;
    11'b00111101011: data <= 32'hbd713b70;
    11'b00111101100: data <= 32'h35823664;
    11'b00111101101: data <= 32'h38f93271;
    11'b00111101110: data <= 32'hb330b56e;
    11'b00111101111: data <= 32'hae9cba12;
    11'b00111110000: data <= 32'h3dc92593;
    11'b00111110001: data <= 32'h40f73dfc;
    11'b00111110010: data <= 32'h3e743edb;
    11'b00111110011: data <= 32'haa542ee1;
    11'b00111110100: data <= 32'hb9e7bda3;
    11'b00111110101: data <= 32'hb734bcaa;
    11'b00111110110: data <= 32'hb423b292;
    11'b00111110111: data <= 32'hb32eb87f;
    11'b00111111000: data <= 32'h3595bfdd;
    11'b00111111001: data <= 32'h3c30c04d;
    11'b00111111010: data <= 32'h3874b54d;
    11'b00111111011: data <= 32'hbc333e27;
    11'b00111111100: data <= 32'hbfc93e46;
    11'b00111111101: data <= 32'hbcbf363d;
    11'b00111111110: data <= 32'hb355b3e6;
    11'b00111111111: data <= 32'hb94aad08;
    11'b01000000000: data <= 32'hbe40a986;
    11'b01000000001: data <= 32'hbabbb1cb;
    11'b01000000010: data <= 32'h3d78362a;
    11'b01000000011: data <= 32'h41273df7;
    11'b01000000100: data <= 32'h3dcc3eeb;
    11'b01000000101: data <= 32'hb614397a;
    11'b01000000110: data <= 32'hba33b223;
    11'b01000000111: data <= 32'h2cf5302e;
    11'b01000001000: data <= 32'h38b6376b;
    11'b01000001001: data <= 32'h36dbb9ad;
    11'b01000001010: data <= 32'h3882c0f1;
    11'b01000001011: data <= 32'h3c74c0e6;
    11'b01000001100: data <= 32'h3befb593;
    11'b01000001101: data <= 32'had1c3d88;
    11'b01000001110: data <= 32'hbb133b57;
    11'b01000001111: data <= 32'hb9c1b8c3;
    11'b01000010000: data <= 32'hb91ebc25;
    11'b01000010001: data <= 32'hbe3fb56f;
    11'b01000010010: data <= 32'hc09c20ce;
    11'b01000010011: data <= 32'hbcadb557;
    11'b01000010100: data <= 32'h3c81b307;
    11'b01000010101: data <= 32'h3fee3a2a;
    11'b01000010110: data <= 32'h38303e1f;
    11'b01000010111: data <= 32'hbc8d3d59;
    11'b01000011000: data <= 32'hbb883bf8;
    11'b01000011001: data <= 32'h360d3cbb;
    11'b01000011010: data <= 32'h3a913be6;
    11'b01000011011: data <= 32'h33a3b811;
    11'b01000011100: data <= 32'h31e3c03a;
    11'b01000011101: data <= 32'h3c93bf2a;
    11'b01000011110: data <= 32'h3f2f32f3;
    11'b01000011111: data <= 32'h3cf53d7f;
    11'b01000100000: data <= 32'h348e3564;
    11'b01000100001: data <= 32'hb18dbce7;
    11'b01000100010: data <= 32'hb8e2bcf9;
    11'b01000100011: data <= 32'hbe43b314;
    11'b01000100100: data <= 32'hc01daf7b;
    11'b01000100101: data <= 32'hbb4dbc86;
    11'b01000100110: data <= 32'h3b57bdfd;
    11'b01000100111: data <= 32'h3cc4b548;
    11'b01000101000: data <= 32'hb67a3c87;
    11'b01000101001: data <= 32'hbe963e5f;
    11'b01000101010: data <= 32'hbbbc3dac;
    11'b01000101011: data <= 32'h35323d87;
    11'b01000101100: data <= 32'h33413c3e;
    11'b01000101101: data <= 32'hba97b06b;
    11'b01000101110: data <= 32'hb9bcbcfa;
    11'b01000101111: data <= 32'h3beaba06;
    11'b01000110000: data <= 32'h40c83ad8;
    11'b01000110001: data <= 32'h40233da5;
    11'b01000110010: data <= 32'h3ae931c6;
    11'b01000110011: data <= 32'h3089bbfc;
    11'b01000110100: data <= 32'hb1fab854;
    11'b01000110101: data <= 32'hba31368d;
    11'b01000110110: data <= 32'hbc76b250;
    11'b01000110111: data <= 32'hb57fc006;
    11'b01000111000: data <= 32'h3aacc14f;
    11'b01000111001: data <= 32'h3a05bcaa;
    11'b01000111010: data <= 32'hb8e139e1;
    11'b01000111011: data <= 32'hbd7c3d21;
    11'b01000111100: data <= 32'hb8ed3aeb;
    11'b01000111101: data <= 32'h2e47399b;
    11'b01000111110: data <= 32'hba4b39ba;
    11'b01000111111: data <= 32'hc04b3133;
    11'b01001000000: data <= 32'hbea5b819;
    11'b01001000001: data <= 32'h395ab119;
    11'b01001000010: data <= 32'h40b93bac;
    11'b01001000011: data <= 32'h3f993d1d;
    11'b01001000100: data <= 32'h385436d4;
    11'b01001000101: data <= 32'h2cdaab0a;
    11'b01001000110: data <= 32'h357d39e4;
    11'b01001000111: data <= 32'h32473d38;
    11'b01001001000: data <= 32'hb416ac00;
    11'b01001001001: data <= 32'h9fbbc0ba;
    11'b01001001010: data <= 32'h3a4ac1e8;
    11'b01001001011: data <= 32'h3b0abcf2;
    11'b01001001100: data <= 32'h2d663881;
    11'b01001001101: data <= 32'hb56538f5;
    11'b01001001110: data <= 32'h2d93b2f2;
    11'b01001001111: data <= 32'h0dfab44e;
    11'b01001010000: data <= 32'hbe073542;
    11'b01001010001: data <= 32'hc1cc34ba;
    11'b01001010010: data <= 32'hc02db631;
    11'b01001010011: data <= 32'h35c2b7d6;
    11'b01001010100: data <= 32'h3ef23484;
    11'b01001010101: data <= 32'h3b303ac7;
    11'b01001010110: data <= 32'hb5dd39f7;
    11'b01001010111: data <= 32'hb2c73b74;
    11'b01001011000: data <= 32'h39923f3d;
    11'b01001011001: data <= 32'h39653fe3;
    11'b01001011010: data <= 32'hb19e3424;
    11'b01001011011: data <= 32'hb52bbfcf;
    11'b01001011100: data <= 32'h38cec07a;
    11'b01001011101: data <= 32'h3d5fb875;
    11'b01001011110: data <= 32'h3cbd3946;
    11'b01001011111: data <= 32'h3add1cb6;
    11'b01001100000: data <= 32'h3a8cbc42;
    11'b01001100001: data <= 32'h327cb9e7;
    11'b01001100010: data <= 32'hbdbc35c5;
    11'b01001100011: data <= 32'hc13c35be;
    11'b01001100100: data <= 32'hbf0bbac7;
    11'b01001100101: data <= 32'h3366be23;
    11'b01001100110: data <= 32'h3b5cbabf;
    11'b01001100111: data <= 32'hb3183361;
    11'b01001101000: data <= 32'hbc813a3e;
    11'b01001101001: data <= 32'hb57e3d03;
    11'b01001101010: data <= 32'h3a6b3ffb;
    11'b01001101011: data <= 32'h367a400d;
    11'b01001101100: data <= 32'hbbf438ae;
    11'b01001101101: data <= 32'hbcf5bc3b;
    11'b01001101110: data <= 32'h32acbc22;
    11'b01001101111: data <= 32'h3eb5351e;
    11'b01001110000: data <= 32'h3f913a8a;
    11'b01001110001: data <= 32'h3dcbb481;
    11'b01001110010: data <= 32'h3cadbc95;
    11'b01001110011: data <= 32'h3905b49e;
    11'b01001110100: data <= 32'hb8e73bf0;
    11'b01001110101: data <= 32'hbe22382b;
    11'b01001110110: data <= 32'hbbc8bdc2;
    11'b01001110111: data <= 32'h346ec118;
    11'b01001111000: data <= 32'h360abed7;
    11'b01001111001: data <= 32'hb9c0b41f;
    11'b01001111010: data <= 32'hbc7336ab;
    11'b01001111011: data <= 32'ha22d3948;
    11'b01001111100: data <= 32'h3a7f3ccf;
    11'b01001111101: data <= 32'hb4d73df9;
    11'b01001111110: data <= 32'hc0503a12;
    11'b01001111111: data <= 32'hc075b3df;
    11'b01010000000: data <= 32'hb40ab146;
    11'b01010000001: data <= 32'h3e2c398e;
    11'b01010000010: data <= 32'h3eac39d7;
    11'b01010000011: data <= 32'h3c2db41e;
    11'b01010000100: data <= 32'h3bacb823;
    11'b01010000101: data <= 32'h3c2f3a82;
    11'b01010000110: data <= 32'h36bb3fc3;
    11'b01010000111: data <= 32'hb6ab3ab2;
    11'b01010001000: data <= 32'hb5bebe8e;
    11'b01010001001: data <= 32'h34d8c18f;
    11'b01010001010: data <= 32'h34dcbeec;
    11'b01010001011: data <= 32'hb580b562;
    11'b01010001100: data <= 32'hb455b139;
    11'b01010001101: data <= 32'h39f5b79c;
    11'b01010001110: data <= 32'h3b69976f;
    11'b01010001111: data <= 32'hbaa73aa1;
    11'b01010010000: data <= 32'hc1a93a57;
    11'b01010010001: data <= 32'hc1472b28;
    11'b01010010010: data <= 32'hb831b198;
    11'b01010010011: data <= 32'h3bb3335f;
    11'b01010010100: data <= 32'h38eb3412;
    11'b01010010101: data <= 32'hac9fb171;
    11'b01010010110: data <= 32'h367f33db;
    11'b01010010111: data <= 32'h3d213f30;
    11'b01010011000: data <= 32'h3c33413f;
    11'b01010011001: data <= 32'ha4ec3cb6;
    11'b01010011010: data <= 32'hb704bceb;
    11'b01010011011: data <= 32'h2dfec006;
    11'b01010011100: data <= 32'h3839baf8;
    11'b01010011101: data <= 32'h380a16fc;
    11'b01010011110: data <= 32'h3a97b941;
    11'b01010011111: data <= 32'h3e15bdd0;
    11'b01010100000: data <= 32'h3cd0ba43;
    11'b01010100001: data <= 32'hb9c238d3;
    11'b01010100010: data <= 32'hc0fd3ad0;
    11'b01010100011: data <= 32'hc054b169;
    11'b01010100100: data <= 32'hb71cbb92;
    11'b01010100101: data <= 32'h342bba3b;
    11'b01010100110: data <= 32'hb8f6b6d7;
    11'b01010100111: data <= 32'hbc8bb42d;
    11'b01010101000: data <= 32'h8a3e37ca;
    11'b01010101001: data <= 32'h3d6b3fba;
    11'b01010101010: data <= 32'h3c044124;
    11'b01010101011: data <= 32'hb8623d5b;
    11'b01010101100: data <= 32'hbcdeb6f9;
    11'b01010101101: data <= 32'hb5f4b99e;
    11'b01010101110: data <= 32'h398d34c7;
    11'b01010101111: data <= 32'h3c5f3720;
    11'b01010110000: data <= 32'h3d75bb10;
    11'b01010110001: data <= 32'h3f3ebef8;
    11'b01010110010: data <= 32'h3e10b917;
    11'b01010110011: data <= 32'h26593c49;
    11'b01010110100: data <= 32'hbd453c54;
    11'b01010110101: data <= 32'hbc67b886;
    11'b01010110110: data <= 32'haf0dbf38;
    11'b01010110111: data <= 32'hb270be60;
    11'b01010111000: data <= 32'hbd40bb30;
    11'b01010111001: data <= 32'hbdc0b890;
    11'b01010111010: data <= 32'h307fab94;
    11'b01010111011: data <= 32'h3dad3c39;
    11'b01010111100: data <= 32'h38123f27;
    11'b01010111101: data <= 32'hbe1b3cee;
    11'b01010111110: data <= 32'hc04d3484;
    11'b01010111111: data <= 32'hbad53599;
    11'b01011000000: data <= 32'h38733c00;
    11'b01011000001: data <= 32'h3b0e38a0;
    11'b01011000010: data <= 32'h3b1ebb25;
    11'b01011000011: data <= 32'h3d8cbd57;
    11'b01011000100: data <= 32'h3eb63417;
    11'b01011000101: data <= 32'h3bad3fd0;
    11'b01011000110: data <= 32'ha7733dcb;
    11'b01011000111: data <= 32'hb0deb9ac;
    11'b01011001000: data <= 32'h314ac008;
    11'b01011001001: data <= 32'hb491be39;
    11'b01011001010: data <= 32'hbca6ba79;
    11'b01011001011: data <= 32'hbaa6bb72;
    11'b01011001100: data <= 32'h3a86bc67;
    11'b01011001101: data <= 32'h3e68b4e5;
    11'b01011001110: data <= 32'h2d0b3a4e;
    11'b01011001111: data <= 32'hc04b3bf0;
    11'b01011010000: data <= 32'hc106388d;
    11'b01011010001: data <= 32'hbc053887;
    11'b01011010010: data <= 32'h30c73a64;
    11'b01011010011: data <= 32'hadc932a9;
    11'b01011010100: data <= 32'hb5eebb0f;
    11'b01011010101: data <= 32'h3810b9a8;
    11'b01011010110: data <= 32'h3e803ca2;
    11'b01011010111: data <= 32'h3e334133;
    11'b01011011000: data <= 32'h38be3ede;
    11'b01011011001: data <= 32'h2bb7b6c6;
    11'b01011011010: data <= 32'h2dfebd3d;
    11'b01011011011: data <= 32'hb057b88b;
    11'b01011011100: data <= 32'hb7a2b14a;
    11'b01011011101: data <= 32'h30fbbc89;
    11'b01011011110: data <= 32'h3e41c00b;
    11'b01011011111: data <= 32'h3f68bd3b;
    11'b01011100000: data <= 32'h2f9533d3;
    11'b01011100001: data <= 32'hbf6a3b03;
    11'b01011100010: data <= 32'hbfb6367c;
    11'b01011100011: data <= 32'hb933a4ca;
    11'b01011100100: data <= 32'hb469ac94;
    11'b01011100101: data <= 32'hbd0cb726;
    11'b01011100110: data <= 32'hbe9abbe4;
    11'b01011100111: data <= 32'hb392b714;
    11'b01011101000: data <= 32'h3df23d45;
    11'b01011101001: data <= 32'h3e2e40eb;
    11'b01011101010: data <= 32'h344a3e91;
    11'b01011101011: data <= 32'hb85f2f8c;
    11'b01011101100: data <= 32'hb55bac1a;
    11'b01011101101: data <= 32'ha2943a80;
    11'b01011101110: data <= 32'h2d9f390a;
    11'b01011101111: data <= 32'h399bbc7a;
    11'b01011110000: data <= 32'h3f29c0ab;
    11'b01011110001: data <= 32'h3fe7bd82;
    11'b01011110010: data <= 32'h3923380a;
    11'b01011110011: data <= 32'hb9e63c31;
    11'b01011110100: data <= 32'hb94d2c79;
    11'b01011110101: data <= 32'h291dba82;
    11'b01011110110: data <= 32'hb79bbaf7;
    11'b01011110111: data <= 32'hbfd7bb09;
    11'b01011111000: data <= 32'hc05cbca3;
    11'b01011111001: data <= 32'hb572ba74;
    11'b01011111010: data <= 32'h3dd937fc;
    11'b01011111011: data <= 32'h3c783df7;
    11'b01011111100: data <= 32'hb8e63cbf;
    11'b01011111101: data <= 32'hbdc0387f;
    11'b01011111110: data <= 32'hba5d3bda;
    11'b01011111111: data <= 32'hac2b3f04;
    11'b01100000000: data <= 32'h23d83c2d;
    11'b01100000001: data <= 32'h3476bc07;
    11'b01100000010: data <= 32'h3cd3bff7;
    11'b01100000011: data <= 32'h3f3cb8e7;
    11'b01100000100: data <= 32'h3d343d45;
    11'b01100000101: data <= 32'h38473d9b;
    11'b01100000110: data <= 32'h384baf59;
    11'b01100000111: data <= 32'h390dbc79;
    11'b01100001000: data <= 32'hb66dbb06;
    11'b01100001001: data <= 32'hbf7ab947;
    11'b01100001010: data <= 32'hbeeabce8;
    11'b01100001011: data <= 32'h337dbe55;
    11'b01100001100: data <= 32'h3e85bab8;
    11'b01100001101: data <= 32'h39713397;
    11'b01100001110: data <= 32'hbd2538cd;
    11'b01100001111: data <= 32'hbf5a393f;
    11'b01100010000: data <= 32'hbaca3cff;
    11'b01100010001: data <= 32'hb3253ef2;
    11'b01100010010: data <= 32'hb9b53a7e;
    11'b01100010011: data <= 32'hbba0bbc5;
    11'b01100010100: data <= 32'h2d03bd87;
    11'b01100010101: data <= 32'h3d9334ed;
    11'b01100010110: data <= 32'h3eae3ff9;
    11'b01100010111: data <= 32'h3cce3e68;
    11'b01100011000: data <= 32'h3bb1a7e2;
    11'b01100011001: data <= 32'h39f0b907;
    11'b01100011010: data <= 32'hb2962cff;
    11'b01100011011: data <= 32'hbce23301;
    11'b01100011100: data <= 32'hba12bc42;
    11'b01100011101: data <= 32'h3bfcc087;
    11'b01100011110: data <= 32'h3f5cbf82;
    11'b01100011111: data <= 32'h3885b85d;
    11'b01100100000: data <= 32'hbcb63412;
    11'b01100100001: data <= 32'hbd2736ab;
    11'b01100100010: data <= 32'hb47d39b7;
    11'b01100100011: data <= 32'hb4b53b5b;
    11'b01100100100: data <= 32'hbe8b3120;
    11'b01100100101: data <= 32'hc086bc39;
    11'b01100100110: data <= 32'hbb69bc05;
    11'b01100100111: data <= 32'h3bd638fb;
    11'b01100101000: data <= 32'h3e393f93;
    11'b01100101001: data <= 32'h3b753d5f;
    11'b01100101010: data <= 32'h372631bb;
    11'b01100101011: data <= 32'h358d35eb;
    11'b01100101100: data <= 32'hacbb3def;
    11'b01100101101: data <= 32'hb8ac3d27;
    11'b01100101110: data <= 32'had98b9e5;
    11'b01100101111: data <= 32'h3d18c0dd;
    11'b01100110000: data <= 32'h3f42c003;
    11'b01100110001: data <= 32'h3a4eb6a8;
    11'b01100110010: data <= 32'hb4d635ab;
    11'b01100110011: data <= 32'h9aec2c7e;
    11'b01100110100: data <= 32'h3986af93;
    11'b01100110101: data <= 32'hb0ef2688;
    11'b01100110110: data <= 32'hc053b53a;
    11'b01100110111: data <= 32'hc1b5bc78;
    11'b01100111000: data <= 32'hbccdbc6e;
    11'b01100111001: data <= 32'h3ab32828;
    11'b01100111010: data <= 32'h3c683b52;
    11'b01100111011: data <= 32'h291838e2;
    11'b01100111100: data <= 32'hb80b3448;
    11'b01100111101: data <= 32'hb1503ce7;
    11'b01100111110: data <= 32'haa9740fc;
    11'b01100111111: data <= 32'hb6fb3fa4;
    11'b01101000000: data <= 32'hb4b7b756;
    11'b01101000001: data <= 32'h398dc015;
    11'b01101000010: data <= 32'h3d8bbcff;
    11'b01101000011: data <= 32'h3c5936bd;
    11'b01101000100: data <= 32'h3a2139f9;
    11'b01101000101: data <= 32'h3d12b12d;
    11'b01101000110: data <= 32'h3e1bb8d1;
    11'b01101000111: data <= 32'h3048b1bb;
    11'b01101001000: data <= 32'hc000b021;
    11'b01101001001: data <= 32'hc0dbbb9c;
    11'b01101001010: data <= 32'hb920be22;
    11'b01101001011: data <= 32'h3c17bc5f;
    11'b01101001100: data <= 32'h3912b698;
    11'b01101001101: data <= 32'hba35b404;
    11'b01101001110: data <= 32'hbc542e8d;
    11'b01101001111: data <= 32'hb4223d99;
    11'b01101010000: data <= 32'ha1da4109;
    11'b01101010001: data <= 32'hbaae3ef3;
    11'b01101010010: data <= 32'hbd3db68c;
    11'b01101010011: data <= 32'hb802bda2;
    11'b01101010100: data <= 32'h3969b300;
    11'b01101010101: data <= 32'h3ca23d02;
    11'b01101010110: data <= 32'h3d433c00;
    11'b01101010111: data <= 32'h3f05b3a2;
    11'b01101011000: data <= 32'h3efbb69f;
    11'b01101011001: data <= 32'h361e387b;
    11'b01101011010: data <= 32'hbd4f3a70;
    11'b01101011011: data <= 32'hbd81b7d6;
    11'b01101011100: data <= 32'h341abf8e;
    11'b01101011101: data <= 32'h3d2dbffa;
    11'b01101011110: data <= 32'h3647bd1a;
    11'b01101011111: data <= 32'hbb84ba0e;
    11'b01101100000: data <= 32'hb9fbb394;
    11'b01101100001: data <= 32'h35903aa5;
    11'b01101100010: data <= 32'h32ab3e98;
    11'b01101100011: data <= 32'hbdad3bdc;
    11'b01101100100: data <= 32'hc0eeb873;
    11'b01101100101: data <= 32'hbe66bb7d;
    11'b01101100110: data <= 32'h2ae8356a;
    11'b01101100111: data <= 32'h3b263d75;
    11'b01101101000: data <= 32'h3c0039cc;
    11'b01101101001: data <= 32'h3cdfb4ce;
    11'b01101101010: data <= 32'h3d2433d6;
    11'b01101101011: data <= 32'h37603f35;
    11'b01101101100: data <= 32'hb8f43fe8;
    11'b01101101101: data <= 32'hb7db2d83;
    11'b01101101110: data <= 32'h39eebf6f;
    11'b01101101111: data <= 32'h3d1bc01f;
    11'b01101110000: data <= 32'h35ecbc9e;
    11'b01101110001: data <= 32'hb659b921;
    11'b01101110010: data <= 32'h35d8b86c;
    11'b01101110011: data <= 32'h3db2ab48;
    11'b01101110100: data <= 32'h3901388f;
    11'b01101110101: data <= 32'hbed434ae;
    11'b01101110110: data <= 32'hc1f6b935;
    11'b01101110111: data <= 32'hbfa6ba96;
    11'b01101111000: data <= 32'hb00b2c86;
    11'b01101111001: data <= 32'h36f8388b;
    11'b01101111010: data <= 32'h2bd7aeec;
    11'b01101111011: data <= 32'h2f33b80e;
    11'b01101111100: data <= 32'h38ab3aa6;
    11'b01101111101: data <= 32'h36e24171;
    11'b01101111110: data <= 32'hb4a74155;
    11'b01101111111: data <= 32'hb63e3754;
    11'b01110000000: data <= 32'h35aebdb0;
    11'b01110000001: data <= 32'h3a1bbd08;
    11'b01110000010: data <= 32'h35e3b243;
    11'b01110000011: data <= 32'h3615ad53;
    11'b01110000100: data <= 32'h3e27b9c5;
    11'b01110000101: data <= 32'h40b5b985;
    11'b01110000110: data <= 32'h3c3e2cc8;
    11'b01110000111: data <= 32'hbdd33489;
    11'b01110001000: data <= 32'hc103b6c8;
    11'b01110001001: data <= 32'hbd0fbba2;
    11'b01110001010: data <= 32'h321ab9fc;
    11'b01110001011: data <= 32'h2778b937;
    11'b01110001100: data <= 32'hbb06bc59;
    11'b01110001101: data <= 32'hb9e1baf5;
    11'b01110001110: data <= 32'h34633afe;
    11'b01110001111: data <= 32'h38024165;
    11'b01110010000: data <= 32'hb69740e2;
    11'b01110010001: data <= 32'hbc5c36b1;
    11'b01110010010: data <= 32'hb9c1bab1;
    11'b01110010011: data <= 32'hacedafc9;
    11'b01110010100: data <= 32'h32613b14;
    11'b01110010101: data <= 32'h3a133646;
    11'b01110010110: data <= 32'h3fe8ba66;
    11'b01110010111: data <= 32'h4121ba09;
    11'b01110011000: data <= 32'h3d1537f1;
    11'b01110011001: data <= 32'hba773c51;
    11'b01110011010: data <= 32'hbd733161;
    11'b01110011011: data <= 32'hb086bc28;
    11'b01110011100: data <= 32'h3974bdc6;
    11'b01110011101: data <= 32'hb216bddc;
    11'b01110011110: data <= 32'hbd14be82;
    11'b01110011111: data <= 32'hb9babce8;
    11'b01110100000: data <= 32'h39ca34d5;
    11'b01110100001: data <= 32'h3ab83efd;
    11'b01110100010: data <= 32'hb9ad3df4;
    11'b01110100011: data <= 32'hc0062be8;
    11'b01110100100: data <= 32'hbf0fb673;
    11'b01110100101: data <= 32'hba333920;
    11'b01110100110: data <= 32'hb0983d3e;
    11'b01110100111: data <= 32'h368234b0;
    11'b01110101000: data <= 32'h3d7cbbb0;
    11'b01110101001: data <= 32'h3fc5b62b;
    11'b01110101010: data <= 32'h3ca63def;
    11'b01110101011: data <= 32'hb0b84062;
    11'b01110101100: data <= 32'hb4ad3ad0;
    11'b01110101101: data <= 32'h393abb00;
    11'b01110101110: data <= 32'h3ae4bdbf;
    11'b01110101111: data <= 32'hb498bd26;
    11'b01110110000: data <= 32'hbc0cbd93;
    11'b01110110001: data <= 32'h300abd90;
    11'b01110110010: data <= 32'h3eebb850;
    11'b01110110011: data <= 32'h3d8c3807;
    11'b01110110100: data <= 32'hba8a37ee;
    11'b01110110101: data <= 32'hc0d6b400;
    11'b01110110110: data <= 32'hc00fb3c6;
    11'b01110110111: data <= 32'hbb173932;
    11'b01110111000: data <= 32'hb7f23a63;
    11'b01110111001: data <= 32'hb7f4b747;
    11'b01110111010: data <= 32'h2f9abd3b;
    11'b01110111011: data <= 32'h3b9da421;
    11'b01110111100: data <= 32'h3b364087;
    11'b01110111101: data <= 32'h327241b0;
    11'b01110111110: data <= 32'h2cbf3cd1;
    11'b01110111111: data <= 32'h388bb7d8;
    11'b01111000000: data <= 32'h3746b931;
    11'b01111000001: data <= 32'hb6e2b267;
    11'b01111000010: data <= 32'hb7a7b892;
    11'b01111000011: data <= 32'h3c8bbd50;
    11'b01111000100: data <= 32'h4144bcad;
    11'b01111000101: data <= 32'h3f67b3c9;
    11'b01111000110: data <= 32'hb880317a;
    11'b01111000111: data <= 32'hbfbdb108;
    11'b01111001000: data <= 32'hbd17b3c5;
    11'b01111001001: data <= 32'hb56a2df0;
    11'b01111001010: data <= 32'hb97bb37d;
    11'b01111001011: data <= 32'hbdaebda5;
    11'b01111001100: data <= 32'hbbb9bef8;
    11'b01111001101: data <= 32'h350ea7c9;
    11'b01111001110: data <= 32'h3a74406a;
    11'b01111001111: data <= 32'h321f410f;
    11'b01111010000: data <= 32'hb5a23bcc;
    11'b01111010001: data <= 32'hb4b7ae23;
    11'b01111010010: data <= 32'hb5c73778;
    11'b01111010011: data <= 32'hb9a53c69;
    11'b01111010100: data <= 32'hb2903380;
    11'b01111010101: data <= 32'h3e14bcdb;
    11'b01111010110: data <= 32'h418dbd48;
    11'b01111010111: data <= 32'h3fadae5d;
    11'b01111011000: data <= 32'hac7f39d5;
    11'b01111011001: data <= 32'hba77365a;
    11'b01111011010: data <= 32'h2b7ab255;
    11'b01111011011: data <= 32'h37aeb741;
    11'b01111011100: data <= 32'hb988bbc6;
    11'b01111011101: data <= 32'hbf7fbfa4;
    11'b01111011110: data <= 32'hbce6c006;
    11'b01111011111: data <= 32'h3802b7d1;
    11'b01111100000: data <= 32'h3c573d12;
    11'b01111100001: data <= 32'h284f3d8b;
    11'b01111100010: data <= 32'hbc5c34d7;
    11'b01111100011: data <= 32'hbcf82f54;
    11'b01111100100: data <= 32'hbc283d18;
    11'b01111100101: data <= 32'hbc113f39;
    11'b01111100110: data <= 32'hb7df36cc;
    11'b01111100111: data <= 32'h3b55bd25;
    11'b01111101000: data <= 32'h3ff3bc5c;
    11'b01111101001: data <= 32'h3e113967;
    11'b01111101010: data <= 32'h35e33ee0;
    11'b01111101011: data <= 32'h34b13c4c;
    11'b01111101100: data <= 32'h3c85a2e1;
    11'b01111101101: data <= 32'h3bc9b765;
    11'b01111101110: data <= 32'hb95aba49;
    11'b01111101111: data <= 32'hbefbbe29;
    11'b01111110000: data <= 32'hb8eabfad;
    11'b01111110001: data <= 32'h3d70bc79;
    11'b01111110010: data <= 32'h3e86182e;
    11'b01111110011: data <= 32'ha26c2f9a;
    11'b01111110100: data <= 32'hbddbb57d;
    11'b01111110101: data <= 32'hbdf42ff5;
    11'b01111110110: data <= 32'hbc313d99;
    11'b01111110111: data <= 32'hbca43e2d;
    11'b01111111000: data <= 32'hbcd4b0bc;
    11'b01111111001: data <= 32'hb5a1be82;
    11'b01111111010: data <= 32'h39d8ba7f;
    11'b01111111011: data <= 32'h3b463d89;
    11'b01111111100: data <= 32'h385040ae;
    11'b01111111101: data <= 32'h3a1b3d6f;
    11'b01111111110: data <= 32'h3d4032e6;
    11'b01111111111: data <= 32'h3a303177;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    