
module memory_rom_2(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hb882bdf1;
    11'b00000000001: data <= 32'hb506b9fa;
    11'b00000000010: data <= 32'h34a73bda;
    11'b00000000011: data <= 32'hb4cc3f68;
    11'b00000000100: data <= 32'hbe8338f0;
    11'b00000000101: data <= 32'hc017bcd0;
    11'b00000000110: data <= 32'hbd0cbcf1;
    11'b00000000111: data <= 32'hb6d73650;
    11'b00000001000: data <= 32'ha31f3d6e;
    11'b00000001001: data <= 32'h39463941;
    11'b00000001010: data <= 32'h3e4fab5c;
    11'b00000001011: data <= 32'h3de139c5;
    11'b00000001100: data <= 32'haa7a3fd3;
    11'b00000001101: data <= 32'hbcfb3ee2;
    11'b00000001110: data <= 32'hb7ba2e2b;
    11'b00000001111: data <= 32'h3cf0bcb2;
    11'b00000010000: data <= 32'h3e70bd53;
    11'b00000010001: data <= 32'h36febcc5;
    11'b00000010010: data <= 32'hb239bccf;
    11'b00000010011: data <= 32'h3a02b95d;
    11'b00000010100: data <= 32'h3e5c37ec;
    11'b00000010101: data <= 32'h38333b6e;
    11'b00000010110: data <= 32'hbe4bb23a;
    11'b00000010111: data <= 32'hc0e3bdfb;
    11'b00000011000: data <= 32'hbe62bcc2;
    11'b00000011001: data <= 32'hb84331c7;
    11'b00000011010: data <= 32'hb2293851;
    11'b00000011011: data <= 32'h2990b6e2;
    11'b00000011100: data <= 32'h388fb98c;
    11'b00000011101: data <= 32'h38713b80;
    11'b00000011110: data <= 32'hb6bc417f;
    11'b00000011111: data <= 32'hbc8640f6;
    11'b00000100000: data <= 32'hb6b13826;
    11'b00000100001: data <= 32'h3a7ebae2;
    11'b00000100010: data <= 32'h3af5b9d7;
    11'b00000100011: data <= 32'h295eb445;
    11'b00000100100: data <= 32'h33e4b5fa;
    11'b00000100101: data <= 32'h3f61b674;
    11'b00000100110: data <= 32'h415c31f4;
    11'b00000100111: data <= 32'h3c98382d;
    11'b00000101000: data <= 32'hbd24b2a1;
    11'b00000101001: data <= 32'hc018bc8f;
    11'b00000101010: data <= 32'hbb67bc19;
    11'b00000101011: data <= 32'h2c4eb606;
    11'b00000101100: data <= 32'hb08cb967;
    11'b00000101101: data <= 32'hb83dbeb0;
    11'b00000101110: data <= 32'hb1c4bd80;
    11'b00000101111: data <= 32'h31373a83;
    11'b00000110000: data <= 32'hb5f6416e;
    11'b00000110001: data <= 32'hbc6b406e;
    11'b00000110010: data <= 32'hbb9e337c;
    11'b00000110011: data <= 32'hb525b971;
    11'b00000110100: data <= 32'hb4f52cbc;
    11'b00000110101: data <= 32'hb85f3a0b;
    11'b00000110110: data <= 32'h35f9347c;
    11'b00000110111: data <= 32'h407eb4c3;
    11'b00000111000: data <= 32'h41c83083;
    11'b00000111001: data <= 32'h3cd03b09;
    11'b00000111010: data <= 32'hbb89396b;
    11'b00000111011: data <= 32'hbc99b23a;
    11'b00000111100: data <= 32'h32e0b936;
    11'b00000111101: data <= 32'h3aa7ba43;
    11'b00000111110: data <= 32'ha986bde5;
    11'b00000111111: data <= 32'hba17c0a0;
    11'b00001000000: data <= 32'hb0a6bedf;
    11'b00001000001: data <= 32'h398636aa;
    11'b00001000010: data <= 32'h342f3fa8;
    11'b00001000011: data <= 32'hbbe43caf;
    11'b00001000100: data <= 32'hbe6bb78c;
    11'b00001000101: data <= 32'hbd9db938;
    11'b00001000110: data <= 32'hbcee38c4;
    11'b00001000111: data <= 32'hbc2b3c8a;
    11'b00001001000: data <= 32'h2ad430f8;
    11'b00001001001: data <= 32'h3ed8b920;
    11'b00001001010: data <= 32'h4048328e;
    11'b00001001011: data <= 32'h39bc3eac;
    11'b00001001100: data <= 32'hb9c03f8d;
    11'b00001001101: data <= 32'hb55d3a92;
    11'b00001001110: data <= 32'h3bfab1d0;
    11'b00001001111: data <= 32'h3c55b96d;
    11'b00001010000: data <= 32'hb1b8bd47;
    11'b00001010001: data <= 32'hb954bfeb;
    11'b00001010010: data <= 32'h38c9be31;
    11'b00001010011: data <= 32'h3f6ba2d7;
    11'b00001010100: data <= 32'h3cd23b27;
    11'b00001010101: data <= 32'hb98d2f45;
    11'b00001010110: data <= 32'hbf4fbbe1;
    11'b00001010111: data <= 32'hbebbb8de;
    11'b00001011000: data <= 32'hbd4f390f;
    11'b00001011001: data <= 32'hbcb7391a;
    11'b00001011010: data <= 32'hb838ba46;
    11'b00001011011: data <= 32'h38fabd96;
    11'b00001011100: data <= 32'h3c0530ec;
    11'b00001011101: data <= 32'h2ff9407f;
    11'b00001011110: data <= 32'hb90e412d;
    11'b00001011111: data <= 32'ha9d13d17;
    11'b00001100000: data <= 32'h3b2230ba;
    11'b00001100001: data <= 32'h380bad2d;
    11'b00001100010: data <= 32'hb97cb52c;
    11'b00001100011: data <= 32'hb812bbaa;
    11'b00001100100: data <= 32'h3dcfbc46;
    11'b00001100101: data <= 32'h41c2b467;
    11'b00001100110: data <= 32'h3f93349c;
    11'b00001100111: data <= 32'hb54eb2d4;
    11'b00001101000: data <= 32'hbd94ba7e;
    11'b00001101001: data <= 32'hbb99b58f;
    11'b00001101010: data <= 32'hb89035db;
    11'b00001101011: data <= 32'hbb82b50e;
    11'b00001101100: data <= 32'hbc2cbfd1;
    11'b00001101101: data <= 32'hb4d5c05a;
    11'b00001101110: data <= 32'h34e2ae4c;
    11'b00001101111: data <= 32'ha7be4048;
    11'b00001110000: data <= 32'hb8474087;
    11'b00001110001: data <= 32'hb4aa3af8;
    11'b00001110010: data <= 32'h28b2318a;
    11'b00001110011: data <= 32'hb8c23956;
    11'b00001110100: data <= 32'hbd953ad0;
    11'b00001110101: data <= 32'hb8799f8d;
    11'b00001110110: data <= 32'h3efab9ee;
    11'b00001110111: data <= 32'h4214b5c4;
    11'b00001111000: data <= 32'h3f8135e5;
    11'b00001111001: data <= 32'hae3f360a;
    11'b00001111010: data <= 32'hb8532914;
    11'b00001111011: data <= 32'h35353128;
    11'b00001111100: data <= 32'h379831a9;
    11'b00001111101: data <= 32'hb8dcbbc8;
    11'b00001111110: data <= 32'hbd24c11b;
    11'b00001111111: data <= 32'hb838c0fc;
    11'b00010000000: data <= 32'h3837b701;
    11'b00010000001: data <= 32'h37cf3d72;
    11'b00010000010: data <= 32'hb4793c65;
    11'b00010000011: data <= 32'hb993adf9;
    11'b00010000100: data <= 32'hbafea7e8;
    11'b00010000101: data <= 32'hbdee3cb5;
    11'b00010000110: data <= 32'hbfa93de5;
    11'b00010000111: data <= 32'hbb0331d8;
    11'b00010001000: data <= 32'h3cd3bb89;
    11'b00010001001: data <= 32'h405eb6bd;
    11'b00010001010: data <= 32'h3ca33b21;
    11'b00010001011: data <= 32'hae283d90;
    11'b00010001100: data <= 32'h33f33c19;
    11'b00010001101: data <= 32'h3d563997;
    11'b00010001110: data <= 32'h3c30355d;
    11'b00010001111: data <= 32'hb896ba53;
    11'b00010010000: data <= 32'hbd2dc044;
    11'b00010010001: data <= 32'hab5dc043;
    11'b00010010010: data <= 32'h3de0b958;
    11'b00010010011: data <= 32'h3d9535f7;
    11'b00010010100: data <= 32'h2f66b178;
    11'b00010010101: data <= 32'hba7ebb76;
    11'b00010010110: data <= 32'hbc65b1d4;
    11'b00010010111: data <= 32'hbe0d3d2d;
    11'b00010011000: data <= 32'hbfa13d01;
    11'b00010011001: data <= 32'hbd2bb81a;
    11'b00010011010: data <= 32'h30bebe99;
    11'b00010011011: data <= 32'h3accb8c7;
    11'b00010011100: data <= 32'h33bc3d46;
    11'b00010011101: data <= 32'hb3364004;
    11'b00010011110: data <= 32'h38c33db9;
    11'b00010011111: data <= 32'h3e033b83;
    11'b00010100000: data <= 32'h39e33a7f;
    11'b00010100001: data <= 32'hbc0e31d5;
    11'b00010100010: data <= 32'hbd17bb76;
    11'b00010100011: data <= 32'h38dfbd58;
    11'b00010100100: data <= 32'h40c6b998;
    11'b00010100101: data <= 32'h401db44c;
    11'b00010100110: data <= 32'h3716ba2a;
    11'b00010100111: data <= 32'hb72cbc32;
    11'b00010101000: data <= 32'hb604a2a0;
    11'b00010101001: data <= 32'hb8cb3ca7;
    11'b00010101010: data <= 32'hbd803816;
    11'b00010101011: data <= 32'hbe4cbe37;
    11'b00010101100: data <= 32'hba5ac0d4;
    11'b00010101101: data <= 32'hafacbaea;
    11'b00010101110: data <= 32'hb3423cea;
    11'b00010101111: data <= 32'hb4053eb8;
    11'b00010110000: data <= 32'h37a23b2f;
    11'b00010110001: data <= 32'h3b1039ab;
    11'b00010110010: data <= 32'hb2c73d5b;
    11'b00010110011: data <= 32'hbedd3d74;
    11'b00010110100: data <= 32'hbd84347e;
    11'b00010110101: data <= 32'h3af5b967;
    11'b00010110110: data <= 32'h410db907;
    11'b00010110111: data <= 32'h3fbeb4d3;
    11'b00010111000: data <= 32'h3774b6eb;
    11'b00010111001: data <= 32'h32bbb60a;
    11'b00010111010: data <= 32'h3b3437c6;
    11'b00010111011: data <= 32'h39963c42;
    11'b00010111100: data <= 32'hb999aca2;
    11'b00010111101: data <= 32'hbe86c03c;
    11'b00010111110: data <= 32'hbc75c150;
    11'b00010111111: data <= 32'hb14cbc2c;
    11'b00011000000: data <= 32'h2d0538e3;
    11'b00011000001: data <= 32'ha4fb3818;
    11'b00011000010: data <= 32'h31f5b4dd;
    11'b00011000011: data <= 32'h2d5d3122;
    11'b00011000100: data <= 32'hbc353e93;
    11'b00011000101: data <= 32'hc0624020;
    11'b00011000110: data <= 32'hbe5b39ff;
    11'b00011000111: data <= 32'h374cb906;
    11'b00011001000: data <= 32'h3eaab921;
    11'b00011001001: data <= 32'h3c002e14;
    11'b00011001010: data <= 32'h305436ef;
    11'b00011001011: data <= 32'h3a463856;
    11'b00011001100: data <= 32'h3fe53c07;
    11'b00011001101: data <= 32'h3e3c3cae;
    11'b00011001110: data <= 32'hb62426ae;
    11'b00011001111: data <= 32'hbe3ebec5;
    11'b00011010000: data <= 32'hba2ec035;
    11'b00011010001: data <= 32'h38c9bbb8;
    11'b00011010010: data <= 32'h3b2fb141;
    11'b00011010011: data <= 32'h3607ba83;
    11'b00011010100: data <= 32'h2c5cbdc0;
    11'b00011010101: data <= 32'hb1deb4d7;
    11'b00011010110: data <= 32'hbc4f3e99;
    11'b00011010111: data <= 32'hc00e3fdb;
    11'b00011011000: data <= 32'hbeed3429;
    11'b00011011001: data <= 32'hb663bce0;
    11'b00011011010: data <= 32'h3484ba96;
    11'b00011011011: data <= 32'hb2d737bf;
    11'b00011011100: data <= 32'hb5463c36;
    11'b00011011101: data <= 32'h3bee3b8c;
    11'b00011011110: data <= 32'h40853c87;
    11'b00011011111: data <= 32'h3dea3dae;
    11'b00011100000: data <= 32'hb9633a84;
    11'b00011100001: data <= 32'hbe27b733;
    11'b00011100010: data <= 32'hb18fbc13;
    11'b00011100011: data <= 32'h3decb929;
    11'b00011100100: data <= 32'h3e32b923;
    11'b00011100101: data <= 32'h3905be1c;
    11'b00011100110: data <= 32'h341abf3f;
    11'b00011100111: data <= 32'h3619b526;
    11'b00011101000: data <= 32'hb02a3e02;
    11'b00011101001: data <= 32'hbce33d3e;
    11'b00011101010: data <= 32'hbea5b9b1;
    11'b00011101011: data <= 32'hbca4bfdb;
    11'b00011101100: data <= 32'hba60bc30;
    11'b00011101101: data <= 32'hbbbd3823;
    11'b00011101110: data <= 32'hb8af3ad3;
    11'b00011101111: data <= 32'h3aae362e;
    11'b00011110000: data <= 32'h3ef8393c;
    11'b00011110001: data <= 32'h39113e6e;
    11'b00011110010: data <= 32'hbd5e3f39;
    11'b00011110011: data <= 32'hbe813af1;
    11'b00011110100: data <= 32'h3136aa75;
    11'b00011110101: data <= 32'h3edeb4d7;
    11'b00011110110: data <= 32'h3da6b8e2;
    11'b00011110111: data <= 32'h3708bd37;
    11'b00011111000: data <= 32'h38d1bd1d;
    11'b00011111001: data <= 32'h3de12fcb;
    11'b00011111010: data <= 32'h3d0f3d9b;
    11'b00011111011: data <= 32'hb339398c;
    11'b00011111100: data <= 32'hbda3bd61;
    11'b00011111101: data <= 32'hbd8dc067;
    11'b00011111110: data <= 32'hbbbabc37;
    11'b00011111111: data <= 32'hbab731a4;
    11'b00100000000: data <= 32'hb70bb05f;
    11'b00100000001: data <= 32'h3862bb3e;
    11'b00100000010: data <= 32'h3b8fb2f3;
    11'b00100000011: data <= 32'hb3f53e50;
    11'b00100000100: data <= 32'hbf4b40c6;
    11'b00100000101: data <= 32'hbed43dde;
    11'b00100000110: data <= 32'ha39f32e3;
    11'b00100000111: data <= 32'h3c17b201;
    11'b00100001000: data <= 32'h3661b2d4;
    11'b00100001001: data <= 32'hb29db786;
    11'b00100001010: data <= 32'h3aa8b592;
    11'b00100001011: data <= 32'h40d0393a;
    11'b00100001100: data <= 32'h40853dab;
    11'b00100001101: data <= 32'h358d38c9;
    11'b00100001110: data <= 32'hbca9bc49;
    11'b00100001111: data <= 32'hbc1fbe57;
    11'b00100010000: data <= 32'hb42db96e;
    11'b00100010001: data <= 32'ha9c4b41b;
    11'b00100010010: data <= 32'ha8dcbd45;
    11'b00100010011: data <= 32'h3603c05b;
    11'b00100010100: data <= 32'h3837bbc3;
    11'b00100010101: data <= 32'hb6943d77;
    11'b00100010110: data <= 32'hbe774082;
    11'b00100010111: data <= 32'hbe523c3b;
    11'b00100011000: data <= 32'hb850b4f5;
    11'b00100011001: data <= 32'hb2c5b5c0;
    11'b00100011010: data <= 32'hbbaa328e;
    11'b00100011011: data <= 32'hbbe93424;
    11'b00100011100: data <= 32'h3a423194;
    11'b00100011101: data <= 32'h41473a10;
    11'b00100011110: data <= 32'h40903dbf;
    11'b00100011111: data <= 32'h31553c4e;
    11'b00100100000: data <= 32'hbc6b2504;
    11'b00100100001: data <= 32'hb6a9b5c0;
    11'b00100100010: data <= 32'h398aa62c;
    11'b00100100011: data <= 32'h39a8b721;
    11'b00100100100: data <= 32'h32d3bfd7;
    11'b00100100101: data <= 32'h360bc159;
    11'b00100100110: data <= 32'h3a7cbc94;
    11'b00100100111: data <= 32'h36203c95;
    11'b00100101000: data <= 32'hb9743e5b;
    11'b00100101001: data <= 32'hbcad2a15;
    11'b00100101010: data <= 32'hbbe9bc87;
    11'b00100101011: data <= 32'hbcd4b8c6;
    11'b00100101100: data <= 32'hbf6c361d;
    11'b00100101101: data <= 32'hbdcb34e5;
    11'b00100101110: data <= 32'h3819b35e;
    11'b00100101111: data <= 32'h40373182;
    11'b00100110000: data <= 32'h3db63d2c;
    11'b00100110001: data <= 32'hb8673efa;
    11'b00100110010: data <= 32'hbcd93cf8;
    11'b00100110011: data <= 32'h27463a2b;
    11'b00100110100: data <= 32'h3c923890;
    11'b00100110101: data <= 32'h39c5b420;
    11'b00100110110: data <= 32'hab5fbede;
    11'b00100110111: data <= 32'h36a6c055;
    11'b00100111000: data <= 32'h3e4cb983;
    11'b00100111001: data <= 32'h3eb13c3c;
    11'b00100111010: data <= 32'h37d23b20;
    11'b00100111011: data <= 32'hb900ba24;
    11'b00100111100: data <= 32'hbc12be11;
    11'b00100111101: data <= 32'hbd66b863;
    11'b00100111110: data <= 32'hbf253514;
    11'b00100111111: data <= 32'hbd57b5e8;
    11'b00101000000: data <= 32'h3328bda3;
    11'b00101000001: data <= 32'h3d00bb01;
    11'b00101000010: data <= 32'h36503b8a;
    11'b00101000011: data <= 32'hbcb0402e;
    11'b00101000100: data <= 32'hbd0d3f3a;
    11'b00101000101: data <= 32'h2de43c86;
    11'b00101000110: data <= 32'h39fa3a28;
    11'b00101000111: data <= 32'hb18d315e;
    11'b00101001000: data <= 32'hbafbbab9;
    11'b00101001001: data <= 32'h34f0bc77;
    11'b00101001010: data <= 32'h407fa6e0;
    11'b00101001011: data <= 32'h41403c46;
    11'b00101001100: data <= 32'h3cc238b8;
    11'b00101001101: data <= 32'hb3b3ba34;
    11'b00101001110: data <= 32'hb8c6bc1c;
    11'b00101001111: data <= 32'hb8e5a4e8;
    11'b00101010000: data <= 32'hbb453323;
    11'b00101010001: data <= 32'hba94bd13;
    11'b00101010010: data <= 32'h2bffc145;
    11'b00101010011: data <= 32'h394abf25;
    11'b00101010100: data <= 32'ha80c3849;
    11'b00101010101: data <= 32'hbc6b3f69;
    11'b00101010110: data <= 32'hbc063d7b;
    11'b00101010111: data <= 32'hae923881;
    11'b00101011000: data <= 32'hb24f3827;
    11'b00101011001: data <= 32'hbde9388d;
    11'b00101011010: data <= 32'hbf572754;
    11'b00101011011: data <= 32'h245db59a;
    11'b00101011100: data <= 32'h40ad3357;
    11'b00101011101: data <= 32'h413f3be7;
    11'b00101011110: data <= 32'h3c083a0d;
    11'b00101011111: data <= 32'hb2ea254f;
    11'b00101100000: data <= 32'h20413069;
    11'b00101100001: data <= 32'h37483aa7;
    11'b00101100010: data <= 32'h2c043507;
    11'b00101100011: data <= 32'hb694bef4;
    11'b00101100100: data <= 32'h9b12c239;
    11'b00101100101: data <= 32'h3944c001;
    11'b00101100110: data <= 32'h377534d3;
    11'b00101100111: data <= 32'hb3c83cb7;
    11'b00101101000: data <= 32'hb6513444;
    11'b00101101001: data <= 32'hb3cab735;
    11'b00101101010: data <= 32'hbbf02fd9;
    11'b00101101011: data <= 32'hc0b93a47;
    11'b00101101100: data <= 32'hc0c33554;
    11'b00101101101: data <= 32'hb51fb75f;
    11'b00101101110: data <= 32'h3f18b43a;
    11'b00101101111: data <= 32'h3ec53938;
    11'b00101110000: data <= 32'h30353c64;
    11'b00101110001: data <= 32'hb78a3c15;
    11'b00101110010: data <= 32'h37883d0a;
    11'b00101110011: data <= 32'h3c883e3a;
    11'b00101110100: data <= 32'h35d838ff;
    11'b00101110101: data <= 32'hb88dbdbd;
    11'b00101110110: data <= 32'hb05ac115;
    11'b00101110111: data <= 32'h3c5fbdb2;
    11'b00101111000: data <= 32'h3e0f3574;
    11'b00101111001: data <= 32'h3b5b3795;
    11'b00101111010: data <= 32'h3515ba03;
    11'b00101111011: data <= 32'hae29bc77;
    11'b00101111100: data <= 32'hbc3028cb;
    11'b00101111101: data <= 32'hc0803ae7;
    11'b00101111110: data <= 32'hc062a541;
    11'b00101111111: data <= 32'hb81cbd89;
    11'b00110000000: data <= 32'h3b4ebd30;
    11'b00110000001: data <= 32'h37a72ee6;
    11'b00110000010: data <= 32'hba163ce2;
    11'b00110000011: data <= 32'hb9623de1;
    11'b00110000100: data <= 32'h392f3e65;
    11'b00110000101: data <= 32'h3c2f3eed;
    11'b00110000110: data <= 32'hb4323bfa;
    11'b00110000111: data <= 32'hbd6db865;
    11'b00110001000: data <= 32'hb730bd55;
    11'b00110001001: data <= 32'h3e07b80d;
    11'b00110001010: data <= 32'h40a7381b;
    11'b00110001011: data <= 32'h3e772d86;
    11'b00110001100: data <= 32'h39ddbc36;
    11'b00110001101: data <= 32'h352bbb3c;
    11'b00110001110: data <= 32'hb4a1382a;
    11'b00110001111: data <= 32'hbcf43bcc;
    11'b00110010000: data <= 32'hbdcab918;
    11'b00110010001: data <= 32'hb813c0e4;
    11'b00110010010: data <= 32'h342dc06f;
    11'b00110010011: data <= 32'hb342b61c;
    11'b00110010100: data <= 32'hbbdb3b71;
    11'b00110010101: data <= 32'hb7c33bf9;
    11'b00110010110: data <= 32'h39333b60;
    11'b00110010111: data <= 32'h36673d24;
    11'b00110011000: data <= 32'hbd8b3cf8;
    11'b00110011001: data <= 32'hc0ad35d3;
    11'b00110011010: data <= 32'hbaf3b4dd;
    11'b00110011011: data <= 32'h3df82a13;
    11'b00110011100: data <= 32'h4089383c;
    11'b00110011101: data <= 32'h3d6a2cad;
    11'b00110011110: data <= 32'h38ddb881;
    11'b00110011111: data <= 32'h3a5d2c08;
    11'b00110100000: data <= 32'h3a7e3d93;
    11'b00110100001: data <= 32'ha5ce3ceb;
    11'b00110100010: data <= 32'hb9dfbba3;
    11'b00110100011: data <= 32'hb734c1b3;
    11'b00110100100: data <= 32'h2e71c0c4;
    11'b00110100101: data <= 32'ha91bb828;
    11'b00110100110: data <= 32'hb56d35aa;
    11'b00110100111: data <= 32'h308fb072;
    11'b00110101000: data <= 32'h3996b506;
    11'b00110101001: data <= 32'hb29338bb;
    11'b00110101010: data <= 32'hc05d3d3e;
    11'b00110101011: data <= 32'hc1b93a67;
    11'b00110101100: data <= 32'hbca8ae9a;
    11'b00110101101: data <= 32'h3bdeb27f;
    11'b00110101110: data <= 32'h3d36323d;
    11'b00110101111: data <= 32'h347432c5;
    11'b00110110000: data <= 32'h2c9832dd;
    11'b00110110001: data <= 32'h3c663c57;
    11'b00110110010: data <= 32'h3e664040;
    11'b00110110011: data <= 32'h38b43e38;
    11'b00110110100: data <= 32'hb8feb94e;
    11'b00110110101: data <= 32'hb873c07b;
    11'b00110110110: data <= 32'h354abe88;
    11'b00110110111: data <= 32'h3a13b336;
    11'b00110111000: data <= 32'h39a5b236;
    11'b00110111001: data <= 32'h3b13bd00;
    11'b00110111010: data <= 32'h3b50bd21;
    11'b00110111011: data <= 32'hb34a32f9;
    11'b00110111100: data <= 32'hc00f3d54;
    11'b00110111101: data <= 32'hc1113926;
    11'b00110111110: data <= 32'hbc90ba0d;
    11'b00110111111: data <= 32'h3447bc63;
    11'b00111000000: data <= 32'h1dc4b643;
    11'b00111000001: data <= 32'hbb4732ff;
    11'b00111000010: data <= 32'hb6f238b2;
    11'b00111000011: data <= 32'h3cc43d84;
    11'b00111000100: data <= 32'h3ec84067;
    11'b00111000101: data <= 32'h33de3f07;
    11'b00111000110: data <= 32'hbcfd2e48;
    11'b00111000111: data <= 32'hbb49bba9;
    11'b00111001000: data <= 32'h38c1b6e2;
    11'b00111001001: data <= 32'h3dd2342a;
    11'b00111001010: data <= 32'h3d6bb78d;
    11'b00111001011: data <= 32'h3cf9bee2;
    11'b00111001100: data <= 32'h3ce0bd7a;
    11'b00111001101: data <= 32'h36f53811;
    11'b00111001110: data <= 32'hbb9b3de6;
    11'b00111001111: data <= 32'hbe183264;
    11'b00111010000: data <= 32'hba97beab;
    11'b00111010001: data <= 32'hb41fbfd8;
    11'b00111010010: data <= 32'hbadabae8;
    11'b00111010011: data <= 32'hbdc5a3db;
    11'b00111010100: data <= 32'hb7833199;
    11'b00111010101: data <= 32'h3cd23926;
    11'b00111010110: data <= 32'h3cef3e12;
    11'b00111010111: data <= 32'hb9923ed0;
    11'b00111011000: data <= 32'hc0533aff;
    11'b00111011001: data <= 32'hbd5f32f4;
    11'b00111011010: data <= 32'h38a6372e;
    11'b00111011011: data <= 32'h3dae3841;
    11'b00111011100: data <= 32'h3c2ab790;
    11'b00111011101: data <= 32'h3b5abdb0;
    11'b00111011110: data <= 32'h3dafb8e2;
    11'b00111011111: data <= 32'h3d983d33;
    11'b00111100000: data <= 32'h36673f0d;
    11'b00111100001: data <= 32'hb7a7ac98;
    11'b00111100010: data <= 32'hb7aac01e;
    11'b00111100011: data <= 32'hb60dc02b;
    11'b00111100100: data <= 32'hbae7bac1;
    11'b00111100101: data <= 32'hbc25b5d0;
    11'b00111100110: data <= 32'h2b02baac;
    11'b00111100111: data <= 32'h3d32b9ba;
    11'b00111101000: data <= 32'h39b737ea;
    11'b00111101001: data <= 32'hbdcd3ddc;
    11'b00111101010: data <= 32'hc14d3cfa;
    11'b00111101011: data <= 32'hbe1c38e3;
    11'b00111101100: data <= 32'h3405376f;
    11'b00111101101: data <= 32'h3880354c;
    11'b00111101110: data <= 32'hb0aeb61a;
    11'b00111101111: data <= 32'h2c35ba1a;
    11'b00111110000: data <= 32'h3da3356a;
    11'b00111110001: data <= 32'h40324001;
    11'b00111110010: data <= 32'h3ccd400b;
    11'b00111110011: data <= 32'hacac2dcd;
    11'b00111110100: data <= 32'hb69ebe26;
    11'b00111110101: data <= 32'hb1f1bcf0;
    11'b00111110110: data <= 32'hb2a8b418;
    11'b00111110111: data <= 32'hae25b8cb;
    11'b00111111000: data <= 32'h3a28bf61;
    11'b00111111001: data <= 32'h3df5bf7b;
    11'b00111111010: data <= 32'h38e7b260;
    11'b00111111011: data <= 32'hbd723d19;
    11'b00111111100: data <= 32'hc07b3c6c;
    11'b00111111101: data <= 32'hbcf62fc5;
    11'b00111111110: data <= 32'hb16cb4a7;
    11'b00111111111: data <= 32'hb90ab30e;
    11'b01000000000: data <= 32'hbe11b61e;
    11'b01000000001: data <= 32'hba3bb5be;
    11'b01000000010: data <= 32'h3d043967;
    11'b01000000011: data <= 32'h40624009;
    11'b01000000100: data <= 32'h3c254000;
    11'b01000000101: data <= 32'hb82b38ab;
    11'b01000000110: data <= 32'hb9b6b5b1;
    11'b01000000111: data <= 32'h2a3130a9;
    11'b01000001000: data <= 32'h379738a4;
    11'b01000001001: data <= 32'h3895b8d1;
    11'b01000001010: data <= 32'h3c5bc095;
    11'b01000001011: data <= 32'h3e7ac04b;
    11'b01000001100: data <= 32'h3c2bafc0;
    11'b01000001101: data <= 32'hb6173d55;
    11'b01000001110: data <= 32'hbc40399b;
    11'b01000001111: data <= 32'hb892b9e9;
    11'b01000010000: data <= 32'hb666bc99;
    11'b01000010001: data <= 32'hbdcfb95d;
    11'b01000010010: data <= 32'hc080b7df;
    11'b01000010011: data <= 32'hbc43b8a3;
    11'b01000010100: data <= 32'h3c99281d;
    11'b01000010101: data <= 32'h3f113cbd;
    11'b01000010110: data <= 32'h319c3e6e;
    11'b01000010111: data <= 32'hbd9c3c39;
    11'b01000011000: data <= 32'hbc883a24;
    11'b01000011001: data <= 32'h2f443cf3;
    11'b01000011010: data <= 32'h38b13c90;
    11'b01000011011: data <= 32'h357eb729;
    11'b01000011100: data <= 32'h391fc00c;
    11'b01000011101: data <= 32'h3e07bdfd;
    11'b01000011110: data <= 32'h3ed238d8;
    11'b01000011111: data <= 32'h3b473e71;
    11'b01000100000: data <= 32'h32883634;
    11'b01000100001: data <= 32'h2e35bcf1;
    11'b01000100010: data <= 32'hb53bbd61;
    11'b01000100011: data <= 32'hbdedb871;
    11'b01000100100: data <= 32'hbfeeb87f;
    11'b01000100101: data <= 32'hb922bd36;
    11'b01000100110: data <= 32'h3ce4bd0b;
    11'b01000100111: data <= 32'h3cefabce;
    11'b01000101000: data <= 32'hb9283c12;
    11'b01000101001: data <= 32'hbfd03cca;
    11'b01000101010: data <= 32'hbd003cb2;
    11'b01000101011: data <= 32'h24983dad;
    11'b01000101100: data <= 32'ha16e3c55;
    11'b01000101101: data <= 32'hba33b510;
    11'b01000101110: data <= 32'hb6d6bd7b;
    11'b01000101111: data <= 32'h3c87b823;
    11'b01000110000: data <= 32'h404c3d6e;
    11'b01000110001: data <= 32'h3ed93f4e;
    11'b01000110010: data <= 32'h3a6c35c6;
    11'b01000110011: data <= 32'h35adbb8d;
    11'b01000110100: data <= 32'hac35b889;
    11'b01000110101: data <= 32'hbac4336b;
    11'b01000110110: data <= 32'hbc2eb700;
    11'b01000110111: data <= 32'h2eb4c015;
    11'b01000111000: data <= 32'h3d91c0d1;
    11'b01000111001: data <= 32'h3be3bbc7;
    11'b01000111010: data <= 32'hba0f38b1;
    11'b01000111011: data <= 32'hbe783ba1;
    11'b01000111100: data <= 32'hba4c39ae;
    11'b01000111101: data <= 32'hab3f39a4;
    11'b01000111110: data <= 32'hbb673837;
    11'b01000111111: data <= 32'hc043b4f4;
    11'b01001000000: data <= 32'hbe08bae4;
    11'b01001000001: data <= 32'h39879fee;
    11'b01001000010: data <= 32'h40323dce;
    11'b01001000011: data <= 32'h3e4c3ea4;
    11'b01001000100: data <= 32'h36f23842;
    11'b01001000101: data <= 32'h2d82a8b6;
    11'b01001000110: data <= 32'h31973a5c;
    11'b01001000111: data <= 32'hadee3d43;
    11'b01001001000: data <= 32'hb387afb0;
    11'b01001001001: data <= 32'h3811c09f;
    11'b01001001010: data <= 32'h3da4c16c;
    11'b01001001011: data <= 32'h3c81bc0c;
    11'b01001001100: data <= 32'ha956388d;
    11'b01001001101: data <= 32'hb76a383e;
    11'b01001001110: data <= 32'h3043b233;
    11'b01001001111: data <= 32'h2b58b431;
    11'b01001010000: data <= 32'hbe2f9f14;
    11'b01001010001: data <= 32'hc1cab57c;
    11'b01001010010: data <= 32'hbfcdbaa7;
    11'b01001010011: data <= 32'h3761b65f;
    11'b01001010100: data <= 32'h3e89393c;
    11'b01001010101: data <= 32'h39853c16;
    11'b01001010110: data <= 32'hb82a392e;
    11'b01001010111: data <= 32'hb6883aeb;
    11'b01001011000: data <= 32'h34983fad;
    11'b01001011001: data <= 32'h33534024;
    11'b01001011010: data <= 32'hb34c32bd;
    11'b01001011011: data <= 32'h2f10bfe9;
    11'b01001011100: data <= 32'h3c4cc01b;
    11'b01001011101: data <= 32'h3dbab3f7;
    11'b01001011110: data <= 32'h3c0d3b36;
    11'b01001011111: data <= 32'h3ab2320c;
    11'b01001100000: data <= 32'h3c1fbae6;
    11'b01001100001: data <= 32'h35b2b967;
    11'b01001100010: data <= 32'hbdec2942;
    11'b01001100011: data <= 32'hc144b309;
    11'b01001100100: data <= 32'hbe20bcd8;
    11'b01001100101: data <= 32'h387fbdc9;
    11'b01001100110: data <= 32'h3c52b8f9;
    11'b01001100111: data <= 32'hb44e31af;
    11'b01001101000: data <= 32'hbd143823;
    11'b01001101001: data <= 32'hb8d83c99;
    11'b01001101010: data <= 32'h359a403f;
    11'b01001101011: data <= 32'ha9fe4020;
    11'b01001101100: data <= 32'hbc6535a0;
    11'b01001101101: data <= 32'hbbd4bd37;
    11'b01001101110: data <= 32'h36e4bbb1;
    11'b01001101111: data <= 32'h3e45396e;
    11'b01001110000: data <= 32'h3eac3cd5;
    11'b01001110001: data <= 32'h3de628d1;
    11'b01001110010: data <= 32'h3d8fbae9;
    11'b01001110011: data <= 32'h3963b095;
    11'b01001110100: data <= 32'hba883aaf;
    11'b01001110101: data <= 32'hbe713188;
    11'b01001110110: data <= 32'hb913be7a;
    11'b01001110111: data <= 32'h3a9bc0da;
    11'b01001111000: data <= 32'h39e9be57;
    11'b01001111001: data <= 32'hb92eb680;
    11'b01001111010: data <= 32'hbcb4314c;
    11'b01001111011: data <= 32'hb0e83925;
    11'b01001111100: data <= 32'h38403d67;
    11'b01001111101: data <= 32'hb8fb3d90;
    11'b01001111110: data <= 32'hc08b344f;
    11'b01001111111: data <= 32'hc03db9cd;
    11'b01010000000: data <= 32'hb2a2b2d8;
    11'b01010000001: data <= 32'h3d6d3c0f;
    11'b01010000010: data <= 32'h3de03c4c;
    11'b01010000011: data <= 32'h3c4ca6a5;
    11'b01010000100: data <= 32'h3c31b4b9;
    11'b01010000101: data <= 32'h3abe3c18;
    11'b01010000110: data <= 32'ha2703ff1;
    11'b01010000111: data <= 32'hb8b639c8;
    11'b01010001000: data <= 32'h1f96beb9;
    11'b01010001001: data <= 32'h3b34c14b;
    11'b01010001010: data <= 32'h395fbe7b;
    11'b01010001011: data <= 32'hb437b66f;
    11'b01010001100: data <= 32'hb349b2fe;
    11'b01010001101: data <= 32'h3aa7b4d5;
    11'b01010001110: data <= 32'h3b39326c;
    11'b01010001111: data <= 32'hbbf73906;
    11'b01010010000: data <= 32'hc1df3107;
    11'b01010010001: data <= 32'hc12bb828;
    11'b01010010010: data <= 32'hb786b489;
    11'b01010010011: data <= 32'h3b1e36f5;
    11'b01010010100: data <= 32'h38593619;
    11'b01010010101: data <= 32'ha850b1d4;
    11'b01010010110: data <= 32'h35823547;
    11'b01010010111: data <= 32'h3ae54012;
    11'b01010011000: data <= 32'h37424193;
    11'b01010011001: data <= 32'hb4693c91;
    11'b01010011010: data <= 32'hb11cbd32;
    11'b01010011011: data <= 32'h383dbfc5;
    11'b01010011100: data <= 32'h39a2b9de;
    11'b01010011101: data <= 32'h37e22f25;
    11'b01010011110: data <= 32'h3b96b76b;
    11'b01010011111: data <= 32'h3f34bc5a;
    11'b01010100000: data <= 32'h3d5fb801;
    11'b01010100001: data <= 32'hbab336ee;
    11'b01010100010: data <= 32'hc13e349a;
    11'b01010100011: data <= 32'hc026b918;
    11'b01010100100: data <= 32'hb337bc14;
    11'b01010100101: data <= 32'h36c5b99f;
    11'b01010100110: data <= 32'hb81db86b;
    11'b01010100111: data <= 32'hbc35b802;
    11'b01010101000: data <= 32'haea637a4;
    11'b01010101001: data <= 32'h3b39405d;
    11'b01010101010: data <= 32'h36b54174;
    11'b01010101011: data <= 32'hba9f3cbd;
    11'b01010101100: data <= 32'hbc5fb989;
    11'b01010101101: data <= 32'hb2b0ba1e;
    11'b01010101110: data <= 32'h38e8371a;
    11'b01010101111: data <= 32'h3bc3395f;
    11'b01010110000: data <= 32'h3e19b889;
    11'b01010110001: data <= 32'h404bbd3a;
    11'b01010110010: data <= 32'h3e77b49f;
    11'b01010110011: data <= 32'hb2c83c36;
    11'b01010110100: data <= 32'hbe163a26;
    11'b01010110101: data <= 32'hbb99ba5a;
    11'b01010110110: data <= 32'h3493bf25;
    11'b01010110111: data <= 32'h30c1be65;
    11'b01010111000: data <= 32'hbc59bca6;
    11'b01010111001: data <= 32'hbd1cbaf3;
    11'b01010111010: data <= 32'h30e2a676;
    11'b01010111011: data <= 32'h3c9f3d5d;
    11'b01010111100: data <= 32'h2eb53f6c;
    11'b01010111101: data <= 32'hbf0a3af5;
    11'b01010111110: data <= 32'hc051b229;
    11'b01010111111: data <= 32'hbb423109;
    11'b01011000000: data <= 32'h353a3c64;
    11'b01011000001: data <= 32'h39e23a09;
    11'b01011000010: data <= 32'h3c41b971;
    11'b01011000011: data <= 32'h3e94bc00;
    11'b01011000100: data <= 32'h3e5238f0;
    11'b01011000101: data <= 32'h3814403b;
    11'b01011000110: data <= 32'hb57f3d9e;
    11'b01011000111: data <= 32'h1ef3b9d3;
    11'b01011001000: data <= 32'h38ccbfba;
    11'b01011001001: data <= 32'h2b6cbe52;
    11'b01011001010: data <= 32'hbbadbc2b;
    11'b01011001011: data <= 32'hb8dbbc5b;
    11'b01011001100: data <= 32'h3c26bb2b;
    11'b01011001101: data <= 32'h3e842a92;
    11'b01011001110: data <= 32'hae4b3a4b;
    11'b01011001111: data <= 32'hc0a03801;
    11'b01011010000: data <= 32'hc1262071;
    11'b01011010001: data <= 32'hbc68355c;
    11'b01011010010: data <= 32'ha7003a80;
    11'b01011010011: data <= 32'hb04a31d0;
    11'b01011010100: data <= 32'hb16abb8b;
    11'b01011010101: data <= 32'h3936b89f;
    11'b01011010110: data <= 32'h3d563df3;
    11'b01011010111: data <= 32'h3b9241c0;
    11'b01011011000: data <= 32'h328f3f34;
    11'b01011011001: data <= 32'h30d7b673;
    11'b01011011010: data <= 32'h3605bd08;
    11'b01011011011: data <= 32'ha113b8a9;
    11'b01011011100: data <= 32'hb6e0b43f;
    11'b01011011101: data <= 32'h366abc4c;
    11'b01011011110: data <= 32'h3fdfbe89;
    11'b01011011111: data <= 32'h402ebaf9;
    11'b01011100000: data <= 32'h2b7b3440;
    11'b01011100001: data <= 32'hc000373c;
    11'b01011100010: data <= 32'hbfe0a638;
    11'b01011100011: data <= 32'hb907b11a;
    11'b01011100100: data <= 32'hb411b02a;
    11'b01011100101: data <= 32'hbc8bb9b2;
    11'b01011100110: data <= 32'hbd95bd49;
    11'b01011100111: data <= 32'hb03ab7b1;
    11'b01011101000: data <= 32'h3ca93e73;
    11'b01011101001: data <= 32'h3bc74179;
    11'b01011101010: data <= 32'hae303ea1;
    11'b01011101011: data <= 32'hb8789d89;
    11'b01011101100: data <= 32'hb4ffb04b;
    11'b01011101101: data <= 32'hb20e3a55;
    11'b01011101110: data <= 32'haa73390e;
    11'b01011101111: data <= 32'h3b6fbb8b;
    11'b01011110000: data <= 32'h4083bf8e;
    11'b01011110001: data <= 32'h4073bb4d;
    11'b01011110010: data <= 32'h381c3913;
    11'b01011110011: data <= 32'hbb973ae6;
    11'b01011110100: data <= 32'hb949acf5;
    11'b01011110101: data <= 32'h32edba4a;
    11'b01011110110: data <= 32'hb46ebba0;
    11'b01011110111: data <= 32'hbee5bd24;
    11'b01011111000: data <= 32'hbf7fbe6c;
    11'b01011111001: data <= 32'hb0eabadf;
    11'b01011111010: data <= 32'h3d473a75;
    11'b01011111011: data <= 32'h3a1c3ecc;
    11'b01011111100: data <= 32'hbadd3c17;
    11'b01011111101: data <= 32'hbe1a338a;
    11'b01011111110: data <= 32'hbbe93a4b;
    11'b01011111111: data <= 32'hb71c3ecb;
    11'b01100000000: data <= 32'hb2c43c14;
    11'b01100000001: data <= 32'h37e3bb67;
    11'b01100000010: data <= 32'h3e73beb8;
    11'b01100000011: data <= 32'h3f98b272;
    11'b01100000100: data <= 32'h3bda3e48;
    11'b01100000101: data <= 32'h32f23dee;
    11'b01100000110: data <= 32'h386618a2;
    11'b01100000111: data <= 32'h3ae0bba4;
    11'b01100001000: data <= 32'hb286bb8d;
    11'b01100001001: data <= 32'hbebabc34;
    11'b01100001010: data <= 32'hbdacbe4b;
    11'b01100001011: data <= 32'h389bbdf9;
    11'b01100001100: data <= 32'h3f18b76b;
    11'b01100001101: data <= 32'h38df3614;
    11'b01100001110: data <= 32'hbd8e34e3;
    11'b01100001111: data <= 32'hbfbe33ba;
    11'b01100010000: data <= 32'hbc653c26;
    11'b01100010001: data <= 32'hb8c33e96;
    11'b01100010010: data <= 32'hbafc3913;
    11'b01100010011: data <= 32'hb9bebca1;
    11'b01100010100: data <= 32'h3610bd52;
    11'b01100010101: data <= 32'h3d2d38dc;
    11'b01100010110: data <= 32'h3cc8409e;
    11'b01100010111: data <= 32'h3a973f4a;
    11'b01100011000: data <= 32'h3b9131a8;
    11'b01100011001: data <= 32'h3ae2b73a;
    11'b01100011010: data <= 32'hb30a281f;
    11'b01100011011: data <= 32'hbcf5aac4;
    11'b01100011100: data <= 32'hb80dbcd3;
    11'b01100011101: data <= 32'h3de0bff8;
    11'b01100011110: data <= 32'h4068bdb9;
    11'b01100011111: data <= 32'h3955b689;
    11'b01100100000: data <= 32'hbcd49fee;
    11'b01100100001: data <= 32'hbd643012;
    11'b01100100010: data <= 32'hb6d93919;
    11'b01100100011: data <= 32'hb7d03aa9;
    11'b01100100100: data <= 32'hbe88b273;
    11'b01100100101: data <= 32'hbfe9be18;
    11'b01100100110: data <= 32'hb976bcb9;
    11'b01100100111: data <= 32'h3a943a98;
    11'b01100101000: data <= 32'h3c6c405f;
    11'b01100101001: data <= 32'h38f03e0b;
    11'b01100101010: data <= 32'h365a3455;
    11'b01100101011: data <= 32'h341f3701;
    11'b01100101100: data <= 32'hb6563dbb;
    11'b01100101101: data <= 32'hbacd3c83;
    11'b01100101110: data <= 32'h2cf5b9ef;
    11'b01100101111: data <= 32'h3f19c031;
    11'b01100110000: data <= 32'h4069be3f;
    11'b01100110001: data <= 32'h3adbb375;
    11'b01100110010: data <= 32'hb5f7347b;
    11'b01100110011: data <= 32'ha45f2c51;
    11'b01100110100: data <= 32'h39992871;
    11'b01100110101: data <= 32'hb115a0b5;
    11'b01100110110: data <= 32'hc016ba54;
    11'b01100110111: data <= 32'hc115bed9;
    11'b01100111000: data <= 32'hbb6bbd5c;
    11'b01100111001: data <= 32'h3a7f32eb;
    11'b01100111010: data <= 32'h3b003c88;
    11'b01100111011: data <= 32'hae1838d3;
    11'b01100111100: data <= 32'hb86a30db;
    11'b01100111101: data <= 32'hb6da3ca6;
    11'b01100111110: data <= 32'hb8bd40d8;
    11'b01100111111: data <= 32'hbaba3f12;
    11'b01101000000: data <= 32'hb1f5b81f;
    11'b01101000001: data <= 32'h3c7ebf5e;
    11'b01101000010: data <= 32'h3e7fbb53;
    11'b01101000011: data <= 32'h3bc03932;
    11'b01101000100: data <= 32'h38b03b28;
    11'b01101000101: data <= 32'h3d182f73;
    11'b01101000110: data <= 32'h3e7bb419;
    11'b01101000111: data <= 32'h3150b0aa;
    11'b01101001000: data <= 32'hbfb6b87f;
    11'b01101001001: data <= 32'hc052bdd4;
    11'b01101001010: data <= 32'hb49ebe8a;
    11'b01101001011: data <= 32'h3cf2babf;
    11'b01101001100: data <= 32'h39a6b43a;
    11'b01101001101: data <= 32'hb9a3b6a0;
    11'b01101001110: data <= 32'hbc50b049;
    11'b01101001111: data <= 32'hb8723d40;
    11'b01101010000: data <= 32'hb87940e9;
    11'b01101010001: data <= 32'hbcc63e0b;
    11'b01101010010: data <= 32'hbcc1b97f;
    11'b01101010011: data <= 32'hb1cdbdee;
    11'b01101010100: data <= 32'h39abac0f;
    11'b01101010101: data <= 32'h3ade3de7;
    11'b01101010110: data <= 32'h3c453d0b;
    11'b01101010111: data <= 32'h3f1130b8;
    11'b01101011000: data <= 32'h3f2ba619;
    11'b01101011001: data <= 32'h33f2390c;
    11'b01101011010: data <= 32'hbde337ee;
    11'b01101011011: data <= 32'hbcf0ba3d;
    11'b01101011100: data <= 32'h3950bf28;
    11'b01101011101: data <= 32'h3ec9bea8;
    11'b01101011110: data <= 32'h3943bca3;
    11'b01101011111: data <= 32'hba08bb8a;
    11'b01101100000: data <= 32'hb96bb646;
    11'b01101100001: data <= 32'h311c3b1c;
    11'b01101100010: data <= 32'hb1043e9e;
    11'b01101100011: data <= 32'hbe67392f;
    11'b01101100100: data <= 32'hc092bc53;
    11'b01101100101: data <= 32'hbd6cbd0a;
    11'b01101100110: data <= 32'ha4ef3585;
    11'b01101100111: data <= 32'h389b3e1b;
    11'b01101101000: data <= 32'h3a8e3b62;
    11'b01101101001: data <= 32'h3d05a75f;
    11'b01101101010: data <= 32'h3ccd382a;
    11'b01101101011: data <= 32'h2b2b3f71;
    11'b01101101100: data <= 32'hbc233f2c;
    11'b01101101101: data <= 32'hb7efa6ac;
    11'b01101101110: data <= 32'h3c85be9d;
    11'b01101101111: data <= 32'h3ec6beee;
    11'b01101110000: data <= 32'h38e1bc2e;
    11'b01101110001: data <= 32'hb3f0b9b1;
    11'b01101110010: data <= 32'h37a8b75a;
    11'b01101110011: data <= 32'h3d9c3415;
    11'b01101110100: data <= 32'h37be3989;
    11'b01101110101: data <= 32'hbeefad9f;
    11'b01101110110: data <= 32'hc189bd23;
    11'b01101110111: data <= 32'hbebdbcdf;
    11'b01101111000: data <= 32'hb0622992;
    11'b01101111001: data <= 32'h34d23930;
    11'b01101111010: data <= 32'h2d52ae00;
    11'b01101111011: data <= 32'h330fb784;
    11'b01101111100: data <= 32'h36373b88;
    11'b01101111101: data <= 32'hb1894180;
    11'b01101111110: data <= 32'hbae94113;
    11'b01101111111: data <= 32'hb7aa35bd;
    11'b01110000000: data <= 32'h3942bd3f;
    11'b01110000001: data <= 32'h3c12bc3d;
    11'b01110000010: data <= 32'h366aaf0a;
    11'b01110000011: data <= 32'h363f135b;
    11'b01110000100: data <= 32'h3ea4b5eb;
    11'b01110000101: data <= 32'h40e5b123;
    11'b01110000110: data <= 32'h3c1034dd;
    11'b01110000111: data <= 32'hbdf2a949;
    11'b01110001000: data <= 32'hc0b4bbad;
    11'b01110001001: data <= 32'hbc19bcd2;
    11'b01110001010: data <= 32'h3599b981;
    11'b01110001011: data <= 32'h3168b90b;
    11'b01110001100: data <= 32'hb8f8bd03;
    11'b01110001101: data <= 32'hb838bc07;
    11'b01110001110: data <= 32'h2d023b54;
    11'b01110001111: data <= 32'hae4c417c;
    11'b01110010000: data <= 32'hbb794095;
    11'b01110010001: data <= 32'hbc9e3160;
    11'b01110010010: data <= 32'hb827bbc9;
    11'b01110010011: data <= 32'haa34b044;
    11'b01110010100: data <= 32'h19113b43;
    11'b01110010101: data <= 32'h3943385f;
    11'b01110010110: data <= 32'h4036b5a1;
    11'b01110010111: data <= 32'h4155b1af;
    11'b01110011000: data <= 32'h3c843a18;
    11'b01110011001: data <= 32'hbc1b3b04;
    11'b01110011010: data <= 32'hbd75b049;
    11'b01110011011: data <= 32'h2dccbc2f;
    11'b01110011100: data <= 32'h3bd5bd0b;
    11'b01110011101: data <= 32'h302ebde3;
    11'b01110011110: data <= 32'hbb16bf75;
    11'b01110011111: data <= 32'hb6e3bd68;
    11'b01110100000: data <= 32'h39223749;
    11'b01110100001: data <= 32'h37043f8e;
    11'b01110100010: data <= 32'hbc133d2f;
    11'b01110100011: data <= 32'hbfe9b612;
    11'b01110100100: data <= 32'hbe89ba35;
    11'b01110100101: data <= 32'hbb283758;
    11'b01110100110: data <= 32'hb6ca3cfd;
    11'b01110100111: data <= 32'h355c35f5;
    11'b01110101000: data <= 32'h3e32b91f;
    11'b01110101001: data <= 32'h3feb2a32;
    11'b01110101010: data <= 32'h3a793ecf;
    11'b01110101011: data <= 32'hb8f94036;
    11'b01110101100: data <= 32'hb77f3a1e;
    11'b01110101101: data <= 32'h3aa3b9b5;
    11'b01110101110: data <= 32'h3c9cbcdc;
    11'b01110101111: data <= 32'h998abd46;
    11'b01110110000: data <= 32'hb979be52;
    11'b01110110001: data <= 32'h36dabd51;
    11'b01110110010: data <= 32'h3f3ab0bc;
    11'b01110110011: data <= 32'h3cf73a59;
    11'b01110110100: data <= 32'hbb4634de;
    11'b01110110101: data <= 32'hc09dba2a;
    11'b01110110110: data <= 32'hbfb6b96b;
    11'b01110110111: data <= 32'hbc053716;
    11'b01110111000: data <= 32'hb943395d;
    11'b01110111001: data <= 32'hb62bb86f;
    11'b01110111010: data <= 32'h366dbd00;
    11'b01110111011: data <= 32'h3b75323b;
    11'b01110111100: data <= 32'h362d40d1;
    11'b01110111101: data <= 32'hb6c141a3;
    11'b01110111110: data <= 32'hb2053cc1;
    11'b01110111111: data <= 32'h394bb5b4;
    11'b01111000000: data <= 32'h38abb846;
    11'b01111000001: data <= 32'hb60bb49f;
    11'b01111000010: data <= 32'hb575b94d;
    11'b01111000011: data <= 32'h3d9abc33;
    11'b01111000100: data <= 32'h41a6b88b;
    11'b01111000101: data <= 32'h3f6c314c;
    11'b01111000110: data <= 32'hb8b829a0;
    11'b01111000111: data <= 32'hbf6bb899;
    11'b01111001000: data <= 32'hbcc0b81a;
    11'b01111001001: data <= 32'hb5992476;
    11'b01111001010: data <= 32'hb8f4b611;
    11'b01111001011: data <= 32'hbc51bec1;
    11'b01111001100: data <= 32'hb87fbfa3;
    11'b01111001101: data <= 32'h350e2987;
    11'b01111001110: data <= 32'h34e740aa;
    11'b01111001111: data <= 32'hb5d44104;
    11'b01111010000: data <= 32'hb8713afa;
    11'b01111010001: data <= 32'hb443b10d;
    11'b01111010010: data <= 32'hb746360f;
    11'b01111010011: data <= 32'hbb6e3b62;
    11'b01111010100: data <= 32'hb3f631d5;
    11'b01111010101: data <= 32'h3f01bad7;
    11'b01111010110: data <= 32'h41feb979;
    11'b01111010111: data <= 32'h3f913525;
    11'b01111011000: data <= 32'hb35a3991;
    11'b01111011001: data <= 32'hbaff32c0;
    11'b01111011010: data <= 32'h2e83b1c9;
    11'b01111011011: data <= 32'h3888b56b;
    11'b01111011100: data <= 32'hb775bc67;
    11'b01111011101: data <= 32'hbda8c08c;
    11'b01111011110: data <= 32'hba0bc075;
    11'b01111011111: data <= 32'h38c6b5d4;
    11'b01111100000: data <= 32'h3a433de6;
    11'b01111100001: data <= 32'hb4533d6f;
    11'b01111100010: data <= 32'hbc852b44;
    11'b01111100011: data <= 32'hbcf3b107;
    11'b01111100100: data <= 32'hbd2a3c13;
    11'b01111100101: data <= 32'hbd8a3e29;
    11'b01111100110: data <= 32'hb88f34e1;
    11'b01111100111: data <= 32'h3cb5bc3a;
    11'b01111101000: data <= 32'h405ab909;
    11'b01111101001: data <= 32'h3d533bee;
    11'b01111101010: data <= 32'ha4163f08;
    11'b01111101011: data <= 32'h2ae93c72;
    11'b01111101100: data <= 32'h3c6e3369;
    11'b01111101101: data <= 32'h3c32b3af;
    11'b01111101110: data <= 32'hb7c2bb50;
    11'b01111101111: data <= 32'hbd79bf89;
    11'b01111110000: data <= 32'hb1bec002;
    11'b01111110001: data <= 32'h3e4aba59;
    11'b01111110010: data <= 32'h3e5b35b7;
    11'b01111110011: data <= 32'ha93d2f29;
    11'b01111110100: data <= 32'hbd6cb93a;
    11'b01111110101: data <= 32'hbdebb268;
    11'b01111110110: data <= 32'hbd4f3c8f;
    11'b01111110111: data <= 32'hbddf3d03;
    11'b01111111000: data <= 32'hbc95b690;
    11'b01111111001: data <= 32'h223ebea9;
    11'b01111111010: data <= 32'h3b1fb90c;
    11'b01111111011: data <= 32'h38af3e34;
    11'b01111111100: data <= 32'h246440cd;
    11'b01111111101: data <= 32'h37373df5;
    11'b01111111110: data <= 32'h3cf037eb;
    11'b01111111111: data <= 32'h39ba355c;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    