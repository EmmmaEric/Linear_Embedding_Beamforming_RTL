
module memory_rom_21(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3e3934ec;
    11'b00000000001: data <= 32'h3acb2ff5;
    11'b00000000010: data <= 32'hbb8bb3b8;
    11'b00000000011: data <= 32'hbdc9bcc5;
    11'b00000000100: data <= 32'h3410bedb;
    11'b00000000101: data <= 32'h4022bc94;
    11'b00000000110: data <= 32'h3f06b712;
    11'b00000000111: data <= 32'habc6b878;
    11'b00000001000: data <= 32'hbc92b9d6;
    11'b00000001001: data <= 32'hbb5831b7;
    11'b00000001010: data <= 32'hba1d3d6e;
    11'b00000001011: data <= 32'hbd723b63;
    11'b00000001100: data <= 32'hbe9bbc06;
    11'b00000001101: data <= 32'hbad4bfe1;
    11'b00000001110: data <= 32'h30cdb840;
    11'b00000001111: data <= 32'h35ca3e7b;
    11'b00000010000: data <= 32'h34a7402c;
    11'b00000010001: data <= 32'h3a283c1d;
    11'b00000010010: data <= 32'h3c883752;
    11'b00000010011: data <= 32'h333b3bc6;
    11'b00000010100: data <= 32'hbce43c75;
    11'b00000010101: data <= 32'hbc6c2019;
    11'b00000010110: data <= 32'h3b56bce0;
    11'b00000010111: data <= 32'h4111bd46;
    11'b00000011000: data <= 32'h3f96ba0a;
    11'b00000011001: data <= 32'h314bb863;
    11'b00000011010: data <= 32'hb5efb74f;
    11'b00000011011: data <= 32'h3532337f;
    11'b00000011100: data <= 32'h351d3ac8;
    11'b00000011101: data <= 32'hbc2a2848;
    11'b00000011110: data <= 32'hc03cbefd;
    11'b00000011111: data <= 32'hbe42c08f;
    11'b00000100000: data <= 32'hb41db98a;
    11'b00000100001: data <= 32'h34f23c70;
    11'b00000100010: data <= 32'h31903c97;
    11'b00000100011: data <= 32'h326f3237;
    11'b00000100100: data <= 32'h326c35fa;
    11'b00000100101: data <= 32'hb8ac3efc;
    11'b00000100110: data <= 32'hbe2c406a;
    11'b00000100111: data <= 32'hbc593a25;
    11'b00000101000: data <= 32'h3a4ebba6;
    11'b00000101001: data <= 32'h4010bcae;
    11'b00000101010: data <= 32'h3d94b483;
    11'b00000101011: data <= 32'h34d333fd;
    11'b00000101100: data <= 32'h38f23366;
    11'b00000101101: data <= 32'h3ebc368d;
    11'b00000101110: data <= 32'h3d3f3890;
    11'b00000101111: data <= 32'hb9b7b3ce;
    11'b00000110000: data <= 32'hc03abecb;
    11'b00000110001: data <= 32'hbd73c03a;
    11'b00000110010: data <= 32'h3425bbd3;
    11'b00000110011: data <= 32'h3a0e2c79;
    11'b00000110100: data <= 32'h2fbab471;
    11'b00000110101: data <= 32'hb5adbae6;
    11'b00000110110: data <= 32'hb6dc2f84;
    11'b00000110111: data <= 32'hbb28400d;
    11'b00000111000: data <= 32'hbe7640d7;
    11'b00000111001: data <= 32'hbd9f3918;
    11'b00000111010: data <= 32'hb015bc86;
    11'b00000111011: data <= 32'h3a12bb52;
    11'b00000111100: data <= 32'h376337c5;
    11'b00000111101: data <= 32'h33203c7a;
    11'b00000111110: data <= 32'h3cf239f7;
    11'b00000111111: data <= 32'h40b8386b;
    11'b00001000000: data <= 32'h3e653a28;
    11'b00001000001: data <= 32'hb9373662;
    11'b00001000010: data <= 32'hbf19b9ec;
    11'b00001000011: data <= 32'hb85abdcb;
    11'b00001000100: data <= 32'h3cd3bc8f;
    11'b00001000101: data <= 32'h3d41bad3;
    11'b00001000110: data <= 32'h315cbd60;
    11'b00001000111: data <= 32'hb6ccbe00;
    11'b00001001000: data <= 32'hb161ae32;
    11'b00001001001: data <= 32'hb5333f08;
    11'b00001001010: data <= 32'hbd0d3f0a;
    11'b00001001011: data <= 32'hbf32b231;
    11'b00001001100: data <= 32'hbd0cbe5c;
    11'b00001001101: data <= 32'hb84fba1f;
    11'b00001001110: data <= 32'hb5de3b44;
    11'b00001001111: data <= 32'ha15f3d2a;
    11'b00001010000: data <= 32'h3cb63872;
    11'b00001010001: data <= 32'h40123728;
    11'b00001010010: data <= 32'h3c423d2b;
    11'b00001010011: data <= 32'hbb443e69;
    11'b00001010100: data <= 32'hbda838d4;
    11'b00001010101: data <= 32'h327bb901;
    11'b00001010110: data <= 32'h3f18bc2c;
    11'b00001010111: data <= 32'h3dbbbc73;
    11'b00001011000: data <= 32'h31bfbdcf;
    11'b00001011001: data <= 32'h2a7fbd70;
    11'b00001011010: data <= 32'h3b61adcf;
    11'b00001011011: data <= 32'h3b283cf6;
    11'b00001011100: data <= 32'hb8d13a93;
    11'b00001011101: data <= 32'hbfdabc0d;
    11'b00001011110: data <= 32'hbf99bf96;
    11'b00001011111: data <= 32'hbc56ba09;
    11'b00001100000: data <= 32'hb8cc394b;
    11'b00001100001: data <= 32'hb2d23802;
    11'b00001100010: data <= 32'h38dbb670;
    11'b00001100011: data <= 32'h3c5a2633;
    11'b00001100100: data <= 32'h32613efc;
    11'b00001100101: data <= 32'hbcf34136;
    11'b00001100110: data <= 32'hbd0e3e12;
    11'b00001100111: data <= 32'h34d8b049;
    11'b00001101000: data <= 32'h3da7ba1f;
    11'b00001101001: data <= 32'h3a9ab910;
    11'b00001101010: data <= 32'ha10cb962;
    11'b00001101011: data <= 32'h39b7b92d;
    11'b00001101100: data <= 32'h405d2e55;
    11'b00001101101: data <= 32'h401c3af5;
    11'b00001101110: data <= 32'h9c213598;
    11'b00001101111: data <= 32'hbf24bc6a;
    11'b00001110000: data <= 32'hbebabe97;
    11'b00001110001: data <= 32'hb8f2b9e7;
    11'b00001110010: data <= 32'hb15aab43;
    11'b00001110011: data <= 32'hb424ba8d;
    11'b00001110100: data <= 32'ha23fbe8a;
    11'b00001110101: data <= 32'h34c9b84d;
    11'b00001110110: data <= 32'hb3e53f40;
    11'b00001110111: data <= 32'hbd064195;
    11'b00001111000: data <= 32'hbd403ddf;
    11'b00001111001: data <= 32'hb4d9b3ec;
    11'b00001111010: data <= 32'h3405b7f4;
    11'b00001111011: data <= 32'hb49631a8;
    11'b00001111100: data <= 32'hb6b73521;
    11'b00001111101: data <= 32'h3c569e3f;
    11'b00001111110: data <= 32'h41a432ef;
    11'b00001111111: data <= 32'h40e73ab4;
    11'b00010000000: data <= 32'h31753998;
    11'b00010000001: data <= 32'hbd9db43c;
    11'b00010000010: data <= 32'hbaa8ba7d;
    11'b00010000011: data <= 32'h36b3b870;
    11'b00010000100: data <= 32'h37ffb9a8;
    11'b00010000101: data <= 32'hb2dfbf5f;
    11'b00010000110: data <= 32'hb45bc0d4;
    11'b00010000111: data <= 32'h349fbb53;
    11'b00010001000: data <= 32'h323b3ddc;
    11'b00010001001: data <= 32'hba004035;
    11'b00010001010: data <= 32'hbd7238a7;
    11'b00010001011: data <= 32'hbc97ba58;
    11'b00010001100: data <= 32'hbbfdb5b6;
    11'b00010001101: data <= 32'hbd253a05;
    11'b00010001110: data <= 32'hbaf239ea;
    11'b00010001111: data <= 32'h3b49ab96;
    11'b00010010000: data <= 32'h40f4a31c;
    11'b00010010001: data <= 32'h3f993c1e;
    11'b00010010010: data <= 32'hb07a3e6b;
    11'b00010010011: data <= 32'hbc373c18;
    11'b00010010100: data <= 32'h28e23292;
    11'b00010010101: data <= 32'h3cd3b241;
    11'b00010010110: data <= 32'h3a19ba82;
    11'b00010010111: data <= 32'hb4c2bfbd;
    11'b00010011000: data <= 32'hae91c098;
    11'b00010011001: data <= 32'h3c52bb2c;
    11'b00010011010: data <= 32'h3d653b9a;
    11'b00010011011: data <= 32'h2f523c45;
    11'b00010011100: data <= 32'hbce6b6f4;
    11'b00010011101: data <= 32'hbe63bcfb;
    11'b00010011110: data <= 32'hbe20b481;
    11'b00010011111: data <= 32'hbe583a43;
    11'b00010100000: data <= 32'hbc6e33bf;
    11'b00010100001: data <= 32'h3533bb84;
    11'b00010100010: data <= 32'h3dccb91d;
    11'b00010100011: data <= 32'h3aeb3ca3;
    11'b00010100100: data <= 32'hb8e840c8;
    11'b00010100101: data <= 32'hbaed3fb6;
    11'b00010100110: data <= 32'h36293a77;
    11'b00010100111: data <= 32'h3c8831a5;
    11'b00010101000: data <= 32'h33eab4b5;
    11'b00010101001: data <= 32'hb96abc60;
    11'b00010101010: data <= 32'h3345bdcb;
    11'b00010101011: data <= 32'h4034b895;
    11'b00010101100: data <= 32'h40ff3880;
    11'b00010101101: data <= 32'h3ae7360a;
    11'b00010101110: data <= 32'hbb2cba6e;
    11'b00010101111: data <= 32'hbd3bbc6d;
    11'b00010110000: data <= 32'hbc15ae18;
    11'b00010110001: data <= 32'hbc3d3658;
    11'b00010110010: data <= 32'hbc2dba9d;
    11'b00010110011: data <= 32'hb4c5c052;
    11'b00010110100: data <= 32'h3788bd88;
    11'b00010110101: data <= 32'h30c33c18;
    11'b00010110110: data <= 32'hba1840f2;
    11'b00010110111: data <= 32'hba2c3f64;
    11'b00010111000: data <= 32'h2e96392e;
    11'b00010111001: data <= 32'h336c35f1;
    11'b00010111010: data <= 32'hbacb3824;
    11'b00010111011: data <= 32'hbd2a2c04;
    11'b00010111100: data <= 32'h35a7b869;
    11'b00010111101: data <= 32'h4139b4ed;
    11'b00010111110: data <= 32'h41c336b7;
    11'b00010111111: data <= 32'h3c2a36b0;
    11'b00011000000: data <= 32'hb853b38a;
    11'b00011000001: data <= 32'hb729b4c2;
    11'b00011000010: data <= 32'h30fa34df;
    11'b00011000011: data <= 32'hb10d25d8;
    11'b00011000100: data <= 32'hbabebec9;
    11'b00011000101: data <= 32'hb91cc1e2;
    11'b00011000110: data <= 32'h3171bf43;
    11'b00011000111: data <= 32'h34f43937;
    11'b00011001000: data <= 32'hb4da3f0a;
    11'b00011001001: data <= 32'hb8d63ac2;
    11'b00011001010: data <= 32'hb711ae9d;
    11'b00011001011: data <= 32'hbac235b6;
    11'b00011001100: data <= 32'hbf753c99;
    11'b00011001101: data <= 32'hbf603a00;
    11'b00011001110: data <= 32'h2e8cb513;
    11'b00011001111: data <= 32'h4071b771;
    11'b00011010000: data <= 32'h4078368d;
    11'b00011010001: data <= 32'h387d3c09;
    11'b00011010010: data <= 32'hb54c3ae2;
    11'b00011010011: data <= 32'h376939f2;
    11'b00011010100: data <= 32'h3cc43a81;
    11'b00011010101: data <= 32'h365329be;
    11'b00011010110: data <= 32'hba99bee8;
    11'b00011010111: data <= 32'hb92fc183;
    11'b00011011000: data <= 32'h3927beaf;
    11'b00011011001: data <= 32'h3d023407;
    11'b00011011010: data <= 32'h38ae3983;
    11'b00011011011: data <= 32'hb487b668;
    11'b00011011100: data <= 32'hb9b9bac2;
    11'b00011011101: data <= 32'hbd3034ef;
    11'b00011011110: data <= 32'hc0413d54;
    11'b00011011111: data <= 32'hc006388b;
    11'b00011100000: data <= 32'hb674bbbc;
    11'b00011100001: data <= 32'h3ca6bc6a;
    11'b00011100010: data <= 32'h3bee3554;
    11'b00011100011: data <= 32'hb2363e52;
    11'b00011100100: data <= 32'hb48c3eaa;
    11'b00011100101: data <= 32'h3b823d5a;
    11'b00011100110: data <= 32'h3db63caf;
    11'b00011100111: data <= 32'h30233837;
    11'b00011101000: data <= 32'hbccdbad1;
    11'b00011101001: data <= 32'hb843bee5;
    11'b00011101010: data <= 32'h3dafbc54;
    11'b00011101011: data <= 32'h40922380;
    11'b00011101100: data <= 32'h3d67aef2;
    11'b00011101101: data <= 32'h2dbebc4b;
    11'b00011101110: data <= 32'hb6a5bbcc;
    11'b00011101111: data <= 32'hb9fc3776;
    11'b00011110000: data <= 32'hbdc93ca2;
    11'b00011110001: data <= 32'hbed8b381;
    11'b00011110010: data <= 32'hbb03c01c;
    11'b00011110011: data <= 32'h2df2bf88;
    11'b00011110100: data <= 32'ha5d12e7b;
    11'b00011110101: data <= 32'hb9093e6a;
    11'b00011110110: data <= 32'hb3e33e29;
    11'b00011110111: data <= 32'h3ade3c3e;
    11'b00011111000: data <= 32'h3a783cb0;
    11'b00011111001: data <= 32'hba873ccf;
    11'b00011111010: data <= 32'hbf6f361b;
    11'b00011111011: data <= 32'hb85ab850;
    11'b00011111100: data <= 32'h3f4db81f;
    11'b00011111101: data <= 32'h413ba97c;
    11'b00011111110: data <= 32'h3dccb41a;
    11'b00011111111: data <= 32'h34d8ba6b;
    11'b00100000000: data <= 32'h355bb56a;
    11'b00100000001: data <= 32'h37ed3b49;
    11'b00100000010: data <= 32'hb4633b9f;
    11'b00100000011: data <= 32'hbccfbbb6;
    11'b00100000100: data <= 32'hbc6cc18e;
    11'b00100000101: data <= 32'hb611c08b;
    11'b00100000110: data <= 32'hb179b1e7;
    11'b00100000111: data <= 32'hb5f53bbb;
    11'b00100001000: data <= 32'ha9d4379d;
    11'b00100001001: data <= 32'h38092bee;
    11'b00100001010: data <= 32'hae123adb;
    11'b00100001011: data <= 32'hbf103ed2;
    11'b00100001100: data <= 32'hc0cf3ce4;
    11'b00100001101: data <= 32'hba1e2344;
    11'b00100001110: data <= 32'h3de6b709;
    11'b00100001111: data <= 32'h3fa5ac36;
    11'b00100010000: data <= 32'h3a02303f;
    11'b00100010001: data <= 32'h336f2dcf;
    11'b00100010010: data <= 32'h3c713905;
    11'b00100010011: data <= 32'h3eaf3dc7;
    11'b00100010100: data <= 32'h38d33bfd;
    11'b00100010101: data <= 32'hbb5ebbfa;
    11'b00100010110: data <= 32'hbc66c114;
    11'b00100010111: data <= 32'haf04bfc9;
    11'b00100011000: data <= 32'h3853b560;
    11'b00100011001: data <= 32'h36c9261e;
    11'b00100011010: data <= 32'h352bbb30;
    11'b00100011011: data <= 32'h34dcbc04;
    11'b00100011100: data <= 32'hb820382a;
    11'b00100011101: data <= 32'hbff13f60;
    11'b00100011110: data <= 32'hc0dd3cf7;
    11'b00100011111: data <= 32'hbc40b60f;
    11'b00100100000: data <= 32'h3842bbb1;
    11'b00100100001: data <= 32'h3861b257;
    11'b00100100010: data <= 32'hb53138b8;
    11'b00100100011: data <= 32'ha6583aa5;
    11'b00100100100: data <= 32'h3e123cbf;
    11'b00100100101: data <= 32'h40343ed7;
    11'b00100100110: data <= 32'h38f13d4a;
    11'b00100100111: data <= 32'hbc97b30a;
    11'b00100101000: data <= 32'hbc24bd97;
    11'b00100101001: data <= 32'h382ebc33;
    11'b00100101010: data <= 32'h3de6b433;
    11'b00100101011: data <= 32'h3ca1b97e;
    11'b00100101100: data <= 32'h3932bf0d;
    11'b00100101101: data <= 32'h3800bdc0;
    11'b00100101110: data <= 32'ha95237f1;
    11'b00100101111: data <= 32'hbcd83ed4;
    11'b00100110000: data <= 32'hbf6638d5;
    11'b00100110001: data <= 32'hbcecbd58;
    11'b00100110010: data <= 32'hb703bed1;
    11'b00100110011: data <= 32'hb93bb6c4;
    11'b00100110100: data <= 32'hbc57394c;
    11'b00100110101: data <= 32'hb28c3a08;
    11'b00100110110: data <= 32'h3dd43aab;
    11'b00100110111: data <= 32'h3ea63ddb;
    11'b00100111000: data <= 32'hb1523eda;
    11'b00100111001: data <= 32'hbf0a3b47;
    11'b00100111010: data <= 32'hbc46a7ee;
    11'b00100111011: data <= 32'h3b6db078;
    11'b00100111100: data <= 32'h3f4fac5c;
    11'b00100111101: data <= 32'h3ccbbaa9;
    11'b00100111110: data <= 32'h394bbebb;
    11'b00100111111: data <= 32'h3bfabbf6;
    11'b00101000000: data <= 32'h3c663b01;
    11'b00101000001: data <= 32'h30493e2b;
    11'b00101000010: data <= 32'hbbe9ad78;
    11'b00101000011: data <= 32'hbcb7c01c;
    11'b00101000100: data <= 32'hbb19c01b;
    11'b00101000101: data <= 32'hbc05b871;
    11'b00101000110: data <= 32'hbc3c3390;
    11'b00101000111: data <= 32'hae18b2f8;
    11'b00101001000: data <= 32'h3c9bb52f;
    11'b00101001001: data <= 32'h3aab3a6b;
    11'b00101001010: data <= 32'hbc5b3fab;
    11'b00101001011: data <= 32'hc0903ed6;
    11'b00101001100: data <= 32'hbcbc39df;
    11'b00101001101: data <= 32'h39f43291;
    11'b00101001110: data <= 32'h3cd02893;
    11'b00101001111: data <= 32'h35bfb7df;
    11'b00101010000: data <= 32'h342fbb2a;
    11'b00101010001: data <= 32'h3de2ad58;
    11'b00101010010: data <= 32'h40703d93;
    11'b00101010011: data <= 32'h3cea3e1b;
    11'b00101010100: data <= 32'hb670b3b9;
    11'b00101010101: data <= 32'hbc06bf8c;
    11'b00101010110: data <= 32'hb942be6e;
    11'b00101010111: data <= 32'hb6d8b67f;
    11'b00101011000: data <= 32'hb595b69c;
    11'b00101011001: data <= 32'h3425be1e;
    11'b00101011010: data <= 32'h3b6bbe71;
    11'b00101011011: data <= 32'h35503039;
    11'b00101011100: data <= 32'hbd773f66;
    11'b00101011101: data <= 32'hc06e3f03;
    11'b00101011110: data <= 32'hbcdf3802;
    11'b00101011111: data <= 32'h2cd0b21a;
    11'b00101100000: data <= 32'hae1dac89;
    11'b00101100001: data <= 32'hbb7ca939;
    11'b00101100010: data <= 32'hb594af6d;
    11'b00101100011: data <= 32'h3e8f3830;
    11'b00101100100: data <= 32'h41533e62;
    11'b00101100101: data <= 32'h3db43e86;
    11'b00101100110: data <= 32'hb75c349a;
    11'b00101100111: data <= 32'hbb25ba7d;
    11'b00101101000: data <= 32'haa52b7fe;
    11'b00101101001: data <= 32'h380f2795;
    11'b00101101010: data <= 32'h36a9bae7;
    11'b00101101011: data <= 32'h3865c0ca;
    11'b00101101100: data <= 32'h3b9fc07f;
    11'b00101101101: data <= 32'h38b6aec9;
    11'b00101101110: data <= 32'hb94a3e87;
    11'b00101101111: data <= 32'hbdbf3c97;
    11'b00101110000: data <= 32'hbc1bb6c1;
    11'b00101110001: data <= 32'hb8f8bb8b;
    11'b00101110010: data <= 32'hbd29b475;
    11'b00101110011: data <= 32'hbfb130f4;
    11'b00101110100: data <= 32'hba4aa121;
    11'b00101110101: data <= 32'h3dda33b9;
    11'b00101110110: data <= 32'h40833cb9;
    11'b00101110111: data <= 32'h39af3eb6;
    11'b00101111000: data <= 32'hbc363c8e;
    11'b00101111001: data <= 32'hbb563859;
    11'b00101111010: data <= 32'h3706393e;
    11'b00101111011: data <= 32'h3c07382f;
    11'b00101111100: data <= 32'h383dbade;
    11'b00101111101: data <= 32'h36ccc0b2;
    11'b00101111110: data <= 32'h3c8dbfa2;
    11'b00101111111: data <= 32'h3dd43301;
    11'b00110000000: data <= 32'h39513dd2;
    11'b00110000001: data <= 32'hb5243683;
    11'b00110000010: data <= 32'hb922bd04;
    11'b00110000011: data <= 32'hbb18bd75;
    11'b00110000100: data <= 32'hbeb5b4f2;
    11'b00110000101: data <= 32'hc01218a8;
    11'b00110000110: data <= 32'hba30b9c6;
    11'b00110000111: data <= 32'h3c8abb1b;
    11'b00110001000: data <= 32'h3d9a3443;
    11'b00110001001: data <= 32'hb4b33e1b;
    11'b00110001010: data <= 32'hbe903ee7;
    11'b00110001011: data <= 32'hbbb13d60;
    11'b00110001100: data <= 32'h37c93cb6;
    11'b00110001101: data <= 32'h38fd3a2f;
    11'b00110001110: data <= 32'hb45bb796;
    11'b00110001111: data <= 32'hb2ddbe38;
    11'b00110010000: data <= 32'h3cfebb97;
    11'b00110010001: data <= 32'h40b03a5c;
    11'b00110010010: data <= 32'h3f2c3d94;
    11'b00110010011: data <= 32'h37a82ba4;
    11'b00110010100: data <= 32'hb451bd39;
    11'b00110010101: data <= 32'hb8afbbbb;
    11'b00110010110: data <= 32'hbc702b5a;
    11'b00110010111: data <= 32'hbd43b4aa;
    11'b00110011000: data <= 32'hb613bf29;
    11'b00110011001: data <= 32'h3b16c069;
    11'b00110011010: data <= 32'h39f6b92c;
    11'b00110011011: data <= 32'hba2d3cd8;
    11'b00110011100: data <= 32'hbe8c3eab;
    11'b00110011101: data <= 32'hba763c89;
    11'b00110011110: data <= 32'h30fb3a87;
    11'b00110011111: data <= 32'hb6e13941;
    11'b00110100000: data <= 32'hbe61a00c;
    11'b00110100001: data <= 32'hbc59b93e;
    11'b00110100010: data <= 32'h3c83b130;
    11'b00110100011: data <= 32'h414f3c49;
    11'b00110100100: data <= 32'h400c3d62;
    11'b00110100101: data <= 32'h38023464;
    11'b00110100110: data <= 32'haff5b796;
    11'b00110100111: data <= 32'h291e313a;
    11'b00110101000: data <= 32'had713a20;
    11'b00110101001: data <= 32'hb656b6c0;
    11'b00110101010: data <= 32'h9cb4c0ff;
    11'b00110101011: data <= 32'h3a59c1c7;
    11'b00110101100: data <= 32'h39bdbc0b;
    11'b00110101101: data <= 32'hb4ef3b4c;
    11'b00110101110: data <= 32'hbaca3c20;
    11'b00110101111: data <= 32'hb58430c2;
    11'b00110110000: data <= 32'hb279aba0;
    11'b00110110001: data <= 32'hbdcc35d1;
    11'b00110110010: data <= 32'hc1473459;
    11'b00110110011: data <= 32'hbecab4c0;
    11'b00110110100: data <= 32'h3a8eb296;
    11'b00110110101: data <= 32'h40663957;
    11'b00110110110: data <= 32'h3d143c8a;
    11'b00110110111: data <= 32'hb1b13a3b;
    11'b00110111000: data <= 32'hb3243988;
    11'b00110111001: data <= 32'h38b33d8a;
    11'b00110111010: data <= 32'h39113de5;
    11'b00110111011: data <= 32'haa6db390;
    11'b00110111100: data <= 32'hae0fc0c4;
    11'b00110111101: data <= 32'h39f7c111;
    11'b00110111110: data <= 32'h3cf7b924;
    11'b00110111111: data <= 32'h3a873a4e;
    11'b00111000000: data <= 32'h356533e3;
    11'b00111000001: data <= 32'h34a5baf9;
    11'b00111000010: data <= 32'hb3b6b9a0;
    11'b00111000011: data <= 32'hbeff3469;
    11'b00111000100: data <= 32'hc186351e;
    11'b00111000101: data <= 32'hbec2b969;
    11'b00111000110: data <= 32'h3817bc7e;
    11'b00111000111: data <= 32'h3d38b501;
    11'b00111001000: data <= 32'h2eb639ae;
    11'b00111001001: data <= 32'hbbcb3c66;
    11'b00111001010: data <= 32'hb57a3d8c;
    11'b00111001011: data <= 32'h3a6a3fc8;
    11'b00111001100: data <= 32'h38833f21;
    11'b00111001101: data <= 32'hb90e315d;
    11'b00111001110: data <= 32'hba49be34;
    11'b00111001111: data <= 32'h3899bdc2;
    11'b00111010000: data <= 32'h3f552fcb;
    11'b00111010001: data <= 32'h3f4c3a81;
    11'b00111010010: data <= 32'h3cccb39a;
    11'b00111010011: data <= 32'h3a38bcdf;
    11'b00111010100: data <= 32'h300bb843;
    11'b00111010101: data <= 32'hbc8d3963;
    11'b00111010110: data <= 32'hbfc134d7;
    11'b00111010111: data <= 32'hbc8abdbb;
    11'b00111011000: data <= 32'h3596c09c;
    11'b00111011001: data <= 32'h384dbd3b;
    11'b00111011010: data <= 32'hb9313339;
    11'b00111011011: data <= 32'hbcd13b69;
    11'b00111011100: data <= 32'hb1d03c82;
    11'b00111011101: data <= 32'h39db3e0e;
    11'b00111011110: data <= 32'hb16a3e2f;
    11'b00111011111: data <= 32'hbf393873;
    11'b00111100000: data <= 32'hbf02b87b;
    11'b00111100001: data <= 32'h33bcb65a;
    11'b00111100010: data <= 32'h3fec391f;
    11'b00111100011: data <= 32'h3ffc3a45;
    11'b00111100100: data <= 32'h3cc3b435;
    11'b00111100101: data <= 32'h3ad3b9ab;
    11'b00111100110: data <= 32'h399136f7;
    11'b00111100111: data <= 32'ha8dc3dea;
    11'b00111101000: data <= 32'hba4836a8;
    11'b00111101001: data <= 32'hb823bfc2;
    11'b00111101010: data <= 32'h34dcc1d7;
    11'b00111101011: data <= 32'h34b3beb6;
    11'b00111101100: data <= 32'hb80eabaa;
    11'b00111101101: data <= 32'hb8c13503;
    11'b00111101110: data <= 32'h35f52ccc;
    11'b00111101111: data <= 32'h391b36ef;
    11'b00111110000: data <= 32'hbba93c12;
    11'b00111110001: data <= 32'hc18c3a25;
    11'b00111110010: data <= 32'hc0cea233;
    11'b00111110011: data <= 32'haf21afc5;
    11'b00111110100: data <= 32'h3e0a36f2;
    11'b00111110101: data <= 32'h3cb737f5;
    11'b00111110110: data <= 32'h356ba82c;
    11'b00111110111: data <= 32'h38533271;
    11'b00111111000: data <= 32'h3ca83e4d;
    11'b00111111001: data <= 32'h3ac44084;
    11'b00111111010: data <= 32'hb006399d;
    11'b00111111011: data <= 32'hb631bf13;
    11'b00111111100: data <= 32'h3292c103;
    11'b00111111101: data <= 32'h385bbcb0;
    11'b00111111110: data <= 32'h35779b72;
    11'b00111111111: data <= 32'h3801b653;
    11'b01000000000: data <= 32'h3c6cbc5c;
    11'b01000000001: data <= 32'h3a01b81c;
    11'b01000000010: data <= 32'hbca63988;
    11'b01000000011: data <= 32'hc1af3ab0;
    11'b01000000100: data <= 32'hc099b01e;
    11'b01000000101: data <= 32'hb482b9f9;
    11'b01000000110: data <= 32'h396fb707;
    11'b01000000111: data <= 32'haf69a92f;
    11'b01000001000: data <= 32'hb9fa2e0b;
    11'b01000001001: data <= 32'h317c3a25;
    11'b01000001010: data <= 32'h3d7b402d;
    11'b01000001011: data <= 32'h3c184109;
    11'b01000001100: data <= 32'hb66f3c12;
    11'b01000001101: data <= 32'hbb96bbd5;
    11'b01000001110: data <= 32'had1abd2e;
    11'b01000001111: data <= 32'h3b48b05f;
    11'b01000010000: data <= 32'h3cc03462;
    11'b01000010001: data <= 32'h3d49bac9;
    11'b01000010010: data <= 32'h3e5ebeab;
    11'b01000010011: data <= 32'h3c58b945;
    11'b01000010100: data <= 32'hb8923b78;
    11'b01000010101: data <= 32'hbfab3b60;
    11'b01000010110: data <= 32'hbdffb91b;
    11'b01000010111: data <= 32'hb25cbef4;
    11'b01000011000: data <= 32'ha974bd92;
    11'b01000011001: data <= 32'hbc58b88c;
    11'b01000011010: data <= 32'hbd35aecb;
    11'b01000011011: data <= 32'h30c337fb;
    11'b01000011100: data <= 32'h3d8a3e48;
    11'b01000011101: data <= 32'h385d4025;
    11'b01000011110: data <= 32'hbd713cb9;
    11'b01000011111: data <= 32'hbf78a94c;
    11'b01000100000: data <= 32'hb7dbaa2c;
    11'b01000100001: data <= 32'h3bd039b3;
    11'b01000100010: data <= 32'h3d483746;
    11'b01000100011: data <= 32'h3cf9bb7b;
    11'b01000100100: data <= 32'h3e04bdaa;
    11'b01000100101: data <= 32'h3dda2c86;
    11'b01000100110: data <= 32'h37a13eb8;
    11'b01000100111: data <= 32'hb8973c8c;
    11'b01000101000: data <= 32'hb864bc12;
    11'b01000101001: data <= 32'ha133c091;
    11'b01000101010: data <= 32'hb52fbed9;
    11'b01000101011: data <= 32'hbcd0b9f1;
    11'b01000101100: data <= 32'hbba1b891;
    11'b01000101101: data <= 32'h3901b812;
    11'b01000101110: data <= 32'h3d9e3513;
    11'b01000101111: data <= 32'had103ce2;
    11'b01000110000: data <= 32'hc0783c92;
    11'b01000110001: data <= 32'hc0f7382c;
    11'b01000110010: data <= 32'hba4737c9;
    11'b01000110011: data <= 32'h38d23a5b;
    11'b01000110100: data <= 32'h38443458;
    11'b01000110101: data <= 32'h33a2ba8f;
    11'b01000110110: data <= 32'h3b1cb997;
    11'b01000110111: data <= 32'h3eb63c5e;
    11'b01000111000: data <= 32'h3d6c40df;
    11'b01000111001: data <= 32'h35773da6;
    11'b01000111010: data <= 32'haebabb24;
    11'b01000111011: data <= 32'h26f4bf86;
    11'b01000111100: data <= 32'hb1cabc4d;
    11'b01000111101: data <= 32'hb891b6a4;
    11'b01000111110: data <= 32'h9a14bc24;
    11'b01000111111: data <= 32'h3d5fbea2;
    11'b01001000000: data <= 32'h3e32bb0a;
    11'b01001000001: data <= 32'hb480387a;
    11'b01001000010: data <= 32'hc0983c28;
    11'b01001000011: data <= 32'hc08b37f5;
    11'b01001000100: data <= 32'hb9cd2e24;
    11'b01001000101: data <= 32'h9fb12e0f;
    11'b01001000110: data <= 32'hb9efb3ea;
    11'b01001000111: data <= 32'hbc5bba16;
    11'b01001001000: data <= 32'h317db1c1;
    11'b01001001001: data <= 32'h3eba3e57;
    11'b01001001010: data <= 32'h3e6e413d;
    11'b01001001011: data <= 32'h35083e2f;
    11'b01001001100: data <= 32'hb758b4ad;
    11'b01001001101: data <= 32'hb32eb982;
    11'b01001001110: data <= 32'h2de5321d;
    11'b01001001111: data <= 32'h31f932d2;
    11'b01001010000: data <= 32'h3a43bd0f;
    11'b01001010001: data <= 32'h3f1fc095;
    11'b01001010010: data <= 32'h3f05bd24;
    11'b01001010011: data <= 32'h31113878;
    11'b01001010100: data <= 32'hbd8c3c44;
    11'b01001010101: data <= 32'hbd092de2;
    11'b01001010110: data <= 32'hb4c9ba29;
    11'b01001010111: data <= 32'hb7e8ba6f;
    11'b01001011000: data <= 32'hbf05ba04;
    11'b01001011001: data <= 32'hbfa9bb16;
    11'b01001011010: data <= 32'hb01bb569;
    11'b01001011011: data <= 32'h3e6c3c53;
    11'b01001011100: data <= 32'h3cf03ff0;
    11'b01001011101: data <= 32'hb7cb3d8b;
    11'b01001011110: data <= 32'hbd33368b;
    11'b01001011111: data <= 32'hb90638bc;
    11'b01001100000: data <= 32'h31e53d48;
    11'b01001100001: data <= 32'h363339a0;
    11'b01001100010: data <= 32'h39bdbcea;
    11'b01001100011: data <= 32'h3e26c048;
    11'b01001100100: data <= 32'h3f5eb9ec;
    11'b01001100101: data <= 32'h3bd33cca;
    11'b01001100110: data <= 32'ha4533d1c;
    11'b01001100111: data <= 32'ha5f9b45d;
    11'b01001101000: data <= 32'h333fbd5f;
    11'b01001101001: data <= 32'hb8fabc87;
    11'b01001101010: data <= 32'hbfe0ba76;
    11'b01001101011: data <= 32'hbf1cbc6b;
    11'b01001101100: data <= 32'h32a2bc8b;
    11'b01001101101: data <= 32'h3e76b226;
    11'b01001101110: data <= 32'h393d3acd;
    11'b01001101111: data <= 32'hbd663bee;
    11'b01001110000: data <= 32'hbfaa3a55;
    11'b01001110001: data <= 32'hbab83cdf;
    11'b01001110010: data <= 32'h1dba3e90;
    11'b01001110011: data <= 32'hb2ea399a;
    11'b01001110100: data <= 32'hb4d1bc5b;
    11'b01001110101: data <= 32'h393bbdf5;
    11'b01001110110: data <= 32'h3ec8338f;
    11'b01001110111: data <= 32'h3ea03fca;
    11'b01001111000: data <= 32'h3be03e03;
    11'b01001111001: data <= 32'h397fb4ae;
    11'b01001111010: data <= 32'h37cdbc5f;
    11'b01001111011: data <= 32'hb6e8b7d2;
    11'b01001111100: data <= 32'hbdabb399;
    11'b01001111101: data <= 32'hbb3ebce0;
    11'b01001111110: data <= 32'h3b39c026;
    11'b01001111111: data <= 32'h3ef1bde0;
    11'b01010000000: data <= 32'h35abae79;
    11'b01010000001: data <= 32'hbe2538f7;
    11'b01010000010: data <= 32'hbed43987;
    11'b01010000011: data <= 32'hb88d3b5d;
    11'b01010000100: data <= 32'hb4723c3a;
    11'b01010000101: data <= 32'hbd1f3333;
    11'b01010000110: data <= 32'hbecfbc16;
    11'b01010000111: data <= 32'hb5e3bb50;
    11'b01010001000: data <= 32'h3d923a97;
    11'b01010001001: data <= 32'h3f344047;
    11'b01010001010: data <= 32'h3c3b3dda;
    11'b01010001011: data <= 32'h37d12360;
    11'b01010001100: data <= 32'h3500ae8f;
    11'b01010001101: data <= 32'hb1003ac3;
    11'b01010001110: data <= 32'hb91f399c;
    11'b01010001111: data <= 32'haaecbc75;
    11'b01010010000: data <= 32'h3d70c125;
    11'b01010010001: data <= 32'h3f3bbfec;
    11'b01010010010: data <= 32'h384fb4c4;
    11'b01010010011: data <= 32'hba86383b;
    11'b01010010100: data <= 32'hb914346f;
    11'b01010010101: data <= 32'h313b2c30;
    11'b01010010110: data <= 32'hb6aa2ff1;
    11'b01010010111: data <= 32'hc048b4d9;
    11'b01010011000: data <= 32'hc147bc36;
    11'b01010011001: data <= 32'hbb38badf;
    11'b01010011010: data <= 32'h3c9c37f3;
    11'b01010011011: data <= 32'h3d9e3dd6;
    11'b01010011100: data <= 32'h34ae3c0a;
    11'b01010011101: data <= 32'hb59a35d4;
    11'b01010011110: data <= 32'haeff3c0e;
    11'b01010011111: data <= 32'h9d09402e;
    11'b01010100000: data <= 32'hb44e3dd8;
    11'b01010100001: data <= 32'h296ebaf3;
    11'b01010100010: data <= 32'h3c5cc0c1;
    11'b01010100011: data <= 32'h3e83bdf7;
    11'b01010100100: data <= 32'h3c0f34ca;
    11'b01010100101: data <= 32'h362139ef;
    11'b01010100110: data <= 32'h39c4afdb;
    11'b01010100111: data <= 32'h3be9b917;
    11'b01010101000: data <= 32'hb4adb591;
    11'b01010101001: data <= 32'hc094b5ab;
    11'b01010101010: data <= 32'hc127bc2c;
    11'b01010101011: data <= 32'hb934bd54;
    11'b01010101100: data <= 32'h3c8bb8d1;
    11'b01010101101: data <= 32'h3a6832a3;
    11'b01010101110: data <= 32'hb94d34b8;
    11'b01010101111: data <= 32'hbc5c3756;
    11'b01010110000: data <= 32'hb55d3e39;
    11'b01010110001: data <= 32'h1b574104;
    11'b01010110010: data <= 32'hb89c3e5b;
    11'b01010110011: data <= 32'hba65b957;
    11'b01010110100: data <= 32'h2e71bed4;
    11'b01010110101: data <= 32'h3c9cb744;
    11'b01010110110: data <= 32'h3d833c99;
    11'b01010110111: data <= 32'h3d233bf2;
    11'b01010111000: data <= 32'h3e33b4a1;
    11'b01010111001: data <= 32'h3db9b933;
    11'b01010111010: data <= 32'h0bd12fb0;
    11'b01010111011: data <= 32'hbedc34df;
    11'b01010111100: data <= 32'hbeb3baae;
    11'b01010111101: data <= 32'h2f8dbfc3;
    11'b01010111110: data <= 32'h3d26bf0f;
    11'b01010111111: data <= 32'h3635bb0b;
    11'b01011000000: data <= 32'hbc52b4e4;
    11'b01011000001: data <= 32'hbc3732bf;
    11'b01011000010: data <= 32'h15773cea;
    11'b01011000011: data <= 32'h25b43fb3;
    11'b01011000100: data <= 32'hbd3c3c4d;
    11'b01011000101: data <= 32'hc027b905;
    11'b01011000110: data <= 32'hbc47bc2f;
    11'b01011000111: data <= 32'h389f3558;
    11'b01011001000: data <= 32'h3d513e0a;
    11'b01011001001: data <= 32'h3d473b4c;
    11'b01011001010: data <= 32'h3d8bb41b;
    11'b01011001011: data <= 32'h3d0c2416;
    11'b01011001100: data <= 32'h34393d49;
    11'b01011001101: data <= 32'hbaff3d94;
    11'b01011001110: data <= 32'hb938b6d5;
    11'b01011001111: data <= 32'h39eac069;
    11'b01011010000: data <= 32'h3d61c074;
    11'b01011010001: data <= 32'h354bbc95;
    11'b01011010010: data <= 32'hb95eb74f;
    11'b01011010011: data <= 32'hafb9b300;
    11'b01011010100: data <= 32'h3b0d3537;
    11'b01011010101: data <= 32'h32953ad4;
    11'b01011010110: data <= 32'hbf9f364a;
    11'b01011010111: data <= 32'hc1e8b958;
    11'b01011011000: data <= 32'hbed1ba46;
    11'b01011011001: data <= 32'h331734da;
    11'b01011011010: data <= 32'h3b0a3bd5;
    11'b01011011011: data <= 32'h381c3533;
    11'b01011011100: data <= 32'h3718b380;
    11'b01011011101: data <= 32'h39a53aca;
    11'b01011011110: data <= 32'h36394100;
    11'b01011011111: data <= 32'hb54d4092;
    11'b01011100000: data <= 32'hb46ea18c;
    11'b01011100001: data <= 32'h390cbfac;
    11'b01011100010: data <= 32'h3c36becd;
    11'b01011100011: data <= 32'h37c1b7b6;
    11'b01011100100: data <= 32'h3368b082;
    11'b01011100101: data <= 32'h3ca7b8b3;
    11'b01011100110: data <= 32'h3f72b823;
    11'b01011100111: data <= 32'h38642fd5;
    11'b01011101000: data <= 32'hbfae3162;
    11'b01011101001: data <= 32'hc1b6b898;
    11'b01011101010: data <= 32'hbdb3bb9b;
    11'b01011101011: data <= 32'h3448b7de;
    11'b01011101100: data <= 32'h34cdb22c;
    11'b01011101101: data <= 32'hb877b880;
    11'b01011101110: data <= 32'hb843b66a;
    11'b01011101111: data <= 32'h34c73ce4;
    11'b01011110000: data <= 32'h373041c6;
    11'b01011110001: data <= 32'hb5b240da;
    11'b01011110010: data <= 32'hba8031a4;
    11'b01011110011: data <= 32'hb43fbd01;
    11'b01011110100: data <= 32'h3663b883;
    11'b01011110101: data <= 32'h387138a0;
    11'b01011110110: data <= 32'h3b7834aa;
    11'b01011110111: data <= 32'h3fdcba39;
    11'b01011111000: data <= 32'h40baba48;
    11'b01011111001: data <= 32'h3b0d3492;
    11'b01011111010: data <= 32'hbd4e39b9;
    11'b01011111011: data <= 32'hbf7ab249;
    11'b01011111100: data <= 32'hb79dbcfc;
    11'b01011111101: data <= 32'h38b9bdb8;
    11'b01011111110: data <= 32'haf6fbd06;
    11'b01011111111: data <= 32'hbcd0bd11;
    11'b01100000000: data <= 32'hba5eb9f8;
    11'b01100000001: data <= 32'h38063ac8;
    11'b01100000010: data <= 32'h38f34078;
    11'b01100000011: data <= 32'hba2a3f13;
    11'b01100000100: data <= 32'hbf5f2c19;
    11'b01100000101: data <= 32'hbda2b8ca;
    11'b01100000110: data <= 32'hb51336d9;
    11'b01100000111: data <= 32'h35a63cee;
    11'b01100001000: data <= 32'h3b1e35ce;
    11'b01100001001: data <= 32'h3effbaf6;
    11'b01100001010: data <= 32'h402fb6e9;
    11'b01100001011: data <= 32'h3c173ce7;
    11'b01100001100: data <= 32'hb7f83f17;
    11'b01100001101: data <= 32'hb9503613;
    11'b01100001110: data <= 32'h36e6bd3d;
    11'b01100001111: data <= 32'h3a8cbf20;
    11'b01100010000: data <= 32'hb455bdf2;
    11'b01100010001: data <= 32'hbc62bd79;
    11'b01100010010: data <= 32'hb058bc62;
    11'b01100010011: data <= 32'h3d5aaa2f;
    11'b01100010100: data <= 32'h3be03c01;
    11'b01100010101: data <= 32'hbc813a81;
    11'b01100010110: data <= 32'hc12ab126;
    11'b01100010111: data <= 32'hc00cb443;
    11'b01100011000: data <= 32'hb96a397e;
    11'b01100011001: data <= 32'hac663be4;
    11'b01100011010: data <= 32'h2cfeb12a;
    11'b01100011011: data <= 32'h3957bc21;
    11'b01100011100: data <= 32'h3d253048;
    11'b01100011101: data <= 32'h3bac407d;
    11'b01100011110: data <= 32'h2dd8414f;
    11'b01100011111: data <= 32'ha29e3acd;
    11'b01100100000: data <= 32'h38f6bbf3;
    11'b01100100001: data <= 32'h38e7bceb;
    11'b01100100010: data <= 32'hb4b6b9a7;
    11'b01100100011: data <= 32'hb7a5baaf;
    11'b01100100100: data <= 32'h3bbebd22;
    11'b01100100101: data <= 32'h40a3bb5a;
    11'b01100100110: data <= 32'h3db5214b;
    11'b01100100111: data <= 32'hbc3e3479;
    11'b01100101000: data <= 32'hc0e0b1de;
    11'b01100101001: data <= 32'hbe9db457;
    11'b01100101010: data <= 32'hb75331fd;
    11'b01100101011: data <= 32'hb7d923c1;
    11'b01100101100: data <= 32'hbc0cbc37;
    11'b01100101101: data <= 32'hb868bd59;
    11'b01100101110: data <= 32'h38863613;
    11'b01100101111: data <= 32'h3aff4121;
    11'b01100110000: data <= 32'h32914177;
    11'b01100110001: data <= 32'hb3e63b4f;
    11'b01100110010: data <= 32'haab1b739;
    11'b01100110011: data <= 32'ha919acee;
    11'b01100110100: data <= 32'hb63c389e;
    11'b01100110101: data <= 32'h2b09ade8;
    11'b01100110110: data <= 32'h3ebfbd3a;
    11'b01100110111: data <= 32'h4192bd34;
    11'b01100111000: data <= 32'h3ec3b01e;
    11'b01100111001: data <= 32'hb86838a0;
    11'b01100111010: data <= 32'hbdb931a8;
    11'b01100111011: data <= 32'hb802b62d;
    11'b01100111100: data <= 32'h3139b85d;
    11'b01100111101: data <= 32'hb9d2bb99;
    11'b01100111110: data <= 32'hbefebf00;
    11'b01100111111: data <= 32'hbc74bead;
    11'b01101000000: data <= 32'h37f2299f;
    11'b01101000001: data <= 32'h3bff3f8c;
    11'b01101000010: data <= 32'ha6a03f94;
    11'b01101000011: data <= 32'hbc2d3836;
    11'b01101000100: data <= 32'hbc50254d;
    11'b01101000101: data <= 32'hba273bee;
    11'b01101000110: data <= 32'hb9113e1c;
    11'b01101000111: data <= 32'h1abd3462;
    11'b01101001000: data <= 32'h3dc3bd4d;
    11'b01101001001: data <= 32'h40bcbc7d;
    11'b01101001010: data <= 32'h3e5d3873;
    11'b01101001011: data <= 32'h2edc3dfb;
    11'b01101001100: data <= 32'hb11f3a37;
    11'b01101001101: data <= 32'h3996b5c2;
    11'b01101001110: data <= 32'h39a2babf;
    11'b01101001111: data <= 32'hba3cbc93;
    11'b01101010000: data <= 32'hbf37bef7;
    11'b01101010001: data <= 32'hb9cebf4b;
    11'b01101010010: data <= 32'h3caab99c;
    11'b01101010011: data <= 32'h3d8e38c2;
    11'b01101010100: data <= 32'hb41f393f;
    11'b01101010101: data <= 32'hbebfa635;
    11'b01101010110: data <= 32'hbe99332d;
    11'b01101010111: data <= 32'hbc3c3d99;
    11'b01101011000: data <= 32'hbb513e46;
    11'b01101011001: data <= 32'hb97dab38;
    11'b01101011010: data <= 32'h34edbe02;
    11'b01101011011: data <= 32'h3d2db9a3;
    11'b01101011100: data <= 32'h3ccb3dc5;
    11'b01101011101: data <= 32'h386140a6;
    11'b01101011110: data <= 32'h39093cdb;
    11'b01101011111: data <= 32'h3cc2b013;
    11'b01101100000: data <= 32'h39cdb60d;
    11'b01101100001: data <= 32'hba64b51c;
    11'b01101100010: data <= 32'hbd64bbc0;
    11'b01101100011: data <= 32'h32e3bec8;
    11'b01101100100: data <= 32'h402bbda4;
    11'b01101100101: data <= 32'h3f50b82d;
    11'b01101100110: data <= 32'hb311b238;
    11'b01101100111: data <= 32'hbe5db4ea;
    11'b01101101000: data <= 32'hbcf53219;
    11'b01101101001: data <= 32'hb9113c48;
    11'b01101101010: data <= 32'hbc303a50;
    11'b01101101011: data <= 32'hbe75baf6;
    11'b01101101100: data <= 32'hbc1abf4c;
    11'b01101101101: data <= 32'h33f0b7a7;
    11'b01101101110: data <= 32'h3a923f19;
    11'b01101101111: data <= 32'h38d440bc;
    11'b01101110000: data <= 32'h388a3c71;
    11'b01101110001: data <= 32'h39e93142;
    11'b01101110010: data <= 32'h319438fd;
    11'b01101110011: data <= 32'hbb663c48;
    11'b01101110100: data <= 32'hbb012e5a;
    11'b01101110101: data <= 32'h3b50bd9a;
    11'b01101110110: data <= 32'h410abed3;
    11'b01101110111: data <= 32'h3fdebaa8;
    11'b01101111000: data <= 32'h2d67b0bf;
    11'b01101111001: data <= 32'hb9bbad32;
    11'b01101111010: data <= 32'h21182eea;
    11'b01101111011: data <= 32'h34d836eb;
    11'b01101111100: data <= 32'hbba4afe7;
    11'b01101111101: data <= 32'hc07cbe2c;
    11'b01101111110: data <= 32'hbf06c026;
    11'b01101111111: data <= 32'hae8ab944;
    11'b01110000000: data <= 32'h3a303cd5;
    11'b01110000001: data <= 32'h364c3dc6;
    11'b01110000010: data <= 32'haee736d0;
    11'b01110000011: data <= 32'hb27334f1;
    11'b01110000100: data <= 32'hb8423e47;
    11'b01110000101: data <= 32'hbc84405f;
    11'b01110000110: data <= 32'hba933a2f;
    11'b01110000111: data <= 32'h3a0ebcd3;
    11'b01110001000: data <= 32'h4010be1e;
    11'b01110001001: data <= 32'h3e64b498;
    11'b01110001010: data <= 32'h36da392f;
    11'b01110001011: data <= 32'h36d437ca;
    11'b01110001100: data <= 32'h3d7d3015;
    11'b01110001101: data <= 32'h3cb02d05;
    11'b01110001110: data <= 32'hba0db625;
    11'b01110001111: data <= 32'hc08dbdee;
    11'b01110010000: data <= 32'hbe16bfff;
    11'b01110010001: data <= 32'h368fbc73;
    11'b01110010010: data <= 32'h3c7129ad;
    11'b01110010011: data <= 32'h31a529ca;
    11'b01110010100: data <= 32'hba19b77e;
    11'b01110010101: data <= 32'hba853363;
    11'b01110010110: data <= 32'hba523fbe;
    11'b01110010111: data <= 32'hbce740c8;
    11'b01110011000: data <= 32'hbd053918;
    11'b01110011001: data <= 32'hb409bd35;
    11'b01110011010: data <= 32'h3a77bc89;
    11'b01110011011: data <= 32'h3adb3896;
    11'b01110011100: data <= 32'h38823df8;
    11'b01110011101: data <= 32'h3ca03b41;
    11'b01110011110: data <= 32'h4015332c;
    11'b01110011111: data <= 32'h3db53544;
    11'b01110100000: data <= 32'hb9493530;
    11'b01110100001: data <= 32'hbf5fb89b;
    11'b01110100010: data <= 32'hb919be1f;
    11'b01110100011: data <= 32'h3d43be04;
    11'b01110100100: data <= 32'h3e2abbfe;
    11'b01110100101: data <= 32'h2fbebbf7;
    11'b01110100110: data <= 32'hbab2bc1a;
    11'b01110100111: data <= 32'hb815296d;
    11'b01110101000: data <= 32'hb40a3e7d;
    11'b01110101001: data <= 32'hbc293eca;
    11'b01110101010: data <= 32'hbf76b040;
    11'b01110101011: data <= 32'hbe01be77;
    11'b01110101100: data <= 32'hb6fdbad1;
    11'b01110101101: data <= 32'h315e3c23;
    11'b01110101110: data <= 32'h36c63e84;
    11'b01110101111: data <= 32'h3c6739bc;
    11'b01110110000: data <= 32'h3ed1336f;
    11'b01110110001: data <= 32'h3ba73c1b;
    11'b01110110010: data <= 32'hba2a3e7e;
    11'b01110110011: data <= 32'hbd5e398b;
    11'b01110110100: data <= 32'h30e0bb2a;
    11'b01110110101: data <= 32'h3f56be42;
    11'b01110110110: data <= 32'h3e7abd35;
    11'b01110110111: data <= 32'h31dcbc5d;
    11'b01110111000: data <= 32'hb3c7bb65;
    11'b01110111001: data <= 32'h392bacd8;
    11'b01110111010: data <= 32'h3b083bd1;
    11'b01110111011: data <= 32'hb8bf39d5;
    11'b01110111100: data <= 32'hc075bb03;
    11'b01110111101: data <= 32'hc06cbf54;
    11'b01110111110: data <= 32'hbba4baa7;
    11'b01110111111: data <= 32'haaf239c4;
    11'b01111000000: data <= 32'h30b83a66;
    11'b01111000001: data <= 32'h36e3b0d4;
    11'b01111000010: data <= 32'h39f32510;
    11'b01111000011: data <= 32'h32513ec2;
    11'b01111000100: data <= 32'hbbaf416b;
    11'b01111000101: data <= 32'hbc863e3b;
    11'b01111000110: data <= 32'h3309b7a1;
    11'b01111000111: data <= 32'h3dc6bd23;
    11'b01111001000: data <= 32'h3c59ba23;
    11'b01111001001: data <= 32'h31c3b4fc;
    11'b01111001010: data <= 32'h38dfb54a;
    11'b01111001011: data <= 32'h3fe4ab58;
    11'b01111001100: data <= 32'h3fd7380c;
    11'b01111001101: data <= 32'hb0033460;
    11'b01111001110: data <= 32'hc03dbb58;
    11'b01111001111: data <= 32'hbff2be7b;
    11'b01111010000: data <= 32'hb7f2bbaf;
    11'b01111010001: data <= 32'h345ab0e2;
    11'b01111010010: data <= 32'hac8ab876;
    11'b01111010011: data <= 32'hb4e7bd15;
    11'b01111010100: data <= 32'ha836b5d7;
    11'b01111010101: data <= 32'hb14f3f82;
    11'b01111010110: data <= 32'hbba541d8;
    11'b01111010111: data <= 32'hbd143e0d;
    11'b01111011000: data <= 32'hb80ab823;
    11'b01111011001: data <= 32'h3445bb01;
    11'b01111011010: data <= 32'h2f5030cb;
    11'b01111011011: data <= 32'ha52d394f;
    11'b01111011100: data <= 32'h3c863232;
    11'b01111011101: data <= 32'h414da765;
    11'b01111011110: data <= 32'h40b037fe;
    11'b01111011111: data <= 32'h2cc539ad;
    11'b01111100000: data <= 32'hbe99ac77;
    11'b01111100001: data <= 32'hbc42bb67;
    11'b01111100010: data <= 32'h380cbbff;
    11'b01111100011: data <= 32'h3a61bbb7;
    11'b01111100100: data <= 32'hb156be6f;
    11'b01111100101: data <= 32'hb8cbbffc;
    11'b01111100110: data <= 32'h23dab9ad;
    11'b01111100111: data <= 32'h34c73e00;
    11'b01111101000: data <= 32'hb87f4068;
    11'b01111101001: data <= 32'hbe193972;
    11'b01111101010: data <= 32'hbe06bb45;
    11'b01111101011: data <= 32'hbbe8b891;
    11'b01111101100: data <= 32'hba3b3a57;
    11'b01111101101: data <= 32'hb5e63c27;
    11'b01111101110: data <= 32'h3bdc2dd0;
    11'b01111101111: data <= 32'h409bb26d;
    11'b01111110000: data <= 32'h3f673ad3;
    11'b01111110001: data <= 32'had783eff;
    11'b01111110010: data <= 32'hbc8b3cd2;
    11'b01111110011: data <= 32'hafebaba5;
    11'b01111110100: data <= 32'h3cfaba6d;
    11'b01111110101: data <= 32'h3bcfbc94;
    11'b01111110110: data <= 32'hb40bbed6;
    11'b01111110111: data <= 32'hb542bfac;
    11'b01111111000: data <= 32'h3b47ba84;
    11'b01111111001: data <= 32'h3db63abc;
    11'b01111111010: data <= 32'h30303c73;
    11'b01111111011: data <= 32'hbe5eb42f;
    11'b01111111100: data <= 32'hc021bcf1;
    11'b01111111101: data <= 32'hbe19b6f6;
    11'b01111111110: data <= 32'hbc4d3a38;
    11'b01111111111: data <= 32'hb96e3787;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    