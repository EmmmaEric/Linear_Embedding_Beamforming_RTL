
module memory_rom_9(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbe063807;
    11'b00000000001: data <= 32'hba3134b5;
    11'b00000000010: data <= 32'h3bc8b40f;
    11'b00000000011: data <= 32'h3f5e35ab;
    11'b00000000100: data <= 32'h38a33e8e;
    11'b00000000101: data <= 32'hbd0f4002;
    11'b00000000110: data <= 32'hbd2c3ce8;
    11'b00000000111: data <= 32'h35c03729;
    11'b00000001000: data <= 32'h3d6c2c61;
    11'b00000001001: data <= 32'h398ab8fd;
    11'b00000001010: data <= 32'h1130be49;
    11'b00000001011: data <= 32'h3a14bdd0;
    11'b00000001100: data <= 32'h3fc82e91;
    11'b00000001101: data <= 32'h3ec03d38;
    11'b00000001110: data <= 32'h2e39380a;
    11'b00000001111: data <= 32'hbc7cbd0c;
    11'b00000010000: data <= 32'hbd17bea8;
    11'b00000010001: data <= 32'hbcb3b7eb;
    11'b00000010010: data <= 32'hbcd730e2;
    11'b00000010011: data <= 32'hb93aba16;
    11'b00000010100: data <= 32'h3854be49;
    11'b00000010101: data <= 32'h3b9fb819;
    11'b00000010110: data <= 32'hb37c3e2f;
    11'b00000010111: data <= 32'hbe4f40c7;
    11'b00000011000: data <= 32'hbd0b3e42;
    11'b00000011001: data <= 32'h30b8385f;
    11'b00000011010: data <= 32'h384e32d8;
    11'b00000011011: data <= 32'hb6adaaea;
    11'b00000011100: data <= 32'hb971b8b9;
    11'b00000011101: data <= 32'h3b77b838;
    11'b00000011110: data <= 32'h41713811;
    11'b00000011111: data <= 32'h40e83ce3;
    11'b00000100000: data <= 32'h3834373c;
    11'b00000100001: data <= 32'hba97baaa;
    11'b00000100010: data <= 32'hb9a1bb3a;
    11'b00000100011: data <= 32'hb445ab81;
    11'b00000100100: data <= 32'hb5cbb3ee;
    11'b00000100101: data <= 32'hb56dbf5c;
    11'b00000100110: data <= 32'h346ec159;
    11'b00000100111: data <= 32'h3889bc9f;
    11'b00000101000: data <= 32'hb3b93d06;
    11'b00000101001: data <= 32'hbcd54004;
    11'b00000101010: data <= 32'hbc433b38;
    11'b00000101011: data <= 32'hb60cacef;
    11'b00000101100: data <= 32'hb95c2f20;
    11'b00000101101: data <= 32'hbeba377d;
    11'b00000101110: data <= 32'hbd963054;
    11'b00000101111: data <= 32'h3a54b04f;
    11'b00000110000: data <= 32'h41623765;
    11'b00000110001: data <= 32'h40623cba;
    11'b00000110010: data <= 32'h32ff3bbd;
    11'b00000110011: data <= 32'hb98b34d2;
    11'b00000110100: data <= 32'h2a8134ee;
    11'b00000110101: data <= 32'h39df389b;
    11'b00000110110: data <= 32'h34d5b581;
    11'b00000110111: data <= 32'hb2dac079;
    11'b00000111000: data <= 32'h339ec1c8;
    11'b00000111001: data <= 32'h3b5cbcca;
    11'b00000111010: data <= 32'h39343b9b;
    11'b00000111011: data <= 32'hb34e3c9c;
    11'b00000111100: data <= 32'hb923b327;
    11'b00000111101: data <= 32'hb9fcbae7;
    11'b00000111110: data <= 32'hbddaa600;
    11'b00000111111: data <= 32'hc0ab3967;
    11'b00001000000: data <= 32'hbef62df4;
    11'b00001000001: data <= 32'h36a9b960;
    11'b00001000010: data <= 32'h3facb281;
    11'b00001000011: data <= 32'h3c9c3c11;
    11'b00001000100: data <= 32'hb8233e58;
    11'b00001000101: data <= 32'hb9b33d87;
    11'b00001000110: data <= 32'h384a3d03;
    11'b00001000111: data <= 32'h3c663c5c;
    11'b00001001000: data <= 32'h3176a77c;
    11'b00001001001: data <= 32'hb89fbedf;
    11'b00001001010: data <= 32'h3445c048;
    11'b00001001011: data <= 32'h3ebbb969;
    11'b00001001100: data <= 32'h3f783a3f;
    11'b00001001101: data <= 32'h3a933612;
    11'b00001001110: data <= 32'hb067bbef;
    11'b00001001111: data <= 32'hb910bc77;
    11'b00001010000: data <= 32'hbd432f72;
    11'b00001010001: data <= 32'hbfff38c9;
    11'b00001010010: data <= 32'hbe27b918;
    11'b00001010011: data <= 32'h28c5bf66;
    11'b00001010100: data <= 32'h3b80bcc1;
    11'b00001010101: data <= 32'h2e9f396d;
    11'b00001010110: data <= 32'hbc2f3f24;
    11'b00001010111: data <= 32'hb9763ea8;
    11'b00001011000: data <= 32'h38953d68;
    11'b00001011001: data <= 32'h38d63cd2;
    11'b00001011010: data <= 32'hba4c3815;
    11'b00001011011: data <= 32'hbd83b94c;
    11'b00001011100: data <= 32'h314cbc04;
    11'b00001011101: data <= 32'h4078ab10;
    11'b00001011110: data <= 32'h412439cd;
    11'b00001011111: data <= 32'h3d252eb8;
    11'b00001100000: data <= 32'h31fcbb0b;
    11'b00001100001: data <= 32'habd7b82a;
    11'b00001100010: data <= 32'hb57a3950;
    11'b00001100011: data <= 32'hbbc437ce;
    11'b00001100100: data <= 32'hbc14bdde;
    11'b00001100101: data <= 32'hb1bfc1c4;
    11'b00001100110: data <= 32'h35babf9e;
    11'b00001100111: data <= 32'hb2e534d6;
    11'b00001101000: data <= 32'hbae33d73;
    11'b00001101001: data <= 32'hb6463b8c;
    11'b00001101010: data <= 32'h357b38aa;
    11'b00001101011: data <= 32'hb5573b60;
    11'b00001101100: data <= 32'hbfe83bcd;
    11'b00001101101: data <= 32'hc0653368;
    11'b00001101110: data <= 32'haf7bb4ee;
    11'b00001101111: data <= 32'h403f2e7a;
    11'b00001110000: data <= 32'h408238ee;
    11'b00001110001: data <= 32'h3aff3546;
    11'b00001110010: data <= 32'h3191a7fe;
    11'b00001110011: data <= 32'h391b38db;
    11'b00001110100: data <= 32'h3a6f3db2;
    11'b00001110101: data <= 32'ha44a38a3;
    11'b00001110110: data <= 32'hb967befa;
    11'b00001110111: data <= 32'hb41dc219;
    11'b00001111000: data <= 32'h36eebf89;
    11'b00001111001: data <= 32'h360c2e1b;
    11'b00001111010: data <= 32'h25783861;
    11'b00001111011: data <= 32'h316cb4f6;
    11'b00001111100: data <= 32'h3264b797;
    11'b00001111101: data <= 32'hbbcd3878;
    11'b00001111110: data <= 32'hc12c3cc4;
    11'b00001111111: data <= 32'hc10c372c;
    11'b00010000000: data <= 32'hb71eb84b;
    11'b00010000001: data <= 32'h3d7ab71d;
    11'b00010000010: data <= 32'h3c673500;
    11'b00010000011: data <= 32'haf053988;
    11'b00010000100: data <= 32'hacaa3af2;
    11'b00010000101: data <= 32'h3c713e11;
    11'b00010000110: data <= 32'h3da33fe1;
    11'b00010000111: data <= 32'h315b3b3b;
    11'b00010001000: data <= 32'hbb26bce0;
    11'b00010001001: data <= 32'hb5abc066;
    11'b00010001010: data <= 32'h3b60bc93;
    11'b00010001011: data <= 32'h3d8c3081;
    11'b00010001100: data <= 32'h3c26b25a;
    11'b00010001101: data <= 32'h39ffbd33;
    11'b00010001110: data <= 32'h361bbc30;
    11'b00010001111: data <= 32'hba5a3837;
    11'b00010010000: data <= 32'hc0573ce0;
    11'b00010010001: data <= 32'hc04894c6;
    11'b00010010010: data <= 32'hb90ebdef;
    11'b00010010011: data <= 32'h36bfbd90;
    11'b00010010100: data <= 32'hb0f1b059;
    11'b00010010101: data <= 32'hbbae3a2b;
    11'b00010010110: data <= 32'hb3a33c5a;
    11'b00010010111: data <= 32'h3ce83e36;
    11'b00010011000: data <= 32'h3cc63fcf;
    11'b00010011001: data <= 32'hb8503d25;
    11'b00010011010: data <= 32'hbe92b233;
    11'b00010011011: data <= 32'hb8b1bafb;
    11'b00010011100: data <= 32'h3d3db282;
    11'b00010011101: data <= 32'h400034d0;
    11'b00010011110: data <= 32'h3dd7b83a;
    11'b00010011111: data <= 32'h3bf7bddb;
    11'b00010100000: data <= 32'h3abcb9c9;
    11'b00010100001: data <= 32'h31033c05;
    11'b00010100010: data <= 32'hbbc03cfe;
    11'b00010100011: data <= 32'hbd44b90e;
    11'b00010100100: data <= 32'hb8f6c0cd;
    11'b00010100101: data <= 32'hb221c029;
    11'b00010100110: data <= 32'hb9f7b7cc;
    11'b00010100111: data <= 32'hbc463681;
    11'b00010101000: data <= 32'ha98a3604;
    11'b00010101001: data <= 32'h3c8a3913;
    11'b00010101010: data <= 32'h37aa3d8b;
    11'b00010101011: data <= 32'hbe5b3e16;
    11'b00010101100: data <= 32'hc0e439b9;
    11'b00010101101: data <= 32'hbb262dc1;
    11'b00010101110: data <= 32'h3cd0344a;
    11'b00010101111: data <= 32'h3eb33514;
    11'b00010110000: data <= 32'h3b62b6f1;
    11'b00010110001: data <= 32'h39e4bae0;
    11'b00010110010: data <= 32'h3d4d33be;
    11'b00010110011: data <= 32'h3d3a3f05;
    11'b00010110100: data <= 32'h33cc3da0;
    11'b00010110101: data <= 32'hb91cbaef;
    11'b00010110110: data <= 32'hb851c115;
    11'b00010110111: data <= 32'hb363bfd8;
    11'b00010111000: data <= 32'hb698b7e5;
    11'b00010111001: data <= 32'hb600b301;
    11'b00010111010: data <= 32'h380ebb03;
    11'b00010111011: data <= 32'h3c5eb95a;
    11'b00010111100: data <= 32'hacda3973;
    11'b00010111101: data <= 32'hc0513e33;
    11'b00010111110: data <= 32'hc1693c1b;
    11'b00010111111: data <= 32'hbc493047;
    11'b00011000000: data <= 32'h38d5ab55;
    11'b00011000001: data <= 32'h382928fe;
    11'b00011000010: data <= 32'hb4aeb237;
    11'b00011000011: data <= 32'h30caad73;
    11'b00011000100: data <= 32'h3e5c3c61;
    11'b00011000101: data <= 32'h3ff34085;
    11'b00011000110: data <= 32'h39ac3e8a;
    11'b00011000111: data <= 32'hb8d3b74c;
    11'b00011001000: data <= 32'hb8b1bebf;
    11'b00011001001: data <= 32'h3000bc0a;
    11'b00011001010: data <= 32'h36ffafc8;
    11'b00011001011: data <= 32'h388ab9fe;
    11'b00011001100: data <= 32'h3c4abfb6;
    11'b00011001101: data <= 32'h3cedbe1f;
    11'b00011001110: data <= 32'h281835d0;
    11'b00011001111: data <= 32'hbef03dfc;
    11'b00011010000: data <= 32'hc04639af;
    11'b00011010001: data <= 32'hbba9b8fc;
    11'b00011010010: data <= 32'hb035bb41;
    11'b00011010011: data <= 32'hba4eb697;
    11'b00011010100: data <= 32'hbdbeafd7;
    11'b00011010101: data <= 32'hb549314c;
    11'b00011010110: data <= 32'h3e5f3c7f;
    11'b00011010111: data <= 32'h3f984030;
    11'b00011011000: data <= 32'h32fe3f02;
    11'b00011011001: data <= 32'hbce735e6;
    11'b00011011010: data <= 32'hba9ab502;
    11'b00011011011: data <= 32'h376c3329;
    11'b00011011100: data <= 32'h3c283600;
    11'b00011011101: data <= 32'h3bd6bb7f;
    11'b00011011110: data <= 32'h3cd6c06c;
    11'b00011011111: data <= 32'h3de6bdc8;
    11'b00011100000: data <= 32'h3a6c3974;
    11'b00011100001: data <= 32'hb7e73e19;
    11'b00011100010: data <= 32'hbc1a310d;
    11'b00011100011: data <= 32'hb8c4bdf8;
    11'b00011100100: data <= 32'hb8a1be51;
    11'b00011100101: data <= 32'hbdf8b989;
    11'b00011100110: data <= 32'hbf3bb528;
    11'b00011100111: data <= 32'hb54bb64e;
    11'b00011101000: data <= 32'h3df03192;
    11'b00011101001: data <= 32'h3d203d0a;
    11'b00011101010: data <= 32'hb9fd3e8b;
    11'b00011101011: data <= 32'hc0023c61;
    11'b00011101100: data <= 32'hbc603a0e;
    11'b00011101101: data <= 32'h37823bde;
    11'b00011101110: data <= 32'h3aac3905;
    11'b00011101111: data <= 32'h36b5ba6c;
    11'b00011110000: data <= 32'h39acbedf;
    11'b00011110001: data <= 32'h3e7cb8c4;
    11'b00011110010: data <= 32'h3f0b3d91;
    11'b00011110011: data <= 32'h3a8f3ead;
    11'b00011110100: data <= 32'ha902b080;
    11'b00011110101: data <= 32'hb39fbee1;
    11'b00011110110: data <= 32'hb869bdc8;
    11'b00011110111: data <= 32'hbd1eb7e4;
    11'b00011111000: data <= 32'hbd0fb91f;
    11'b00011111001: data <= 32'h30ffbdd5;
    11'b00011111010: data <= 32'h3dc5bce5;
    11'b00011111011: data <= 32'h39a3337a;
    11'b00011111100: data <= 32'hbd803d6a;
    11'b00011111101: data <= 32'hc0823d3e;
    11'b00011111110: data <= 32'hbc6d3b6f;
    11'b00011111111: data <= 32'h30763ac5;
    11'b00100000000: data <= 32'hb092371a;
    11'b00100000001: data <= 32'hbb0fb88f;
    11'b00100000010: data <= 32'hb25fbba8;
    11'b00100000011: data <= 32'h3e343494;
    11'b00100000100: data <= 32'h40a43f98;
    11'b00100000101: data <= 32'h3dac3f18;
    11'b00100000110: data <= 32'h33272977;
    11'b00100000111: data <= 32'hb0c8bc1c;
    11'b00100001000: data <= 32'hb24ab6af;
    11'b00100001001: data <= 32'hb799321c;
    11'b00100001010: data <= 32'hb532ba9b;
    11'b00100001011: data <= 32'h39d3c0be;
    11'b00100001100: data <= 32'h3dffc071;
    11'b00100001101: data <= 32'h3908b590;
    11'b00100001110: data <= 32'hbc643c79;
    11'b00100001111: data <= 32'hbe823bd7;
    11'b00100010000: data <= 32'hb99933bd;
    11'b00100010001: data <= 32'hb40f2882;
    11'b00100010010: data <= 32'hbd359fe3;
    11'b00100010011: data <= 32'hc054b734;
    11'b00100010100: data <= 32'hbbcbb88a;
    11'b00100010101: data <= 32'h3d50371f;
    11'b00100010110: data <= 32'h40643ec2;
    11'b00100010111: data <= 32'h3c123e83;
    11'b00100011000: data <= 32'hb524384f;
    11'b00100011001: data <= 32'hb5f53235;
    11'b00100011010: data <= 32'h314b3ba7;
    11'b00100011011: data <= 32'h332c3c08;
    11'b00100011100: data <= 32'h3265ba00;
    11'b00100011101: data <= 32'h3ac1c132;
    11'b00100011110: data <= 32'h3e12c07d;
    11'b00100011111: data <= 32'h3c5fb0ce;
    11'b00100100000: data <= 32'ha18c3c69;
    11'b00100100001: data <= 32'hb60736ac;
    11'b00100100010: data <= 32'h9533b97c;
    11'b00100100011: data <= 32'hb681b9d3;
    11'b00100100100: data <= 32'hbfbcb499;
    11'b00100100101: data <= 32'hc154b787;
    11'b00100100110: data <= 32'hbc90bad0;
    11'b00100100111: data <= 32'h3c90b5a0;
    11'b00100101000: data <= 32'h3e4a39d5;
    11'b00100101001: data <= 32'h26433caf;
    11'b00100101010: data <= 32'hbca83b96;
    11'b00100101011: data <= 32'hb9393cb6;
    11'b00100101100: data <= 32'h34ec3f74;
    11'b00100101101: data <= 32'h34223de5;
    11'b00100101110: data <= 32'hb2b6b7ef;
    11'b00100101111: data <= 32'h33a2c02f;
    11'b00100110000: data <= 32'h3d56bd98;
    11'b00100110001: data <= 32'h3ee638c3;
    11'b00100110010: data <= 32'h3cd13d0d;
    11'b00100110011: data <= 32'h3a30248c;
    11'b00100110100: data <= 32'h38edbc77;
    11'b00100110101: data <= 32'hb2ebb9ec;
    11'b00100110110: data <= 32'hbed0a033;
    11'b00100110111: data <= 32'hc050b7b9;
    11'b00100111000: data <= 32'hb93bbe5c;
    11'b00100111001: data <= 32'h3c6fbe91;
    11'b00100111010: data <= 32'h3b61b787;
    11'b00100111011: data <= 32'hba2d38b7;
    11'b00100111100: data <= 32'hbe393bab;
    11'b00100111101: data <= 32'hb8e63d4b;
    11'b00100111110: data <= 32'h34013f2e;
    11'b00100111111: data <= 32'hb6793d56;
    11'b00101000000: data <= 32'hbd95b41b;
    11'b00101000001: data <= 32'hbac2bd20;
    11'b00101000010: data <= 32'h3b7fb60d;
    11'b00101000011: data <= 32'h40153cf1;
    11'b00101000100: data <= 32'h3f113d5b;
    11'b00101000101: data <= 32'h3c8ea874;
    11'b00101000110: data <= 32'h3a67b9c4;
    11'b00101000111: data <= 32'h317f3151;
    11'b00101001000: data <= 32'hbae53abf;
    11'b00101001001: data <= 32'hbc70b53f;
    11'b00101001010: data <= 32'h2902c076;
    11'b00101001011: data <= 32'h3ca3c130;
    11'b00101001100: data <= 32'h392ebcbf;
    11'b00101001101: data <= 32'hba2b327a;
    11'b00101001110: data <= 32'hbc393878;
    11'b00101001111: data <= 32'haac138de;
    11'b00101010000: data <= 32'h32513b4f;
    11'b00101010001: data <= 32'hbd1c3a41;
    11'b00101010010: data <= 32'hc140b0bb;
    11'b00101010011: data <= 32'hbf21b9d2;
    11'b00101010100: data <= 32'h381528c4;
    11'b00101010101: data <= 32'h3f3b3ca9;
    11'b00101010110: data <= 32'h3d5f3c42;
    11'b00101010111: data <= 32'h38823031;
    11'b00101011000: data <= 32'h38143298;
    11'b00101011001: data <= 32'h38243def;
    11'b00101011010: data <= 32'ha80f3f60;
    11'b00101011011: data <= 32'hb59f9552;
    11'b00101011100: data <= 32'h34dfc09f;
    11'b00101011101: data <= 32'h3c51c131;
    11'b00101011110: data <= 32'h3a6abbfe;
    11'b00101011111: data <= 32'h24a932c8;
    11'b00101100000: data <= 32'h302d1b33;
    11'b00101100001: data <= 32'h3abfb6c8;
    11'b00101100010: data <= 32'h3553ab6b;
    11'b00101100011: data <= 32'hbee9358d;
    11'b00101100100: data <= 32'hc237ae8d;
    11'b00101100101: data <= 32'hc000b9d4;
    11'b00101100110: data <= 32'h34c1b767;
    11'b00101100111: data <= 32'h3cb0347c;
    11'b00101101000: data <= 32'h343e3683;
    11'b00101101001: data <= 32'hb7563335;
    11'b00101101010: data <= 32'h2ce13bda;
    11'b00101101011: data <= 32'h399240c1;
    11'b00101101100: data <= 32'h341340cf;
    11'b00101101101: data <= 32'hb77e354e;
    11'b00101101110: data <= 32'hb2a6bf14;
    11'b00101101111: data <= 32'h39a5beb9;
    11'b00101110000: data <= 32'h3c68aeda;
    11'b00101110001: data <= 32'h3c033819;
    11'b00101110010: data <= 32'h3d16b694;
    11'b00101110011: data <= 32'h3e65bc4e;
    11'b00101110100: data <= 32'h3942b5ad;
    11'b00101110101: data <= 32'hbdbb3819;
    11'b00101110110: data <= 32'hc1172b00;
    11'b00101110111: data <= 32'hbd9ebc89;
    11'b00101111000: data <= 32'h3622be04;
    11'b00101111001: data <= 32'h3823bb46;
    11'b00101111010: data <= 32'hb9cfb596;
    11'b00101111011: data <= 32'hbc802a35;
    11'b00101111100: data <= 32'ha4183c22;
    11'b00101111101: data <= 32'h3a3d408b;
    11'b00101111110: data <= 32'had6d4067;
    11'b00101111111: data <= 32'hbd9237c2;
    11'b00110000000: data <= 32'hbd18bba3;
    11'b00110000001: data <= 32'h2efab7cf;
    11'b00110000010: data <= 32'h3cbd3a5d;
    11'b00110000011: data <= 32'h3dc639e6;
    11'b00110000100: data <= 32'h3e79b89a;
    11'b00110000101: data <= 32'h3f15bbe9;
    11'b00110000110: data <= 32'h3c02347e;
    11'b00110000111: data <= 32'hb8a93d55;
    11'b00110001000: data <= 32'hbd6636b8;
    11'b00110001001: data <= 32'hb775be07;
    11'b00110001010: data <= 32'h38c0c09d;
    11'b00110001011: data <= 32'h3112be7e;
    11'b00110001100: data <= 32'hbc11ba38;
    11'b00110001101: data <= 32'hbb3ab5c5;
    11'b00110001110: data <= 32'h37ec34c4;
    11'b00110001111: data <= 32'h3b7d3d0f;
    11'b00110010000: data <= 32'hb9523db7;
    11'b00110010001: data <= 32'hc0e736ea;
    11'b00110010010: data <= 32'hc071b575;
    11'b00110010011: data <= 32'hb6923272;
    11'b00110010100: data <= 32'h3b183c0c;
    11'b00110010101: data <= 32'h3bd73846;
    11'b00110010110: data <= 32'h3b8bb8dc;
    11'b00110010111: data <= 32'h3d2fb5de;
    11'b00110011000: data <= 32'h3cca3da4;
    11'b00110011001: data <= 32'h34a040b4;
    11'b00110011010: data <= 32'hb55c3b11;
    11'b00110011011: data <= 32'h2e05bde0;
    11'b00110011100: data <= 32'h38e5c080;
    11'b00110011101: data <= 32'h303dbd73;
    11'b00110011110: data <= 32'hb84fb90c;
    11'b00110011111: data <= 32'h2cf8ba50;
    11'b00110100000: data <= 32'h3da6ba1f;
    11'b00110100001: data <= 32'h3cf92b50;
    11'b00110100010: data <= 32'hbb9f3993;
    11'b00110100011: data <= 32'hc1b635a4;
    11'b00110100100: data <= 32'hc0cab1f3;
    11'b00110100101: data <= 32'hb85023dc;
    11'b00110100110: data <= 32'h357635a3;
    11'b00110100111: data <= 32'hb00eb06e;
    11'b00110101000: data <= 32'hb4b0b9ad;
    11'b00110101001: data <= 32'h389332a2;
    11'b00110101010: data <= 32'h3ceb406b;
    11'b00110101011: data <= 32'h39a441cb;
    11'b00110101100: data <= 32'hb07c3cbf;
    11'b00110101101: data <= 32'hb178bbcb;
    11'b00110101110: data <= 32'h33adbd35;
    11'b00110101111: data <= 32'h332ab47d;
    11'b00110110000: data <= 32'h32ceab5e;
    11'b00110110001: data <= 32'h3c71bc30;
    11'b00110110010: data <= 32'h405abe18;
    11'b00110110011: data <= 32'h3e60b85e;
    11'b00110110100: data <= 32'hb94638be;
    11'b00110110101: data <= 32'hc08237b5;
    11'b00110110110: data <= 32'hbe8bb61c;
    11'b00110110111: data <= 32'hb2a7ba23;
    11'b00110111000: data <= 32'hb117b9b3;
    11'b00110111001: data <= 32'hbcd4bb69;
    11'b00110111010: data <= 32'hbd08bbbb;
    11'b00110111011: data <= 32'h321d32e6;
    11'b00110111100: data <= 32'h3d04401f;
    11'b00110111101: data <= 32'h38854120;
    11'b00110111110: data <= 32'hba4b3c88;
    11'b00110111111: data <= 32'hbc5db4ce;
    11'b00111000000: data <= 32'hb665a7f4;
    11'b00111000001: data <= 32'h31ca3b4b;
    11'b00111000010: data <= 32'h38843785;
    11'b00111000011: data <= 32'h3da4bc7f;
    11'b00111000100: data <= 32'h4084be7b;
    11'b00111000101: data <= 32'h3f1eb276;
    11'b00111000110: data <= 32'h2c923cf9;
    11'b00111000111: data <= 32'hbbe93b1c;
    11'b00111001000: data <= 32'hb6b6b8c1;
    11'b00111001001: data <= 32'h3500bdc4;
    11'b00111001010: data <= 32'hb682bd7e;
    11'b00111001011: data <= 32'hbeaabd38;
    11'b00111001100: data <= 32'hbd5bbd16;
    11'b00111001101: data <= 32'h3808b6e3;
    11'b00111001110: data <= 32'h3dc33bed;
    11'b00111001111: data <= 32'h314f3e21;
    11'b00111010000: data <= 32'hbebb3a2f;
    11'b00111010001: data <= 32'hbfe831eb;
    11'b00111010010: data <= 32'hbb423a82;
    11'b00111010011: data <= 32'hacad3dc4;
    11'b00111010100: data <= 32'h30f637e9;
    11'b00111010101: data <= 32'h396dbcab;
    11'b00111010110: data <= 32'h3e38bcc3;
    11'b00111010111: data <= 32'h3eba39e0;
    11'b00111011000: data <= 32'h3a724060;
    11'b00111011001: data <= 32'h31693d7a;
    11'b00111011010: data <= 32'h376eb85e;
    11'b00111011011: data <= 32'h38b5bd98;
    11'b00111011100: data <= 32'hb6b5bc40;
    11'b00111011101: data <= 32'hbd8abbbd;
    11'b00111011110: data <= 32'hb89ebdc1;
    11'b00111011111: data <= 32'h3d54bd6e;
    11'b00111100000: data <= 32'h3f25b590;
    11'b00111100001: data <= 32'habfb378b;
    11'b00111100010: data <= 32'hc0203680;
    11'b00111100011: data <= 32'hc03634c8;
    11'b00111100100: data <= 32'hbb1a3a98;
    11'b00111100101: data <= 32'hb6643c1c;
    11'b00111100110: data <= 32'hba9eac5d;
    11'b00111100111: data <= 32'hb969bd46;
    11'b00111101000: data <= 32'h380cb9b8;
    11'b00111101001: data <= 32'h3da03dea;
    11'b00111101010: data <= 32'h3c9d4164;
    11'b00111101011: data <= 32'h38773e48;
    11'b00111101100: data <= 32'h3791b30c;
    11'b00111101101: data <= 32'h35b4b871;
    11'b00111101110: data <= 32'hb609300e;
    11'b00111101111: data <= 32'hba1bad51;
    11'b00111110000: data <= 32'h35ecbd86;
    11'b00111110001: data <= 32'h4021c00d;
    11'b00111110010: data <= 32'h4028bc90;
    11'b00111110011: data <= 32'h2f3e2c4d;
    11'b00111110100: data <= 32'hbe2c35bc;
    11'b00111110101: data <= 32'hbd023087;
    11'b00111110110: data <= 32'hb44e324d;
    11'b00111110111: data <= 32'hb8b92d1a;
    11'b00111111000: data <= 32'hbf38ba99;
    11'b00111111001: data <= 32'hbf4dbe3a;
    11'b00111111010: data <= 32'hb254b91e;
    11'b00111111011: data <= 32'h3cdd3d8d;
    11'b00111111100: data <= 32'h3c214090;
    11'b00111111101: data <= 32'h2d673d0b;
    11'b00111111110: data <= 32'hb4bf3135;
    11'b00111111111: data <= 32'hb3c838e1;
    11'b01000000000: data <= 32'hb6f53dfe;
    11'b01000000001: data <= 32'hb64a3a46;
    11'b01000000010: data <= 32'h39a2bcd4;
    11'b01000000011: data <= 32'h402cc03c;
    11'b01000000100: data <= 32'h4019bbd9;
    11'b01000000101: data <= 32'h38a63841;
    11'b01000000110: data <= 32'hb61539a6;
    11'b01000000111: data <= 32'h3067a87d;
    11'b01000001000: data <= 32'h38cdb738;
    11'b01000001001: data <= 32'hb87bb8bb;
    11'b01000001010: data <= 32'hc07abca8;
    11'b01000001011: data <= 32'hc033bec9;
    11'b01000001100: data <= 32'haed4bc3d;
    11'b01000001101: data <= 32'h3d4236a3;
    11'b01000001110: data <= 32'h396a3c5b;
    11'b01000001111: data <= 32'hb9fb386a;
    11'b01000010000: data <= 32'hbcaa35a1;
    11'b01000010001: data <= 32'hb9d33da6;
    11'b01000010010: data <= 32'hb8964077;
    11'b01000010011: data <= 32'hb8f73c44;
    11'b01000010100: data <= 32'h2bedbc83;
    11'b01000010101: data <= 32'h3cf4beeb;
    11'b01000010110: data <= 32'h3e76b072;
    11'b01000010111: data <= 32'h3c0c3dbb;
    11'b01000011000: data <= 32'h39c93cb1;
    11'b01000011001: data <= 32'h3cf1ab38;
    11'b01000011010: data <= 32'h3cafb85b;
    11'b01000011011: data <= 32'hb699b5c3;
    11'b01000011100: data <= 32'hbff7b9a5;
    11'b01000011101: data <= 32'hbdd6be37;
    11'b01000011110: data <= 32'h392abebf;
    11'b01000011111: data <= 32'h3e94bae2;
    11'b01000100000: data <= 32'h36a8b22c;
    11'b01000100001: data <= 32'hbce1b090;
    11'b01000100010: data <= 32'hbd733447;
    11'b01000100011: data <= 32'hb8ec3dca;
    11'b01000100100: data <= 32'hb9073fdc;
    11'b01000100101: data <= 32'hbd4838ee;
    11'b01000100110: data <= 32'hbce5bd05;
    11'b01000100111: data <= 32'ha7d6bcfe;
    11'b01000101000: data <= 32'h3be73944;
    11'b01000101001: data <= 32'h3c803ff9;
    11'b01000101010: data <= 32'h3c803d3b;
    11'b01000101011: data <= 32'h3dab297b;
    11'b01000101100: data <= 32'h3c5f2982;
    11'b01000101101: data <= 32'hb53b3a11;
    11'b01000101110: data <= 32'hbd89363b;
    11'b01000101111: data <= 32'hb7ecbc88;
    11'b01000110000: data <= 32'h3dacc030;
    11'b01000110001: data <= 32'h3f95be9d;
    11'b01000110010: data <= 32'h3693ba5e;
    11'b01000110011: data <= 32'hbb66b647;
    11'b01000110100: data <= 32'hb8a328c5;
    11'b01000110101: data <= 32'h32573ac4;
    11'b01000110110: data <= 32'hb75a3c23;
    11'b01000110111: data <= 32'hc00bb12c;
    11'b01000111000: data <= 32'hc0babde4;
    11'b01000111001: data <= 32'hbba4bc26;
    11'b01000111010: data <= 32'h38613a14;
    11'b01000111011: data <= 32'h3b2a3e9c;
    11'b01000111100: data <= 32'h39743a9c;
    11'b01000111101: data <= 32'h399e2d43;
    11'b01000111110: data <= 32'h37fb3b6d;
    11'b01000111111: data <= 32'hb608403a;
    11'b01001000000: data <= 32'hbb573dfa;
    11'b01001000001: data <= 32'h0fc4b956;
    11'b01001000010: data <= 32'h3e10c014;
    11'b01001000011: data <= 32'h3ee6be19;
    11'b01001000100: data <= 32'h387eb6c5;
    11'b01001000101: data <= 32'ha89fad90;
    11'b01001000110: data <= 32'h3a50b0ae;
    11'b01001000111: data <= 32'h3d433061;
    11'b01001001000: data <= 32'haea53381;
    11'b01001001001: data <= 32'hc08cb8a4;
    11'b01001001010: data <= 32'hc156be04;
    11'b01001001011: data <= 32'hbbf1bcb2;
    11'b01001001100: data <= 32'h38782a7b;
    11'b01001001101: data <= 32'h382937c5;
    11'b01001001110: data <= 32'hb1deb045;
    11'b01001001111: data <= 32'hb433acf2;
    11'b01001010000: data <= 32'hac0d3e17;
    11'b01001010001: data <= 32'hb71341c1;
    11'b01001010010: data <= 32'hbb383fc4;
    11'b01001010011: data <= 32'hb647b739;
    11'b01001010100: data <= 32'h39a2be70;
    11'b01001010101: data <= 32'h3c32b959;
    11'b01001010110: data <= 32'h390d384c;
    11'b01001010111: data <= 32'h3ab83727;
    11'b01001011000: data <= 32'h3fabb2c8;
    11'b01001011001: data <= 32'h402cb10a;
    11'b01001011010: data <= 32'h335c3380;
    11'b01001011011: data <= 32'hbfd4b18a;
    11'b01001011100: data <= 32'hc00dbc8f;
    11'b01001011101: data <= 32'hb2f4bdc5;
    11'b01001011110: data <= 32'h3b7ebbdf;
    11'b01001011111: data <= 32'h337aba9e;
    11'b01001100000: data <= 32'hba8bbc3f;
    11'b01001100001: data <= 32'hb95bb658;
    11'b01001100010: data <= 32'ha4543dd7;
    11'b01001100011: data <= 32'hb4e9413e;
    11'b01001100100: data <= 32'hbd083e08;
    11'b01001100101: data <= 32'hbdb9b8c6;
    11'b01001100110: data <= 32'hb8bdbc70;
    11'b01001100111: data <= 32'h3135341e;
    11'b01001101000: data <= 32'h37773d24;
    11'b01001101001: data <= 32'h3c763948;
    11'b01001101010: data <= 32'h4041b448;
    11'b01001101011: data <= 32'h40252f23;
    11'b01001101100: data <= 32'h355b3c6a;
    11'b01001101101: data <= 32'hbd523b86;
    11'b01001101110: data <= 32'hbbafb72f;
    11'b01001101111: data <= 32'h39c2be25;
    11'b01001110000: data <= 32'h3d18be80;
    11'b01001110001: data <= 32'h2ee8bde4;
    11'b01001110010: data <= 32'hba7dbdb1;
    11'b01001110011: data <= 32'hb037b98a;
    11'b01001110100: data <= 32'h3a6a3aa4;
    11'b01001110101: data <= 32'h302d3e78;
    11'b01001110110: data <= 32'hbe7f38be;
    11'b01001110111: data <= 32'hc0cabb3b;
    11'b01001111000: data <= 32'hbe48ba77;
    11'b01001111001: data <= 32'hb70738f0;
    11'b01001111010: data <= 32'h2f8a3cbe;
    11'b01001111011: data <= 32'h3908321a;
    11'b01001111100: data <= 32'h3d74b7bd;
    11'b01001111101: data <= 32'h3d7f393a;
    11'b01001111110: data <= 32'h3273408a;
    11'b01001111111: data <= 32'hba654036;
    11'b01010000000: data <= 32'hb389331d;
    11'b01010000001: data <= 32'h3c37bd3c;
    11'b01010000010: data <= 32'h3c8bbdba;
    11'b01010000011: data <= 32'h2675bc4f;
    11'b01010000100: data <= 32'hb438bc3b;
    11'b01010000101: data <= 32'h3c25ba7e;
    11'b01010000110: data <= 32'h3ff02ccc;
    11'b01010000111: data <= 32'h39ce38ed;
    11'b01010001000: data <= 32'hbea1ab49;
    11'b01010001001: data <= 32'hc13abbf0;
    11'b01010001010: data <= 32'hbe71b9ec;
    11'b01010001011: data <= 32'hb6b533b4;
    11'b01010001100: data <= 32'hb334334c;
    11'b01010001101: data <= 32'hb461baa7;
    11'b01010001110: data <= 32'h3341bb40;
    11'b01010001111: data <= 32'h38bc3bee;
    11'b01010010000: data <= 32'h2b7b41db;
    11'b01010010001: data <= 32'hb8e4412a;
    11'b01010010010: data <= 32'hb4f237ba;
    11'b01010010011: data <= 32'h3763baf3;
    11'b01010010100: data <= 32'h3684b84d;
    11'b01010010101: data <= 32'hb1c42691;
    11'b01010010110: data <= 32'h353db531;
    11'b01010010111: data <= 32'h4018ba49;
    11'b01010011000: data <= 32'h419eb5c1;
    11'b01010011001: data <= 32'h3ca33505;
    11'b01010011010: data <= 32'hbd222fa0;
    11'b01010011011: data <= 32'hbfb7b8c2;
    11'b01010011100: data <= 32'hb9c8b9de;
    11'b01010011101: data <= 32'h301fb7d1;
    11'b01010011110: data <= 32'hb6b1bba3;
    11'b01010011111: data <= 32'hbc15bf57;
    11'b01010100000: data <= 32'hb765bd82;
    11'b01010100001: data <= 32'h365b3a9a;
    11'b01010100010: data <= 32'h3263413e;
    11'b01010100011: data <= 32'hb9a24022;
    11'b01010100100: data <= 32'hbc1e3293;
    11'b01010100101: data <= 32'hb986b73e;
    11'b01010100110: data <= 32'hb88f37b4;
    11'b01010100111: data <= 32'hb8593c24;
    11'b01010101000: data <= 32'h374a3057;
    11'b01010101001: data <= 32'h4065ba8c;
    11'b01010101010: data <= 32'h417eb54d;
    11'b01010101011: data <= 32'h3cb63ae2;
    11'b01010101100: data <= 32'hb9c03c4a;
    11'b01010101101: data <= 32'hba423225;
    11'b01010101110: data <= 32'h3744b8bb;
    11'b01010101111: data <= 32'h39b6bb87;
    11'b01010110000: data <= 32'hb7eebe24;
    11'b01010110001: data <= 32'hbcebc061;
    11'b01010110010: data <= 32'hb3e2be90;
    11'b01010110011: data <= 32'h3c26334f;
    11'b01010110100: data <= 32'h39ce3e2e;
    11'b01010110101: data <= 32'hba7e3b7b;
    11'b01010110110: data <= 32'hbf15b57c;
    11'b01010110111: data <= 32'hbe64b2fd;
    11'b01010111000: data <= 32'hbcd13c21;
    11'b01010111001: data <= 32'hbb5c3d03;
    11'b01010111010: data <= 32'ha861b056;
    11'b01010111011: data <= 32'h3d7abc6c;
    11'b01010111100: data <= 32'h3f73ab51;
    11'b01010111101: data <= 32'h3a8f3f1a;
    11'b01010111110: data <= 32'hb4454050;
    11'b01010111111: data <= 32'h2f333b6f;
    11'b01011000000: data <= 32'h3c69b471;
    11'b01011000001: data <= 32'h3a5ab9a3;
    11'b01011000010: data <= 32'hb904bc53;
    11'b01011000011: data <= 32'hbb96beb4;
    11'b01011000100: data <= 32'h3938be42;
    11'b01011000101: data <= 32'h4041b721;
    11'b01011000110: data <= 32'h3da53649;
    11'b01011000111: data <= 32'hb9a5a632;
    11'b01011001000: data <= 32'hbf9fb959;
    11'b01011001001: data <= 32'hbe56b01b;
    11'b01011001010: data <= 32'hbc513b50;
    11'b01011001011: data <= 32'hbc7038a5;
    11'b01011001100: data <= 32'hbaebbc36;
    11'b01011001101: data <= 32'h2e5ebe88;
    11'b01011001110: data <= 32'h3a3f2e61;
    11'b01011001111: data <= 32'h36c440a0;
    11'b01011010000: data <= 32'had6d412a;
    11'b01011010001: data <= 32'h34953c86;
    11'b01011010010: data <= 32'h3a7b2be3;
    11'b01011010011: data <= 32'h32133065;
    11'b01011010100: data <= 32'hbb883076;
    11'b01011010101: data <= 32'hb88fb94a;
    11'b01011010110: data <= 32'h3e0bbd1c;
    11'b01011010111: data <= 32'h41d0baca;
    11'b01011011000: data <= 32'h3f53b094;
    11'b01011011001: data <= 32'hb608b131;
    11'b01011011010: data <= 32'hbcfab6c2;
    11'b01011011011: data <= 32'hb8bba4dc;
    11'b01011011100: data <= 32'hb47136ba;
    11'b01011011101: data <= 32'hbc32b6c5;
    11'b01011011110: data <= 32'hbe3fc007;
    11'b01011011111: data <= 32'hba76c044;
    11'b01011100000: data <= 32'h3429acf0;
    11'b01011100001: data <= 32'h361e4002;
    11'b01011100010: data <= 32'hadeb3fea;
    11'b01011100011: data <= 32'hb1e33914;
    11'b01011100100: data <= 32'hb06133d2;
    11'b01011100101: data <= 32'hb9f23c65;
    11'b01011100110: data <= 32'hbd7c3d69;
    11'b01011100111: data <= 32'hb80a3039;
    11'b01011101000: data <= 32'h3e86bc65;
    11'b01011101001: data <= 32'h418bbb0c;
    11'b01011101010: data <= 32'h3eb130bb;
    11'b01011101011: data <= 32'ha30d3878;
    11'b01011101100: data <= 32'hb0eb34f6;
    11'b01011101101: data <= 32'h3a3532f8;
    11'b01011101110: data <= 32'h39222d12;
    11'b01011101111: data <= 32'hbb1fbb94;
    11'b01011110000: data <= 32'hbf38c0a1;
    11'b01011110001: data <= 32'hbac8c08a;
    11'b01011110010: data <= 32'h3922b81a;
    11'b01011110011: data <= 32'h3aaa3bc9;
    11'b01011110100: data <= 32'hadce3959;
    11'b01011110101: data <= 32'hba31b3b4;
    11'b01011110110: data <= 32'hbbaf3346;
    11'b01011110111: data <= 32'hbd5e3ea6;
    11'b01011111000: data <= 32'hbeb23f4c;
    11'b01011111001: data <= 32'hbb0b309d;
    11'b01011111010: data <= 32'h3ab3bd22;
    11'b01011111011: data <= 32'h3ee7b9bc;
    11'b01011111100: data <= 32'h3c033b0a;
    11'b01011111101: data <= 32'h31ce3e23;
    11'b01011111110: data <= 32'h39e63c19;
    11'b01011111111: data <= 32'h3eb53814;
    11'b01100000000: data <= 32'h3c1d340d;
    11'b01100000001: data <= 32'hbb19b81d;
    11'b01100000010: data <= 32'hbe80bea6;
    11'b01100000011: data <= 32'hb0f3bfa4;
    11'b01100000100: data <= 32'h3e61bb7d;
    11'b01100000101: data <= 32'h3e01b142;
    11'b01100000110: data <= 32'h28f7b855;
    11'b01100000111: data <= 32'hbb5abb2d;
    11'b01100001000: data <= 32'hbb9d30d3;
    11'b01100001001: data <= 32'hbc6e3e88;
    11'b01100001010: data <= 32'hbe7b3d80;
    11'b01100001011: data <= 32'hbdeab8dc;
    11'b01100001100: data <= 32'hb694bf28;
    11'b01100001101: data <= 32'h3661b8f0;
    11'b01100001110: data <= 32'h34223d87;
    11'b01100001111: data <= 32'h314f3fca;
    11'b01100010000: data <= 32'h3bdf3c95;
    11'b01100010001: data <= 32'h3e7f393e;
    11'b01100010010: data <= 32'h38f93b26;
    11'b01100010011: data <= 32'hbcac3977;
    11'b01100010100: data <= 32'hbd4fb69f;
    11'b01100010101: data <= 32'h3907bd12;
    11'b01100010110: data <= 32'h40b0bc76;
    11'b01100010111: data <= 32'h3f78ba0f;
    11'b01100011000: data <= 32'h3343bb7c;
    11'b01100011001: data <= 32'hb6bdbb10;
    11'b01100011010: data <= 32'h24f33294;
    11'b01100011011: data <= 32'hadc33cef;
    11'b01100011100: data <= 32'hbcd737b2;
    11'b01100011101: data <= 32'hbfbfbe16;
    11'b01100011110: data <= 32'hbd71c085;
    11'b01100011111: data <= 32'hb643b9a5;
    11'b01100100000: data <= 32'haac33cc6;
    11'b01100100001: data <= 32'h2cbb3d70;
    11'b01100100010: data <= 32'h38ea3757;
    11'b01100100011: data <= 32'h3a8d3813;
    11'b01100100100: data <= 32'hb3d13e74;
    11'b01100100101: data <= 32'hbe593fb5;
    11'b01100100110: data <= 32'hbce33943;
    11'b01100100111: data <= 32'h3aa3ba40;
    11'b01100101000: data <= 32'h4072bc1d;
    11'b01100101001: data <= 32'h3e31b886;
    11'b01100101010: data <= 32'h34b1b631;
    11'b01100101011: data <= 32'h36feb3de;
    11'b01100101100: data <= 32'h3da43707;
    11'b01100101101: data <= 32'h3c713b24;
    11'b01100101110: data <= 32'hb9bbad80;
    11'b01100101111: data <= 32'hc00dbf57;
    11'b01100110000: data <= 32'hbdf9c08a;
    11'b01100110001: data <= 32'hb2cebb13;
    11'b01100110010: data <= 32'h3443360a;
    11'b01100110011: data <= 32'h2c6827ab;
    11'b01100110100: data <= 32'h2b93b993;
    11'b01100110101: data <= 32'ha1513076;
    11'b01100110110: data <= 32'hbad23ffb;
    11'b01100110111: data <= 32'hbf3340f8;
    11'b01100111000: data <= 32'hbd8c3b34;
    11'b01100111001: data <= 32'h334dba57;
    11'b01100111010: data <= 32'h3ca7baba;
    11'b01100111011: data <= 32'h38df2ee5;
    11'b01100111100: data <= 32'h301f3873;
    11'b01100111101: data <= 32'h3c843789;
    11'b01100111110: data <= 32'h40c9396a;
    11'b01100111111: data <= 32'h3f053b41;
    11'b01101000000: data <= 32'hb7f431cc;
    11'b01101000001: data <= 32'hbf32bcb5;
    11'b01101000010: data <= 32'hbafebea4;
    11'b01101000011: data <= 32'h3962bba1;
    11'b01101000100: data <= 32'h3b5eb866;
    11'b01101000101: data <= 32'h317abd08;
    11'b01101000110: data <= 32'hb248be89;
    11'b01101000111: data <= 32'hb06fb243;
    11'b01101001000: data <= 32'hb8fc3f8f;
    11'b01101001001: data <= 32'hbe1c403c;
    11'b01101001010: data <= 32'hbe9a340a;
    11'b01101001011: data <= 32'hba76bd0c;
    11'b01101001100: data <= 32'hb3a7b9d8;
    11'b01101001101: data <= 32'hb6fe396a;
    11'b01101001110: data <= 32'hb1e23c4d;
    11'b01101001111: data <= 32'h3d1638dd;
    11'b01101010000: data <= 32'h40dc3926;
    11'b01101010001: data <= 32'h3df43cf9;
    11'b01101010010: data <= 32'hb9ad3cae;
    11'b01101010011: data <= 32'hbdfa3077;
    11'b01101010100: data <= 32'hab93b9a6;
    11'b01101010101: data <= 32'h3dfeba6f;
    11'b01101010110: data <= 32'h3d3ebc0e;
    11'b01101010111: data <= 32'h3316bf02;
    11'b01101011000: data <= 32'h28c3bf34;
    11'b01101011001: data <= 32'h3913b3ee;
    11'b01101011010: data <= 32'h37363dea;
    11'b01101011011: data <= 32'hba793ce2;
    11'b01101011100: data <= 32'hbf09b9aa;
    11'b01101011101: data <= 32'hbe6cbf08;
    11'b01101011110: data <= 32'hbc8cb9bf;
    11'b01101011111: data <= 32'hbbc639ad;
    11'b01101100000: data <= 32'hb6d9395d;
    11'b01101100001: data <= 32'h3b08afcc;
    11'b01101100010: data <= 32'h3e983290;
    11'b01101100011: data <= 32'h38de3e6f;
    11'b01101100100: data <= 32'hbc9a407e;
    11'b01101100101: data <= 32'hbd473d4c;
    11'b01101100110: data <= 32'h352c2976;
    11'b01101100111: data <= 32'h3e2db822;
    11'b01101101000: data <= 32'h3bb9ba3e;
    11'b01101101001: data <= 32'h2569bd01;
    11'b01101101010: data <= 32'h3867bcc1;
    11'b01101101011: data <= 32'h3f679c19;
    11'b01101101100: data <= 32'h3f113c62;
    11'b01101101101: data <= 32'ha57a3816;
    11'b01101101110: data <= 32'hbe68bcb1;
    11'b01101101111: data <= 32'hbeb4bf0b;
    11'b01101110000: data <= 32'hbc1db94f;
    11'b01101110001: data <= 32'hb9c63310;
    11'b01101110010: data <= 32'hb729b7b5;
    11'b01101110011: data <= 32'h34c3bd8f;
    11'b01101110100: data <= 32'h39b1b7ab;
    11'b01101110101: data <= 32'hb05d3ed4;
    11'b01101110110: data <= 32'hbd824170;
    11'b01101110111: data <= 32'hbd283ea1;
    11'b01101111000: data <= 32'h262630cf;
    11'b01101111001: data <= 32'h394ab474;
    11'b01101111010: data <= 32'had1ead99;
    11'b01101111011: data <= 32'hb778b380;
    11'b01101111100: data <= 32'h3b75b5b3;
    11'b01101111101: data <= 32'h41763439;
    11'b01101111110: data <= 32'h410a3ba2;
    11'b01101111111: data <= 32'h35de3807;
    11'b01110000000: data <= 32'hbd1eb98d;
    11'b01110000001: data <= 32'hbc21bc3d;
    11'b01110000010: data <= 32'hae8bb696;
    11'b01110000011: data <= 32'h24c8b61c;
    11'b01110000100: data <= 32'hb4eabea1;
    11'b01110000101: data <= 32'hace1c0e9;
    11'b01110000110: data <= 32'h3571bc1f;
    11'b01110000111: data <= 32'had813dd8;
    11'b01110001000: data <= 32'hbc2640a4;
    11'b01110001001: data <= 32'hbcfc3bfe;
    11'b01110001010: data <= 32'hb972b5e2;
    11'b01110001011: data <= 32'hb8f3b26c;
    11'b01110001100: data <= 32'hbd13388f;
    11'b01110001101: data <= 32'hbc2737ef;
    11'b01110001110: data <= 32'h3b24a94c;
    11'b01110001111: data <= 32'h4175321e;
    11'b01110010000: data <= 32'h408c3c0a;
    11'b01110010001: data <= 32'h30be3ca8;
    11'b01110010010: data <= 32'hbbee37dc;
    11'b01110010011: data <= 32'hb0ce29ba;
    11'b01110010100: data <= 32'h3b382829;
    11'b01110010101: data <= 32'h38a4b8fd;
    11'b01110010110: data <= 32'hb44dc034;
    11'b01110010111: data <= 32'hada5c15a;
    11'b01110011000: data <= 32'h3a5dbc81;
    11'b01110011001: data <= 32'h3ac43c2a;
    11'b01110011010: data <= 32'hb17a3d79;
    11'b01110011011: data <= 32'hbc26af1b;
    11'b01110011100: data <= 32'hbce5bc1a;
    11'b01110011101: data <= 32'hbdd8b261;
    11'b01110011110: data <= 32'hbf933a80;
    11'b01110011111: data <= 32'hbd863646;
    11'b01110100000: data <= 32'h374cb8f1;
    11'b01110100001: data <= 32'h3f98b617;
    11'b01110100010: data <= 32'h3d1a3c33;
    11'b01110100011: data <= 32'hb6fc3fd7;
    11'b01110100100: data <= 32'hbabe3e73;
    11'b01110100101: data <= 32'h368e3b56;
    11'b01110100110: data <= 32'h3ced379a;
    11'b01110100111: data <= 32'h3663b4ef;
    11'b01110101000: data <= 32'hb8a4be3c;
    11'b01110101001: data <= 32'h2eaebfec;
    11'b01110101010: data <= 32'h3edeba1f;
    11'b01110101011: data <= 32'h402d3984;
    11'b01110101100: data <= 32'h3a203811;
    11'b01110101101: data <= 32'hb960babd;
    11'b01110101110: data <= 32'hbcaebccf;
    11'b01110101111: data <= 32'hbd43abbd;
    11'b01110110000: data <= 32'hbe693906;
    11'b01110110001: data <= 32'hbd49b755;
    11'b01110110010: data <= 32'hae32bf37;
    11'b01110110011: data <= 32'h3ab0bceb;
    11'b01110110100: data <= 32'h348a3b2b;
    11'b01110110101: data <= 32'hbac7408b;
    11'b01110110110: data <= 32'hba0f3fa5;
    11'b01110110111: data <= 32'h364f3c1d;
    11'b01110111000: data <= 32'h39393979;
    11'b01110111001: data <= 32'hb86c35f1;
    11'b01110111010: data <= 32'hbcf4b701;
    11'b01110111011: data <= 32'h3283bb67;
    11'b01110111100: data <= 32'h40ceb4ef;
    11'b01110111101: data <= 32'h419f382b;
    11'b01110111110: data <= 32'h3ccf33b9;
    11'b01110111111: data <= 32'hb528b957;
    11'b01111000000: data <= 32'hb81fb8e3;
    11'b01111000001: data <= 32'hb4d535ba;
    11'b01111000010: data <= 32'hb959353f;
    11'b01111000011: data <= 32'hbbfdbda9;
    11'b01111000100: data <= 32'hb792c1ae;
    11'b01111000101: data <= 32'h335cbf7d;
    11'b01111000110: data <= 32'h278e3887;
    11'b01111000111: data <= 32'hb91a3f52;
    11'b01111001000: data <= 32'hb87f3cb8;
    11'b01111001001: data <= 32'h159835a9;
    11'b01111001010: data <= 32'hb63b38c9;
    11'b01111001011: data <= 32'hbedb3c11;
    11'b01111001100: data <= 32'hbfc23803;
    11'b01111001101: data <= 32'h2686b4f1;
    11'b01111001110: data <= 32'h40a7b343;
    11'b01111001111: data <= 32'h41033734;
    11'b01111010000: data <= 32'h3af738b7;
    11'b01111010001: data <= 32'hb14f3433;
    11'b01111010010: data <= 32'h35a13765;
    11'b01111010011: data <= 32'h3b1c3bb0;
    11'b01111010100: data <= 32'h31f2345d;
    11'b01111010101: data <= 32'hba47bf08;
    11'b01111010110: data <= 32'hb8a9c209;
    11'b01111010111: data <= 32'h361bbf9b;
    11'b01111011000: data <= 32'h39843390;
    11'b01111011001: data <= 32'h31ec3b17;
    11'b01111011010: data <= 32'hb19dae25;
    11'b01111011011: data <= 32'hb505b8a9;
    11'b01111011100: data <= 32'hbc6a3691;
    11'b01111011101: data <= 32'hc0a13d4f;
    11'b01111011110: data <= 32'hc0883980;
    11'b01111011111: data <= 32'hb5e3b8cc;
    11'b01111100000: data <= 32'h3df8b9e1;
    11'b01111100001: data <= 32'h3d7134eb;
    11'b01111100010: data <= 32'h26ff3c82;
    11'b01111100011: data <= 32'hb2ba3cec;
    11'b01111100100: data <= 32'h3ba83d4d;
    11'b01111100101: data <= 32'h3df93dc5;
    11'b01111100110: data <= 32'h34d638c8;
    11'b01111100111: data <= 32'hbc06bcc8;
    11'b01111101000: data <= 32'hb883c065;
    11'b01111101001: data <= 32'h3c18bd3e;
    11'b01111101010: data <= 32'h3f072c91;
    11'b01111101011: data <= 32'h3c7e9a40;
    11'b01111101100: data <= 32'h3476bc5b;
    11'b01111101101: data <= 32'hb247bc45;
    11'b01111101110: data <= 32'hbb5c36ed;
    11'b01111101111: data <= 32'hbfb23d33;
    11'b01111110000: data <= 32'hc009300e;
    11'b01111110001: data <= 32'hba05be5a;
    11'b01111110010: data <= 32'h3690be59;
    11'b01111110011: data <= 32'h2fb2267c;
    11'b01111110100: data <= 32'hb9973d4a;
    11'b01111110101: data <= 32'hb4483de4;
    11'b01111110110: data <= 32'h3c503d78;
    11'b01111110111: data <= 32'h3cd53e0d;
    11'b01111111000: data <= 32'hb6e43c8e;
    11'b01111111001: data <= 32'hbea5ab91;
    11'b01111111010: data <= 32'hb8f6bb48;
    11'b01111111011: data <= 32'h3e34b84b;
    11'b01111111100: data <= 32'h40ce2c70;
    11'b01111111101: data <= 32'h3e13b62b;
    11'b01111111110: data <= 32'h385ebcd8;
    11'b01111111111: data <= 32'h35c7b9be;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    