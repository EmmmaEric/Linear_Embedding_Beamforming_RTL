
module memory_rom_60(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hb9c8bd9a;
    11'b00000000001: data <= 32'hb806ba78;
    11'b00000000010: data <= 32'h36333a35;
    11'b00000000011: data <= 32'h2cff3f78;
    11'b00000000100: data <= 32'hbd923c07;
    11'b00000000101: data <= 32'hc068ba37;
    11'b00000000110: data <= 32'hbe21bc7a;
    11'b00000000111: data <= 32'hb71834d5;
    11'b00000001000: data <= 32'h30913d5b;
    11'b00000001001: data <= 32'h396b3958;
    11'b00000001010: data <= 32'h3df7b43d;
    11'b00000001011: data <= 32'h3e7b35e6;
    11'b00000001100: data <= 32'h361c3f64;
    11'b00000001101: data <= 32'hbb793fe7;
    11'b00000001110: data <= 32'hb8ad3588;
    11'b00000001111: data <= 32'h3b79bd04;
    11'b00000010000: data <= 32'h3dcdbe47;
    11'b00000010001: data <= 32'h3617bd0d;
    11'b00000010010: data <= 32'hb614bcac;
    11'b00000010011: data <= 32'h381dbab7;
    11'b00000010100: data <= 32'h3e7c312b;
    11'b00000010101: data <= 32'h3aa43ac5;
    11'b00000010110: data <= 32'hbd9430e1;
    11'b00000010111: data <= 32'hc141bc3e;
    11'b00000011000: data <= 32'hbf82bc21;
    11'b00000011001: data <= 32'hb8ae30ed;
    11'b00000011010: data <= 32'haf9e38d4;
    11'b00000011011: data <= 32'ha977b54a;
    11'b00000011100: data <= 32'h369fba8f;
    11'b00000011101: data <= 32'h399e3924;
    11'b00000011110: data <= 32'h2c604154;
    11'b00000011111: data <= 32'hb9e0417a;
    11'b00000100000: data <= 32'hb6d53a3a;
    11'b00000100001: data <= 32'h38dbbb2f;
    11'b00000100010: data <= 32'h3a6dbb3e;
    11'b00000100011: data <= 32'h2bc1b4c8;
    11'b00000100100: data <= 32'h2e6db5e6;
    11'b00000100101: data <= 32'h3e70b955;
    11'b00000100110: data <= 32'h4160b445;
    11'b00000100111: data <= 32'h3dbb3550;
    11'b00000101000: data <= 32'hbc6c2aa8;
    11'b00000101001: data <= 32'hc06cba3a;
    11'b00000101010: data <= 32'hbccebb56;
    11'b00000101011: data <= 32'ha813b69c;
    11'b00000101100: data <= 32'hb1a2b89c;
    11'b00000101101: data <= 32'hb9fcbe0b;
    11'b00000101110: data <= 32'hb71ebdc9;
    11'b00000101111: data <= 32'h33e03864;
    11'b00000110000: data <= 32'h2d844148;
    11'b00000110001: data <= 32'hb9b940fb;
    11'b00000110010: data <= 32'hbb7c385d;
    11'b00000110011: data <= 32'hb756b8f7;
    11'b00000110100: data <= 32'hb47f2412;
    11'b00000110101: data <= 32'hb7193a83;
    11'b00000110110: data <= 32'h34633518;
    11'b00000110111: data <= 32'h400db8a1;
    11'b00000111000: data <= 32'h41d4b5b6;
    11'b00000111001: data <= 32'h3e1e3903;
    11'b00000111010: data <= 32'hb9823ac9;
    11'b00000111011: data <= 32'hbcec2b69;
    11'b00000111100: data <= 32'h9de5b923;
    11'b00000111101: data <= 32'h39d8baf7;
    11'b00000111110: data <= 32'hb058bd83;
    11'b00000111111: data <= 32'hbc46c048;
    11'b00001000000: data <= 32'hb80abf36;
    11'b00001000001: data <= 32'h396c2f01;
    11'b00001000010: data <= 32'h38f93f2d;
    11'b00001000011: data <= 32'hb9743db8;
    11'b00001000100: data <= 32'hbe82afe4;
    11'b00001000101: data <= 32'hbe15b80d;
    11'b00001000110: data <= 32'hbc9f3932;
    11'b00001000111: data <= 32'hbb473d36;
    11'b00001001000: data <= 32'haa99348b;
    11'b00001001001: data <= 32'h3de5bacf;
    11'b00001001010: data <= 32'h405bb3df;
    11'b00001001011: data <= 32'h3c6a3db0;
    11'b00001001100: data <= 32'hb5db4006;
    11'b00001001101: data <= 32'hb4e13bed;
    11'b00001001110: data <= 32'h3afdb3d0;
    11'b00001001111: data <= 32'h3c33ba5d;
    11'b00001010000: data <= 32'hb39bbce6;
    11'b00001010001: data <= 32'hbbcbbf4f;
    11'b00001010010: data <= 32'h326dbec9;
    11'b00001010011: data <= 32'h3f0eb6ae;
    11'b00001010100: data <= 32'h3dd63970;
    11'b00001010101: data <= 32'hb7c534e8;
    11'b00001010110: data <= 32'hbf9ab951;
    11'b00001010111: data <= 32'hbf3ab745;
    11'b00001011000: data <= 32'hbd0439d7;
    11'b00001011001: data <= 32'hbc583b11;
    11'b00001011010: data <= 32'hb9a8b868;
    11'b00001011011: data <= 32'h350ebdf8;
    11'b00001011100: data <= 32'h3c0cb26e;
    11'b00001011101: data <= 32'h383e401a;
    11'b00001011110: data <= 32'hb346416b;
    11'b00001011111: data <= 32'h2bb53dad;
    11'b00001100000: data <= 32'h3aee2d70;
    11'b00001100001: data <= 32'h38b0b132;
    11'b00001100010: data <= 32'hb917b20a;
    11'b00001100011: data <= 32'hb9efba73;
    11'b00001100100: data <= 32'h3c4fbd15;
    11'b00001100101: data <= 32'h4184ba21;
    11'b00001100110: data <= 32'h4030a521;
    11'b00001100111: data <= 32'hb147af64;
    11'b00001101000: data <= 32'hbde7b8b5;
    11'b00001101001: data <= 32'hbc42b473;
    11'b00001101010: data <= 32'hb81c36b7;
    11'b00001101011: data <= 32'hbb4daaf3;
    11'b00001101100: data <= 32'hbd4bbe9c;
    11'b00001101101: data <= 32'hb9a8c05e;
    11'b00001101110: data <= 32'h3389b619;
    11'b00001101111: data <= 32'h350f3fec;
    11'b00001110000: data <= 32'hb18840cc;
    11'b00001110001: data <= 32'hb2203c27;
    11'b00001110010: data <= 32'h2c213158;
    11'b00001110011: data <= 32'hb68b3964;
    11'b00001110100: data <= 32'hbce93c48;
    11'b00001110101: data <= 32'hb99f323c;
    11'b00001110110: data <= 32'h3da6bb71;
    11'b00001110111: data <= 32'h41dcbae4;
    11'b00001111000: data <= 32'h402b2652;
    11'b00001111001: data <= 32'h2e763659;
    11'b00001111010: data <= 32'hb8883077;
    11'b00001111011: data <= 32'h34362e44;
    11'b00001111100: data <= 32'h3868306c;
    11'b00001111101: data <= 32'hb8dbb9ed;
    11'b00001111110: data <= 32'hbe7dc07a;
    11'b00001111111: data <= 32'hbc05c0f6;
    11'b00010000000: data <= 32'h35d9b9c2;
    11'b00010000001: data <= 32'h39be3cbc;
    11'b00010000010: data <= 32'ha8e43cde;
    11'b00010000011: data <= 32'hb9662d79;
    11'b00010000100: data <= 32'hbacf22f6;
    11'b00010000101: data <= 32'hbcfa3d0f;
    11'b00010000110: data <= 32'hbebc3f23;
    11'b00010000111: data <= 32'hbbdd37a0;
    11'b00010001000: data <= 32'h3b18bc28;
    11'b00010001001: data <= 32'h402cbab5;
    11'b00010001010: data <= 32'h3d9c38bd;
    11'b00010001011: data <= 32'h31453d89;
    11'b00010001100: data <= 32'h34de3c23;
    11'b00010001101: data <= 32'h3d6d383c;
    11'b00010001110: data <= 32'h3ccb332e;
    11'b00010001111: data <= 32'hb81eb8b5;
    11'b00010010000: data <= 32'hbe62bf57;
    11'b00010010001: data <= 32'hb84cc04f;
    11'b00010010010: data <= 32'h3cfebc09;
    11'b00010010011: data <= 32'h3e0a301e;
    11'b00010010100: data <= 32'h3331af0b;
    11'b00010010101: data <= 32'hbb15ba5a;
    11'b00010010110: data <= 32'hbc72b101;
    11'b00010010111: data <= 32'hbd1a3d90;
    11'b00010011000: data <= 32'hbec03e6e;
    11'b00010011001: data <= 32'hbdbcb023;
    11'b00010011010: data <= 32'hb2d5be7b;
    11'b00010011011: data <= 32'h39d6bb0d;
    11'b00010011100: data <= 32'h37cb3c74;
    11'b00010011101: data <= 32'h2b54400e;
    11'b00010011110: data <= 32'h398c3da9;
    11'b00010011111: data <= 32'h3e6339e8;
    11'b00010100000: data <= 32'h3bed3993;
    11'b00010100001: data <= 32'hbaa6365a;
    11'b00010100010: data <= 32'hbdd7b91a;
    11'b00010100011: data <= 32'h3249bd94;
    11'b00010100100: data <= 32'h4054bc61;
    11'b00010100101: data <= 32'h4039b89a;
    11'b00010100110: data <= 32'h37a4ba44;
    11'b00010100111: data <= 32'hb891bc04;
    11'b00010101000: data <= 32'hb681add1;
    11'b00010101001: data <= 32'hb6133cb6;
    11'b00010101010: data <= 32'hbccd3abc;
    11'b00010101011: data <= 32'hbf24bc82;
    11'b00010101100: data <= 32'hbce6c094;
    11'b00010101101: data <= 32'hb4ccbc2a;
    11'b00010101110: data <= 32'ha96c3c6a;
    11'b00010101111: data <= 32'ha83e3ef5;
    11'b00010110000: data <= 32'h38413b37;
    11'b00010110001: data <= 32'h3bed3852;
    11'b00010110010: data <= 32'h30083d1d;
    11'b00010110011: data <= 32'hbda03e89;
    11'b00010110100: data <= 32'hbdc438e7;
    11'b00010110101: data <= 32'h385eb9b6;
    11'b00010110110: data <= 32'h40b0bc0a;
    11'b00010110111: data <= 32'h3ffeb8dc;
    11'b00010111000: data <= 32'h380bb7d0;
    11'b00010111001: data <= 32'h2ee8b701;
    11'b00010111010: data <= 32'h3b2c3439;
    11'b00010111011: data <= 32'h3b6c3b97;
    11'b00010111100: data <= 32'hb85231d7;
    11'b00010111101: data <= 32'hbf7cbed4;
    11'b00010111110: data <= 32'hbe54c105;
    11'b00010111111: data <= 32'hb67ebcc2;
    11'b00011000000: data <= 32'h3119380c;
    11'b00011000001: data <= 32'h2c0c38a9;
    11'b00011000010: data <= 32'h2fe1b485;
    11'b00011000011: data <= 32'h30832788;
    11'b00011000100: data <= 32'hb9863e8b;
    11'b00011000101: data <= 32'hbf4440c9;
    11'b00011000110: data <= 32'hbe553c96;
    11'b00011000111: data <= 32'h31e4b8ab;
    11'b00011001000: data <= 32'h3e18bb5f;
    11'b00011001001: data <= 32'h3c68b006;
    11'b00011001010: data <= 32'h330f3658;
    11'b00011001011: data <= 32'h39e136b2;
    11'b00011001100: data <= 32'h400c3963;
    11'b00011001101: data <= 32'h3f5d3b96;
    11'b00011001110: data <= 32'hb17632b1;
    11'b00011001111: data <= 32'hbefcbd4f;
    11'b00011010000: data <= 32'hbccfbffc;
    11'b00011010001: data <= 32'h3578bc9a;
    11'b00011010010: data <= 32'h3b19b4e3;
    11'b00011010011: data <= 32'h3519ba2e;
    11'b00011010100: data <= 32'hb00cbdc1;
    11'b00011010101: data <= 32'hb293b73d;
    11'b00011010110: data <= 32'hb9f73e85;
    11'b00011010111: data <= 32'hbea9409a;
    11'b00011011000: data <= 32'hbef439a6;
    11'b00011011001: data <= 32'hb973bc45;
    11'b00011011010: data <= 32'h3094bbaa;
    11'b00011011011: data <= 32'hae353658;
    11'b00011011100: data <= 32'hb3423c5a;
    11'b00011011101: data <= 32'h3bb23a94;
    11'b00011011110: data <= 32'h40b13a22;
    11'b00011011111: data <= 32'h3f513cad;
    11'b00011100000: data <= 32'hb5a73bcf;
    11'b00011100001: data <= 32'hbe61af60;
    11'b00011100010: data <= 32'hb7ecbba6;
    11'b00011100011: data <= 32'h3d13bb07;
    11'b00011100100: data <= 32'h3e07ba93;
    11'b00011100101: data <= 32'h37dfbe1a;
    11'b00011100110: data <= 32'ha3e6bf81;
    11'b00011100111: data <= 32'h34dfb880;
    11'b00011101000: data <= 32'h31013d8a;
    11'b00011101001: data <= 32'hbb4e3e53;
    11'b00011101010: data <= 32'hbee7b44f;
    11'b00011101011: data <= 32'hbdf1befb;
    11'b00011101100: data <= 32'hbbb6bc46;
    11'b00011101101: data <= 32'hbb143857;
    11'b00011101110: data <= 32'hb84f3bbc;
    11'b00011101111: data <= 32'h39f33500;
    11'b00011110000: data <= 32'h3f353541;
    11'b00011110001: data <= 32'h3c163d97;
    11'b00011110010: data <= 32'hbb5e3ffd;
    11'b00011110011: data <= 32'hbe323cd6;
    11'b00011110100: data <= 32'ha858208f;
    11'b00011110101: data <= 32'h3e5ab835;
    11'b00011110110: data <= 32'h3da1ba27;
    11'b00011110111: data <= 32'h3502bd39;
    11'b00011111000: data <= 32'h3557bda0;
    11'b00011111001: data <= 32'h3d91b3b3;
    11'b00011111010: data <= 32'h3e213c92;
    11'b00011111011: data <= 32'h2a383aca;
    11'b00011111100: data <= 32'hbe06bbb6;
    11'b00011111101: data <= 32'hbeebbff7;
    11'b00011111110: data <= 32'hbc9fbc31;
    11'b00011111111: data <= 32'hba9433bd;
    11'b00100000000: data <= 32'hb81624d1;
    11'b00100000001: data <= 32'h3535bb77;
    11'b00100000010: data <= 32'h3b4db7d5;
    11'b00100000011: data <= 32'h2f7e3daf;
    11'b00100000100: data <= 32'hbd75413c;
    11'b00100000101: data <= 32'hbe3e3f59;
    11'b00100000110: data <= 32'hb04f352b;
    11'b00100000111: data <= 32'h3bbdb530;
    11'b00100001000: data <= 32'h3758b455;
    11'b00100001001: data <= 32'hb462b695;
    11'b00100001010: data <= 32'h38e7b7e1;
    11'b00100001011: data <= 32'h40b9329d;
    11'b00100001100: data <= 32'h41183c31;
    11'b00100001101: data <= 32'h39263938;
    11'b00100001110: data <= 32'hbcdfba2e;
    11'b00100001111: data <= 32'hbd44bdc3;
    11'b00100010000: data <= 32'hb6cbb9c7;
    11'b00100010001: data <= 32'hacbcb307;
    11'b00100010010: data <= 32'hb32ebcac;
    11'b00100010011: data <= 32'h2358c065;
    11'b00100010100: data <= 32'h361ebcef;
    11'b00100010101: data <= 32'haf6d3cd3;
    11'b00100010110: data <= 32'hbccb40f1;
    11'b00100010111: data <= 32'hbdd33dbe;
    11'b00100011000: data <= 32'hb942b079;
    11'b00100011001: data <= 32'hb3a2b5f7;
    11'b00100011010: data <= 32'hbad234aa;
    11'b00100011011: data <= 32'hbc0e36d1;
    11'b00100011100: data <= 32'h38b72cd1;
    11'b00100011101: data <= 32'h413834ef;
    11'b00100011110: data <= 32'h41313c2e;
    11'b00100011111: data <= 32'h383a3c60;
    11'b00100100000: data <= 32'hbc333428;
    11'b00100100001: data <= 32'hb8a2b4a4;
    11'b00100100010: data <= 32'h38eab05d;
    11'b00100100011: data <= 32'h3988b737;
    11'b00100100100: data <= 32'ha5c9bf54;
    11'b00100100101: data <= 32'hab78c170;
    11'b00100100110: data <= 32'h38bbbdd8;
    11'b00100100111: data <= 32'h38d03b3d;
    11'b00100101000: data <= 32'hb5913ee4;
    11'b00100101001: data <= 32'hbc7c3612;
    11'b00100101010: data <= 32'hbc9bbb84;
    11'b00100101011: data <= 32'hbcf8b830;
    11'b00100101100: data <= 32'hbeff38ab;
    11'b00100101101: data <= 32'hbdfb389d;
    11'b00100101110: data <= 32'h345fb3ee;
    11'b00100101111: data <= 32'h4011b2a6;
    11'b00100110000: data <= 32'h3ef43bad;
    11'b00100110001: data <= 32'hb03e3f28;
    11'b00100110010: data <= 32'hbc2f3de0;
    11'b00100110011: data <= 32'h9b3f3a6e;
    11'b00100110100: data <= 32'h3cb536fa;
    11'b00100110101: data <= 32'h3a3bb413;
    11'b00100110110: data <= 32'hb413be4c;
    11'b00100110111: data <= 32'h9ae5c077;
    11'b00100111000: data <= 32'h3d65bc54;
    11'b00100111001: data <= 32'h3f673996;
    11'b00100111010: data <= 32'h3a093b32;
    11'b00100111011: data <= 32'hb91bb83f;
    11'b00100111100: data <= 32'hbcd3bd7d;
    11'b00100111101: data <= 32'hbd8eb79e;
    11'b00100111110: data <= 32'hbed23865;
    11'b00100111111: data <= 32'hbdd4aa18;
    11'b00101000000: data <= 32'hb011bd6d;
    11'b00101000001: data <= 32'h3c4bbcad;
    11'b00101000010: data <= 32'h39283983;
    11'b00101000011: data <= 32'hba13405c;
    11'b00101000100: data <= 32'hbc3a4016;
    11'b00101000101: data <= 32'h30373cb1;
    11'b00101000110: data <= 32'h3af33976;
    11'b00101000111: data <= 32'ha5cf3413;
    11'b00101001000: data <= 32'hbbd5b8fa;
    11'b00101001001: data <= 32'ha88bbca3;
    11'b00101001010: data <= 32'h4020b75e;
    11'b00101001011: data <= 32'h419c3901;
    11'b00101001100: data <= 32'h3dc237fa;
    11'b00101001101: data <= 32'hb3eeb922;
    11'b00101001110: data <= 32'hb9f6bbd8;
    11'b00101001111: data <= 32'hb8dea71f;
    11'b00101010000: data <= 32'hbaa93678;
    11'b00101010001: data <= 32'hbc11bbaa;
    11'b00101010010: data <= 32'hb670c11c;
    11'b00101010011: data <= 32'h35e6c011;
    11'b00101010100: data <= 32'h2fd0350b;
    11'b00101010101: data <= 32'hba263fc9;
    11'b00101010110: data <= 32'hbad13e63;
    11'b00101010111: data <= 32'had1e3901;
    11'b00101011000: data <= 32'ha9fd381a;
    11'b00101011001: data <= 32'hbd0b3a3a;
    11'b00101011010: data <= 32'hbf7535cd;
    11'b00101011011: data <= 32'hb443b517;
    11'b00101011100: data <= 32'h405eb16b;
    11'b00101011101: data <= 32'h419f386a;
    11'b00101011110: data <= 32'h3d203924;
    11'b00101011111: data <= 32'hb1022dd8;
    11'b00101100000: data <= 32'ha8b42d95;
    11'b00101100001: data <= 32'h387139c1;
    11'b00101100010: data <= 32'h31f436bb;
    11'b00101100011: data <= 32'hb8edbdd8;
    11'b00101100100: data <= 32'hb81cc214;
    11'b00101100101: data <= 32'h34d3c086;
    11'b00101100110: data <= 32'h38462938;
    11'b00101100111: data <= 32'ha4473cd3;
    11'b00101101000: data <= 32'hb5a336ea;
    11'b00101101001: data <= 32'hb4b8b670;
    11'b00101101010: data <= 32'hbae33137;
    11'b00101101011: data <= 32'hc0413c54;
    11'b00101101100: data <= 32'hc0c93a1f;
    11'b00101101101: data <= 32'hb8e2b552;
    11'b00101101110: data <= 32'h3e5cb884;
    11'b00101101111: data <= 32'h3f7034f4;
    11'b00101110000: data <= 32'h36c13c29;
    11'b00101110001: data <= 32'hb57b3c57;
    11'b00101110010: data <= 32'h38433c9e;
    11'b00101110011: data <= 32'h3d623d89;
    11'b00101110100: data <= 32'h38a7399d;
    11'b00101110101: data <= 32'hb99fbca3;
    11'b00101110110: data <= 32'hb8c3c0f2;
    11'b00101110111: data <= 32'h3a09bee3;
    11'b00101111000: data <= 32'h3e2f185f;
    11'b00101111001: data <= 32'h3c3b365f;
    11'b00101111010: data <= 32'h342db97e;
    11'b00101111011: data <= 32'hb2c2bc90;
    11'b00101111100: data <= 32'hbb7b2984;
    11'b00101111101: data <= 32'hc00c3ca2;
    11'b00101111110: data <= 32'hc07a3710;
    11'b00101111111: data <= 32'hbb00bcbe;
    11'b00110000000: data <= 32'h3929bdf4;
    11'b00110000001: data <= 32'h389caf7a;
    11'b00110000010: data <= 32'hb80a3cfa;
    11'b00110000011: data <= 32'hb84f3e3b;
    11'b00110000100: data <= 32'h3a043df1;
    11'b00110000101: data <= 32'h3d533e45;
    11'b00110000110: data <= 32'h2a903c79;
    11'b00110000111: data <= 32'hbd80b2e9;
    11'b00110001000: data <= 32'hba5dbcec;
    11'b00110001001: data <= 32'h3cf9ba7f;
    11'b00110001010: data <= 32'h40be3021;
    11'b00110001011: data <= 32'h3ee2abf1;
    11'b00110001100: data <= 32'h3924bc53;
    11'b00110001101: data <= 32'h32b6bc24;
    11'b00110001110: data <= 32'hb0d436b1;
    11'b00110001111: data <= 32'hbc033cba;
    11'b00110010000: data <= 32'hbe20b2fd;
    11'b00110010001: data <= 32'hbb93c077;
    11'b00110010010: data <= 32'hae43c0b0;
    11'b00110010011: data <= 32'hb311b844;
    11'b00110010100: data <= 32'hba893bf8;
    11'b00110010101: data <= 32'hb6f13c5d;
    11'b00110010110: data <= 32'h399b3a84;
    11'b00110010111: data <= 32'h39773ca9;
    11'b00110011000: data <= 32'hbc103dca;
    11'b00110011001: data <= 32'hc0843a54;
    11'b00110011010: data <= 32'hbc74b009;
    11'b00110011011: data <= 32'h3d32b27a;
    11'b00110011100: data <= 32'h40ad31ea;
    11'b00110011101: data <= 32'h3dddac0c;
    11'b00110011110: data <= 32'h3861b908;
    11'b00110011111: data <= 32'h39fbb12b;
    11'b00110100000: data <= 32'h3c1b3caa;
    11'b00110100001: data <= 32'h34383d49;
    11'b00110100010: data <= 32'hba6eb8e1;
    11'b00110100011: data <= 32'hbb32c152;
    11'b00110100100: data <= 32'hb4a2c102;
    11'b00110100101: data <= 32'hae58b960;
    11'b00110100110: data <= 32'hb48e3646;
    11'b00110100111: data <= 32'h2b73ad9a;
    11'b00110101000: data <= 32'h3913b71e;
    11'b00110101001: data <= 32'h253737db;
    11'b00110101010: data <= 32'hbf3d3e48;
    11'b00110101011: data <= 32'hc17f3d2f;
    11'b00110101100: data <= 32'hbd8130f8;
    11'b00110101101: data <= 32'h3a68b596;
    11'b00110101110: data <= 32'h3d7aa7b5;
    11'b00110101111: data <= 32'h3657317e;
    11'b00110110000: data <= 32'h2a6731bc;
    11'b00110110001: data <= 32'h3c803a8d;
    11'b00110110010: data <= 32'h3f9b3f47;
    11'b00110110011: data <= 32'h3ba83e4e;
    11'b00110110100: data <= 32'hb8e8b5c1;
    11'b00110110101: data <= 32'hbb66c025;
    11'b00110110110: data <= 32'h96a0bf1e;
    11'b00110110111: data <= 32'h3995b6c6;
    11'b00110111000: data <= 32'h3976b333;
    11'b00110111001: data <= 32'h3973bd1b;
    11'b00110111010: data <= 32'h39f6bdec;
    11'b00110111011: data <= 32'habdb2c60;
    11'b00110111100: data <= 32'hbeba3e3c;
    11'b00110111101: data <= 32'hc0e23c86;
    11'b00110111110: data <= 32'hbd8eb759;
    11'b00110111111: data <= 32'h288abc91;
    11'b00111000000: data <= 32'h25f5b79c;
    11'b00111000001: data <= 32'hba9d34db;
    11'b00111000010: data <= 32'hb78138ef;
    11'b00111000011: data <= 32'h3ce93c7d;
    11'b00111000100: data <= 32'h40113f8e;
    11'b00111000101: data <= 32'h397c3f25;
    11'b00111000110: data <= 32'hbc8036c5;
    11'b00111000111: data <= 32'hbc91ba32;
    11'b00111001000: data <= 32'h3619b8a5;
    11'b00111001001: data <= 32'h3dca28fd;
    11'b00111001010: data <= 32'h3d41b85a;
    11'b00111001011: data <= 32'h3becbf3c;
    11'b00111001100: data <= 32'h3c0ebe9e;
    11'b00111001101: data <= 32'h38b83401;
    11'b00111001110: data <= 32'hb8e83e58;
    11'b00111001111: data <= 32'hbdd938cb;
    11'b00111010000: data <= 32'hbc7ebd94;
    11'b00111010001: data <= 32'hb862bfd3;
    11'b00111010010: data <= 32'hbb39bad8;
    11'b00111010011: data <= 32'hbdbf30d3;
    11'b00111010100: data <= 32'hb8bd33f2;
    11'b00111010101: data <= 32'h3ca33692;
    11'b00111010110: data <= 32'h3e1d3cf7;
    11'b00111010111: data <= 32'hb39e3f29;
    11'b00111011000: data <= 32'hbfd23d0a;
    11'b00111011001: data <= 32'hbdce3738;
    11'b00111011010: data <= 32'h37ab3581;
    11'b00111011011: data <= 32'h3de935c2;
    11'b00111011100: data <= 32'h3c1ab807;
    11'b00111011101: data <= 32'h397abe07;
    11'b00111011110: data <= 32'h3d03bba1;
    11'b00111011111: data <= 32'h3e653b69;
    11'b00111100000: data <= 32'h3a213ef2;
    11'b00111100001: data <= 32'hb68932b9;
    11'b00111100010: data <= 32'hba36bf68;
    11'b00111100011: data <= 32'hb95cc02e;
    11'b00111100100: data <= 32'hbb7eba9a;
    11'b00111100101: data <= 32'hbc71b234;
    11'b00111100110: data <= 32'hb254ba2a;
    11'b00111100111: data <= 32'h3c75bb9d;
    11'b00111101000: data <= 32'h3b3f33a9;
    11'b00111101001: data <= 32'hbc203e5a;
    11'b00111101010: data <= 32'hc0da3eac;
    11'b00111101011: data <= 32'hbe5a3b20;
    11'b00111101100: data <= 32'h32433705;
    11'b00111101101: data <= 32'h3934346f;
    11'b00111101110: data <= 32'hb065b49f;
    11'b00111101111: data <= 32'hb02fba2d;
    11'b00111110000: data <= 32'h3d2e9cad;
    11'b00111110001: data <= 32'h40b53e45;
    11'b00111110010: data <= 32'h3e793fa2;
    11'b00111110011: data <= 32'h2b4234b0;
    11'b00111110100: data <= 32'hb906bd8d;
    11'b00111110101: data <= 32'hb63fbd23;
    11'b00111110110: data <= 32'hb3a9b472;
    11'b00111110111: data <= 32'hb2a3b7a2;
    11'b00111111000: data <= 32'h3697bf51;
    11'b00111111001: data <= 32'h3cb8c04a;
    11'b00111111010: data <= 32'h39a1b7cc;
    11'b00111111011: data <= 32'hbc073d71;
    11'b00111111100: data <= 32'hc01c3df8;
    11'b00111111101: data <= 32'hbd533657;
    11'b00111111110: data <= 32'hb3fdb40a;
    11'b00111111111: data <= 32'hb87db099;
    11'b01000000000: data <= 32'hbe12b090;
    11'b01000000001: data <= 32'hbbd1b429;
    11'b01000000010: data <= 32'h3c91361f;
    11'b01000000011: data <= 32'h40e83e60;
    11'b01000000100: data <= 32'h3def3f8c;
    11'b01000000101: data <= 32'hb5033a3c;
    11'b01000000110: data <= 32'hba61b31c;
    11'b01000000111: data <= 32'ha20e2c74;
    11'b01000001000: data <= 32'h38563838;
    11'b01000001001: data <= 32'h37c3b814;
    11'b01000001010: data <= 32'h3997c09e;
    11'b01000001011: data <= 32'h3d0dc0f1;
    11'b01000001100: data <= 32'h3c5db7cf;
    11'b01000001101: data <= 32'hac733d3c;
    11'b01000001110: data <= 32'hbb713bc5;
    11'b01000001111: data <= 32'hb9bbb847;
    11'b01000010000: data <= 32'hb832bc69;
    11'b01000010001: data <= 32'hbdadb823;
    11'b01000010010: data <= 32'hc097b0fe;
    11'b01000010011: data <= 32'hbd4eb671;
    11'b01000010100: data <= 32'h3ba9b277;
    11'b01000010101: data <= 32'h3fd33a8b;
    11'b01000010110: data <= 32'h38c03e34;
    11'b01000010111: data <= 32'hbc9b3d2f;
    11'b01000011000: data <= 32'hbc6f3b63;
    11'b01000011001: data <= 32'h31e13cb5;
    11'b01000011010: data <= 32'h3a113c77;
    11'b01000011011: data <= 32'h3515b4fe;
    11'b01000011100: data <= 32'h34a1c005;
    11'b01000011101: data <= 32'h3cbdbf55;
    11'b01000011110: data <= 32'h3f1e3136;
    11'b01000011111: data <= 32'h3ce23dd5;
    11'b01000100000: data <= 32'h35123825;
    11'b01000100001: data <= 32'hac01bc8e;
    11'b01000100010: data <= 32'hb72cbd66;
    11'b01000100011: data <= 32'hbdc9b68f;
    11'b01000100100: data <= 32'hc020b2fc;
    11'b01000100101: data <= 32'hbbf8bc75;
    11'b01000100110: data <= 32'h3b32bddf;
    11'b01000100111: data <= 32'h3d2eb614;
    11'b01000101000: data <= 32'hb4f93c0c;
    11'b01000101001: data <= 32'hbee63ddf;
    11'b01000101010: data <= 32'hbcc73d63;
    11'b01000101011: data <= 32'h30923d96;
    11'b01000101100: data <= 32'h32f43c95;
    11'b01000101101: data <= 32'hb9f6ac08;
    11'b01000101110: data <= 32'hb9b9bd03;
    11'b01000101111: data <= 32'h3affba74;
    11'b01000110000: data <= 32'h408a3b26;
    11'b01000110001: data <= 32'h40173e69;
    11'b01000110010: data <= 32'h3b813662;
    11'b01000110011: data <= 32'h33febb7e;
    11'b01000110100: data <= 32'hae8bb92d;
    11'b01000110101: data <= 32'hb9eb3500;
    11'b01000110110: data <= 32'hbc78b0c0;
    11'b01000110111: data <= 32'hb506bf8e;
    11'b01000111000: data <= 32'h3babc141;
    11'b01000111001: data <= 32'h3b72bd28;
    11'b01000111010: data <= 32'hb830388c;
    11'b01000111011: data <= 32'hbdda3cbf;
    11'b01000111100: data <= 32'hba443ac9;
    11'b01000111101: data <= 32'h290e399b;
    11'b01000111110: data <= 32'hb9a03972;
    11'b01000111111: data <= 32'hc02b2d14;
    11'b01001000000: data <= 32'hbf0fb8ec;
    11'b01001000001: data <= 32'h3758b2a7;
    11'b01001000010: data <= 32'h40733c26;
    11'b01001000011: data <= 32'h3fa23dd4;
    11'b01001000100: data <= 32'h38d23883;
    11'b01001000101: data <= 32'h2cd2abf8;
    11'b01001000110: data <= 32'h3464394a;
    11'b01001000111: data <= 32'h305d3d58;
    11'b01001001000: data <= 32'hb3b72f9e;
    11'b01001001001: data <= 32'h2e2fc061;
    11'b01001001010: data <= 32'h3b98c1e6;
    11'b01001001011: data <= 32'h3c19bd75;
    11'b01001001100: data <= 32'h30123795;
    11'b01001001101: data <= 32'hb6463939;
    11'b01001001110: data <= 32'h2af2b0ea;
    11'b01001001111: data <= 32'h2debb4d8;
    11'b01001010000: data <= 32'hbd6b31e0;
    11'b01001010001: data <= 32'hc1ba2fff;
    11'b01001010010: data <= 32'hc076b7fe;
    11'b01001010011: data <= 32'h31c8b81b;
    11'b01001010100: data <= 32'h3ec33546;
    11'b01001010101: data <= 32'h3bbb3b3b;
    11'b01001010110: data <= 32'hb5ac39e5;
    11'b01001010111: data <= 32'hb5963ad6;
    11'b01001011000: data <= 32'h38063f17;
    11'b01001011001: data <= 32'h38994029;
    11'b01001011010: data <= 32'hb083376c;
    11'b01001011011: data <= 32'hb34abf4d;
    11'b01001011100: data <= 32'h3965c08c;
    11'b01001011101: data <= 32'h3d76b90c;
    11'b01001011110: data <= 32'h3cb039bc;
    11'b01001011111: data <= 32'h3ae331d5;
    11'b01001100000: data <= 32'h3b36bb94;
    11'b01001100001: data <= 32'h35e5ba6a;
    11'b01001100010: data <= 32'hbd283205;
    11'b01001100011: data <= 32'hc1373369;
    11'b01001100100: data <= 32'hbf6fbafc;
    11'b01001100101: data <= 32'h31fabe17;
    11'b01001100110: data <= 32'h3c11baf5;
    11'b01001100111: data <= 32'hae6f30a0;
    11'b01001101000: data <= 32'hbca9394a;
    11'b01001101001: data <= 32'hb86c3ca0;
    11'b01001101010: data <= 32'h38cb3ff3;
    11'b01001101011: data <= 32'h35a7403c;
    11'b01001101100: data <= 32'hbb853981;
    11'b01001101101: data <= 32'hbce5bc38;
    11'b01001101110: data <= 32'h301dbc71;
    11'b01001101111: data <= 32'h3e493518;
    11'b01001110000: data <= 32'h3f653bec;
    11'b01001110001: data <= 32'h3df8a97e;
    11'b01001110010: data <= 32'h3d18bc2a;
    11'b01001110011: data <= 32'h39e7b5de;
    11'b01001110100: data <= 32'hb8763b18;
    11'b01001110101: data <= 32'hbe32384d;
    11'b01001110110: data <= 32'hbbdbbd5a;
    11'b01001110111: data <= 32'h360dc105;
    11'b01001111000: data <= 32'h3897bf36;
    11'b01001111001: data <= 32'hb8b5b695;
    11'b01001111010: data <= 32'hbcb134d4;
    11'b01001111011: data <= 32'hb1ec38f0;
    11'b01001111100: data <= 32'h39c63cd1;
    11'b01001111101: data <= 32'hb3d63df7;
    11'b01001111110: data <= 32'hc02e39a3;
    11'b01001111111: data <= 32'hc09db5c3;
    11'b01010000000: data <= 32'hb71eb424;
    11'b01010000001: data <= 32'h3d9339e2;
    11'b01010000010: data <= 32'h3e993b49;
    11'b01010000011: data <= 32'h3c63ad77;
    11'b01010000100: data <= 32'h3bdcb7e6;
    11'b01010000101: data <= 32'h3c0839e8;
    11'b01010000110: data <= 32'h35c13fca;
    11'b01010000111: data <= 32'hb7183bff;
    11'b01010001000: data <= 32'hb4c5bdd5;
    11'b01010001001: data <= 32'h3763c180;
    11'b01010001010: data <= 32'h37c4bf61;
    11'b01010001011: data <= 32'hb431b70c;
    11'b01010001100: data <= 32'hb51db117;
    11'b01010001101: data <= 32'h3980b6b6;
    11'b01010001110: data <= 32'h3bf79c88;
    11'b01010001111: data <= 32'hb96939d2;
    11'b01010010000: data <= 32'hc18a3914;
    11'b01010010001: data <= 32'hc187adc1;
    11'b01010010010: data <= 32'hb9b4b3da;
    11'b01010010011: data <= 32'h3b203430;
    11'b01010010100: data <= 32'h395e355b;
    11'b01010010101: data <= 32'ha902b0c2;
    11'b01010010110: data <= 32'h34ee317d;
    11'b01010010111: data <= 32'h3c6e3ef3;
    11'b01010011000: data <= 32'h3b66416d;
    11'b01010011001: data <= 32'ha84e3d8f;
    11'b01010011010: data <= 32'hb5ebbc50;
    11'b01010011011: data <= 32'h31eec011;
    11'b01010011100: data <= 32'h38b2bbae;
    11'b01010011101: data <= 32'h380c2683;
    11'b01010011110: data <= 32'h3a73b7fb;
    11'b01010011111: data <= 32'h3e50bd45;
    11'b01010100000: data <= 32'h3d7cba68;
    11'b01010100001: data <= 32'hb8643769;
    11'b01010100010: data <= 32'hc0ee39b7;
    11'b01010100011: data <= 32'hc08cb37a;
    11'b01010100100: data <= 32'hb829bbad;
    11'b01010100101: data <= 32'h3566ba59;
    11'b01010100110: data <= 32'hb7c0b7c0;
    11'b01010100111: data <= 32'hbc88b5f4;
    11'b01010101000: data <= 32'hb1a735dd;
    11'b01010101001: data <= 32'h3c963f96;
    11'b01010101010: data <= 32'h3b534155;
    11'b01010101011: data <= 32'hb8373de4;
    11'b01010101100: data <= 32'hbcceb686;
    11'b01010101101: data <= 32'hb6c9ba51;
    11'b01010101110: data <= 32'h38d93420;
    11'b01010101111: data <= 32'h3c2338ae;
    11'b01010110000: data <= 32'h3d84b922;
    11'b01010110001: data <= 32'h3fa2be6a;
    11'b01010110010: data <= 32'h3e9db96c;
    11'b01010110011: data <= 32'h2f173bca;
    11'b01010110100: data <= 32'hbd573c4d;
    11'b01010110101: data <= 32'hbc97b7ce;
    11'b01010110110: data <= 32'ha9bcbf0d;
    11'b01010110111: data <= 32'h9ceebea4;
    11'b01010111000: data <= 32'hbc96bc26;
    11'b01010111001: data <= 32'hbdd6b9a3;
    11'b01010111010: data <= 32'ha590b05c;
    11'b01010111011: data <= 32'h3d3c3c33;
    11'b01010111100: data <= 32'h38523f46;
    11'b01010111101: data <= 32'hbddb3ce0;
    11'b01010111110: data <= 32'hc06a3192;
    11'b01010111111: data <= 32'hbc1c330d;
    11'b01011000000: data <= 32'h365c3bfa;
    11'b01011000001: data <= 32'h3aa839f6;
    11'b01011000010: data <= 32'h3b68b99a;
    11'b01011000011: data <= 32'h3dbabd21;
    11'b01011000100: data <= 32'h3eb9320f;
    11'b01011000101: data <= 32'h3b4f3fc7;
    11'b01011000110: data <= 32'had7c3e5e;
    11'b01011000111: data <= 32'hb076b832;
    11'b01011001000: data <= 32'h34dbbfd8;
    11'b01011001001: data <= 32'had48be9a;
    11'b01011001010: data <= 32'hbc2dbb65;
    11'b01011001011: data <= 32'hbaebbbb3;
    11'b01011001100: data <= 32'h39f4bc45;
    11'b01011001101: data <= 32'h3e9ab49e;
    11'b01011001110: data <= 32'h338039e1;
    11'b01011001111: data <= 32'hc0213ae8;
    11'b01011010000: data <= 32'hc13d367e;
    11'b01011010001: data <= 32'hbccc373f;
    11'b01011010010: data <= 32'h29fc3a72;
    11'b01011010011: data <= 32'habaf34ca;
    11'b01011010100: data <= 32'hb53ebab1;
    11'b01011010101: data <= 32'h3739ba34;
    11'b01011010110: data <= 32'h3def3c51;
    11'b01011010111: data <= 32'h3da94156;
    11'b01011011000: data <= 32'h38473fba;
    11'b01011011001: data <= 32'h2dfcb3d0;
    11'b01011011010: data <= 32'h320ebd37;
    11'b01011011011: data <= 32'ha9fdb948;
    11'b01011011100: data <= 32'hb75eb1a1;
    11'b01011011101: data <= 32'h2fdfbc0a;
    11'b01011011110: data <= 32'h3e63bf8a;
    11'b01011011111: data <= 32'h4009bd25;
    11'b01011100000: data <= 32'h350f30aa;
    11'b01011100001: data <= 32'hbf2f39f6;
    11'b01011100010: data <= 32'hc01234fa;
    11'b01011100011: data <= 32'hba0dab94;
    11'b01011100100: data <= 32'hb36dad30;
    11'b01011100101: data <= 32'hbc84b7a5;
    11'b01011100110: data <= 32'hbe75bc5a;
    11'b01011100111: data <= 32'hb5f1b8b0;
    11'b01011101000: data <= 32'h3d2a3cff;
    11'b01011101001: data <= 32'h3dba4119;
    11'b01011101010: data <= 32'h34143f37;
    11'b01011101011: data <= 32'hb84b31cc;
    11'b01011101100: data <= 32'hb5d4b0a3;
    11'b01011101101: data <= 32'had4b39f0;
    11'b01011101110: data <= 32'h23a039d6;
    11'b01011101111: data <= 32'h3973bb27;
    11'b01011110000: data <= 32'h3f7fc059;
    11'b01011110001: data <= 32'h4046bd88;
    11'b01011110010: data <= 32'h3a2336c6;
    11'b01011110011: data <= 32'hb9f13c1b;
    11'b01011110100: data <= 32'hb9e43001;
    11'b01011110101: data <= 32'h2c1dba26;
    11'b01011110110: data <= 32'hb4bdbb42;
    11'b01011110111: data <= 32'hbf18bbf9;
    11'b01011111000: data <= 32'hc054bd3d;
    11'b01011111001: data <= 32'hb7b5bb66;
    11'b01011111010: data <= 32'h3d5d3785;
    11'b01011111011: data <= 32'h3c803e2b;
    11'b01011111100: data <= 32'hb8733cdd;
    11'b01011111101: data <= 32'hbde6379e;
    11'b01011111110: data <= 32'hbb933aaa;
    11'b01011111111: data <= 32'hb3603ed8;
    11'b01100000000: data <= 32'hac8d3cbe;
    11'b01100000001: data <= 32'h348dba73;
    11'b01100000010: data <= 32'h3d0cbfa7;
    11'b01100000011: data <= 32'h3f6cb956;
    11'b01100000100: data <= 32'h3d253d30;
    11'b01100000101: data <= 32'h37713e19;
    11'b01100000110: data <= 32'h380d2c79;
    11'b01100000111: data <= 32'h39eabc23;
    11'b01100001000: data <= 32'hb227bb85;
    11'b01100001001: data <= 32'hbee3ba35;
    11'b01100001010: data <= 32'hbefabd2f;
    11'b01100001011: data <= 32'h30f5be59;
    11'b01100001100: data <= 32'h3ea4ba8f;
    11'b01100001101: data <= 32'h3aab3332;
    11'b01100001110: data <= 32'hbcb93813;
    11'b01100001111: data <= 32'hbfa837df;
    11'b01100010000: data <= 32'hbc273c6a;
    11'b01100010001: data <= 32'hb5b23edd;
    11'b01100010010: data <= 32'hb9c63b40;
    11'b01100010011: data <= 32'hbb57bb3c;
    11'b01100010100: data <= 32'h2b24bdc6;
    11'b01100010101: data <= 32'h3d2e32af;
    11'b01100010110: data <= 32'h3e2d4011;
    11'b01100010111: data <= 32'h3c713f3e;
    11'b01100011000: data <= 32'h3bab3196;
    11'b01100011001: data <= 32'h3aaab8af;
    11'b01100011010: data <= 32'hae099221;
    11'b01100011011: data <= 32'hbcc131d9;
    11'b01100011100: data <= 32'hba71bbdb;
    11'b01100011101: data <= 32'h3c03c049;
    11'b01100011110: data <= 32'h3ffcbf53;
    11'b01100011111: data <= 32'h3a4cb8d3;
    11'b01100100000: data <= 32'hbc55306c;
    11'b01100100001: data <= 32'hbd8634d7;
    11'b01100100010: data <= 32'hb6853931;
    11'b01100100011: data <= 32'hb4a13b4e;
    11'b01100100100: data <= 32'hbe1830ff;
    11'b01100100101: data <= 32'hc06abc91;
    11'b01100100110: data <= 32'hbc15bcae;
    11'b01100100111: data <= 32'h3a77381f;
    11'b01100101000: data <= 32'h3db63fd9;
    11'b01100101001: data <= 32'h3b1b3e18;
    11'b01100101010: data <= 32'h37253481;
    11'b01100101011: data <= 32'h356834ff;
    11'b01100101100: data <= 32'hafdb3d99;
    11'b01100101101: data <= 32'hb9593d67;
    11'b01100101110: data <= 32'hb0aab84d;
    11'b01100101111: data <= 32'h3d52c087;
    11'b01100110000: data <= 32'h3ff6bfed;
    11'b01100110001: data <= 32'h3ba4b7a8;
    11'b01100110010: data <= 32'hb4763522;
    11'b01100110011: data <= 32'had8e2e8c;
    11'b01100110100: data <= 32'h396dacac;
    11'b01100110101: data <= 32'h997d2556;
    11'b01100110110: data <= 32'hbfe3b699;
    11'b01100110111: data <= 32'hc19ebd18;
    11'b01100111000: data <= 32'hbd45bd11;
    11'b01100111001: data <= 32'h39b5a842;
    11'b01100111010: data <= 32'h3c5b3bc1;
    11'b01100111011: data <= 32'h2d9b3969;
    11'b01100111100: data <= 32'hb82b32d8;
    11'b01100111101: data <= 32'hb4943c4c;
    11'b01100111110: data <= 32'hb2db40d6;
    11'b01100111111: data <= 32'hb879400d;
    11'b01101000000: data <= 32'hb551b421;
    11'b01101000001: data <= 32'h39f1bfc7;
    11'b01101000010: data <= 32'h3ddfbd2a;
    11'b01101000011: data <= 32'h3c723636;
    11'b01101000100: data <= 32'h399a3ac1;
    11'b01101000101: data <= 32'h3cd323bd;
    11'b01101000110: data <= 32'h3e69b7d7;
    11'b01101000111: data <= 32'h3570b257;
    11'b01101001000: data <= 32'hbf55b354;
    11'b01101001001: data <= 32'hc0dabc32;
    11'b01101001010: data <= 32'hb9cebe53;
    11'b01101001011: data <= 32'h3c20bc5a;
    11'b01101001100: data <= 32'h3a38b658;
    11'b01101001101: data <= 32'hb932b4dd;
    11'b01101001110: data <= 32'hbc7baab5;
    11'b01101001111: data <= 32'hb6d93cec;
    11'b01101010000: data <= 32'hb14940f2;
    11'b01101010001: data <= 32'hbb1a3f55;
    11'b01101010010: data <= 32'hbd32b527;
    11'b01101010011: data <= 32'hb809bdd5;
    11'b01101010100: data <= 32'h38f3b55a;
    11'b01101010101: data <= 32'h3c343d09;
    11'b01101010110: data <= 32'h3cd23cc1;
    11'b01101010111: data <= 32'h3ee1a461;
    11'b01101011000: data <= 32'h3f50b543;
    11'b01101011001: data <= 32'h381c3818;
    11'b01101011010: data <= 32'hbd1c3a12;
    11'b01101011011: data <= 32'hbdbcb724;
    11'b01101011100: data <= 32'h3355bf2e;
    11'b01101011101: data <= 32'h3db9bfbd;
    11'b01101011110: data <= 32'h3908bd30;
    11'b01101011111: data <= 32'hba70bad6;
    11'b01101100000: data <= 32'hba75b5df;
    11'b01101100001: data <= 32'h32f339ec;
    11'b01101100010: data <= 32'h31b43e92;
    11'b01101100011: data <= 32'hbd5a3c08;
    11'b01101100100: data <= 32'hc0d1b8f3;
    11'b01101100101: data <= 32'hbea6bc72;
    11'b01101100110: data <= 32'hadd73217;
    11'b01101100111: data <= 32'h3a123d98;
    11'b01101101000: data <= 32'h3b6e3b40;
    11'b01101101001: data <= 32'h3cd4b147;
    11'b01101101010: data <= 32'h3d313312;
    11'b01101101011: data <= 32'h370c3ee3;
    11'b01101101100: data <= 32'hb9a84006;
    11'b01101101101: data <= 32'hb8b43419;
    11'b01101101110: data <= 32'h3a11bec4;
    11'b01101101111: data <= 32'h3dcdc005;
    11'b01101110000: data <= 32'h3892bcc9;
    11'b01101110001: data <= 32'hb55eb97a;
    11'b01101110010: data <= 32'h34a2b864;
    11'b01101110011: data <= 32'h3d8da4c2;
    11'b01101110100: data <= 32'h39fc38c5;
    11'b01101110101: data <= 32'hbe1633f9;
    11'b01101110110: data <= 32'hc1d4ba61;
    11'b01101110111: data <= 32'hc003bc11;
    11'b01101111000: data <= 32'hb405a909;
    11'b01101111001: data <= 32'h366338dd;
    11'b01101111010: data <= 32'h2e0fa4b8;
    11'b01101111011: data <= 32'h2f7ab83b;
    11'b01101111100: data <= 32'h38063983;
    11'b01101111101: data <= 32'h34904142;
    11'b01101111110: data <= 32'hb7114183;
    11'b01101111111: data <= 32'hb7a1393d;
    11'b01110000000: data <= 32'h3615bd3a;
    11'b01110000001: data <= 32'h3aecbd20;
    11'b01110000010: data <= 32'h36e2b3a1;
    11'b01110000011: data <= 32'h3546a499;
    11'b01110000100: data <= 32'h3dd6b887;
    11'b01110000101: data <= 32'h40ceb878;
    11'b01110000110: data <= 32'h3d0a2ea3;
    11'b01110000111: data <= 32'hbd1632eb;
    11'b01110001000: data <= 32'hc0f8b848;
    11'b01110001001: data <= 32'hbd6abc2d;
    11'b01110001010: data <= 32'h3192ba26;
    11'b01110001011: data <= 32'h30ddb8fb;
    11'b01110001100: data <= 32'hb9ebbc6f;
    11'b01110001101: data <= 32'hb9d8bc0c;
    11'b01110001110: data <= 32'h30833981;
    11'b01110001111: data <= 32'h357c4142;
    11'b01110010000: data <= 32'hb80c4112;
    11'b01110010001: data <= 32'hbc763838;
    11'b01110010010: data <= 32'hb9c1baed;
    11'b01110010011: data <= 32'hae80b3d7;
    11'b01110010100: data <= 32'h2f4d3ad8;
    11'b01110010101: data <= 32'h3917385d;
    11'b01110010110: data <= 32'h3fa6b8a2;
    11'b01110010111: data <= 32'h4146b910;
    11'b01110011000: data <= 32'h3db037d4;
    11'b01110011001: data <= 32'hb9e03c2a;
    11'b01110011010: data <= 32'hbdb131d5;
    11'b01110011011: data <= 32'hb26fbbcf;
    11'b01110011100: data <= 32'h3a46bd87;
    11'b01110011101: data <= 32'h2993bdd4;
    11'b01110011110: data <= 32'hbc67bed3;
    11'b01110011111: data <= 32'hb9debd7c;
    11'b01110100000: data <= 32'h38dc31dd;
    11'b01110100001: data <= 32'h3a4c3ef2;
    11'b01110100010: data <= 32'hb94e3e2b;
    11'b01110100011: data <= 32'hbfda2864;
    11'b01110100100: data <= 32'hbf36b896;
    11'b01110100101: data <= 32'hbb27375b;
    11'b01110100110: data <= 32'hb4873d34;
    11'b01110100111: data <= 32'h34e53751;
    11'b01110101000: data <= 32'h3d60ba73;
    11'b01110101001: data <= 32'h3fe7b5ff;
    11'b01110101010: data <= 32'h3cb63dac;
    11'b01110101011: data <= 32'hb32a406b;
    11'b01110101100: data <= 32'hb6b73bf5;
    11'b01110101101: data <= 32'h38ffb9b3;
    11'b01110101110: data <= 32'h3c0ebd72;
    11'b01110101111: data <= 32'hac48bd39;
    11'b01110110000: data <= 32'hbb4fbdc9;
    11'b01110110001: data <= 32'h2c88bdaf;
    11'b01110110010: data <= 32'h3ebbb82a;
    11'b01110110011: data <= 32'h3def386c;
    11'b01110110100: data <= 32'hb92237ff;
    11'b01110110101: data <= 32'hc0abb5ea;
    11'b01110110110: data <= 32'hc032b744;
    11'b01110110111: data <= 32'hbc0a37f7;
    11'b01110111000: data <= 32'hb87b3a80;
    11'b01110111001: data <= 32'hb7d2b5b6;
    11'b01110111010: data <= 32'h304dbd37;
    11'b01110111011: data <= 32'h3b51b0a3;
    11'b01110111100: data <= 32'h3a514051;
    11'b01110111101: data <= 32'h28f941d3;
    11'b01110111110: data <= 32'hab6b3d94;
    11'b01110111111: data <= 32'h3876b5a9;
    11'b01111000000: data <= 32'h387cb92d;
    11'b01111000001: data <= 32'hb56ab3cf;
    11'b01111000010: data <= 32'hb814b854;
    11'b01111000011: data <= 32'h3c30bcd6;
    11'b01111000100: data <= 32'h4151bc24;
    11'b01111000101: data <= 32'h4015b178;
    11'b01111000110: data <= 32'hb5c330b8;
    11'b01111000111: data <= 32'hbf8eb43b;
    11'b01111001000: data <= 32'hbd6db5d8;
    11'b01111001001: data <= 32'hb61a2991;
    11'b01111001010: data <= 32'hb8c5b274;
    11'b01111001011: data <= 32'hbd25bda1;
    11'b01111001100: data <= 32'hbb66bf7c;
    11'b01111001101: data <= 32'h3357b366;
    11'b01111001110: data <= 32'h394c403a;
    11'b01111001111: data <= 32'h2c57413b;
    11'b01111010000: data <= 32'hb6a73c6c;
    11'b01111010001: data <= 32'hb4d5ae03;
    11'b01111010010: data <= 32'hb5c8359f;
    11'b01111010011: data <= 32'hba293c2d;
    11'b01111010100: data <= 32'hb567357f;
    11'b01111010101: data <= 32'h3db6bc0d;
    11'b01111010110: data <= 32'h41acbcb4;
    11'b01111010111: data <= 32'h402dac1a;
    11'b01111011000: data <= 32'h288039ae;
    11'b01111011001: data <= 32'hbadc364a;
    11'b01111011010: data <= 32'ha68fb12e;
    11'b01111011011: data <= 32'h3856b648;
    11'b01111011100: data <= 32'hb7a9bb7e;
    11'b01111011101: data <= 32'hbebfbfdf;
    11'b01111011110: data <= 32'hbcccc056;
    11'b01111011111: data <= 32'h3699b921;
    11'b01111100000: data <= 32'h3c173cf5;
    11'b01111100001: data <= 32'h2a803dd7;
    11'b01111100010: data <= 32'hbc36350a;
    11'b01111100011: data <= 32'hbd0aa858;
    11'b01111100100: data <= 32'hbc873c4d;
    11'b01111100101: data <= 32'hbca33f05;
    11'b01111100110: data <= 32'hb9003878;
    11'b01111100111: data <= 32'h3ae7bc82;
    11'b01111101000: data <= 32'h4010bc33;
    11'b01111101001: data <= 32'h3e4a390c;
    11'b01111101010: data <= 32'h35173ee9;
    11'b01111101011: data <= 32'h30d93cc5;
    11'b01111101100: data <= 32'h3c3c3090;
    11'b01111101101: data <= 32'h3c5fb5c7;
    11'b01111101110: data <= 32'hb725ba30;
    11'b01111101111: data <= 32'hbe79be60;
    11'b01111110000: data <= 32'hb929bff1;
    11'b01111110001: data <= 32'h3d3ebc88;
    11'b01111110010: data <= 32'h3ed32b7d;
    11'b01111110011: data <= 32'h30db314c;
    11'b01111110100: data <= 32'hbd73b6cb;
    11'b01111110101: data <= 32'hbe1bad8c;
    11'b01111110110: data <= 32'hbca73cdd;
    11'b01111110111: data <= 32'hbd023e1c;
    11'b01111111000: data <= 32'hbcf2aac2;
    11'b01111111001: data <= 32'hb571be6a;
    11'b01111111010: data <= 32'h39dabb6b;
    11'b01111111011: data <= 32'h3aba3d12;
    11'b01111111100: data <= 32'h362040c3;
    11'b01111111101: data <= 32'h38c73e25;
    11'b01111111110: data <= 32'h3d0f35f4;
    11'b01111111111: data <= 32'h3af932ad;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    