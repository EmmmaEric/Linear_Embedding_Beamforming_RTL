
module memory_rom_20(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3dcf391a;
    11'b00000000001: data <= 32'h3a6534e2;
    11'b00000000010: data <= 32'hbaf6b713;
    11'b00000000011: data <= 32'hbc9bbdeb;
    11'b00000000100: data <= 32'h38febe77;
    11'b00000000101: data <= 32'h4089b955;
    11'b00000000110: data <= 32'h3f3baa5a;
    11'b00000000111: data <= 32'h2b9fb87a;
    11'b00000001000: data <= 32'hbba9bbaf;
    11'b00000001001: data <= 32'hbb7aa5e5;
    11'b00000001010: data <= 32'hbc2b3ca4;
    11'b00000001011: data <= 32'hbe1f38d2;
    11'b00000001100: data <= 32'hbd91bd60;
    11'b00000001101: data <= 32'hb674c037;
    11'b00000001110: data <= 32'h3432b7b7;
    11'b00000001111: data <= 32'h0b853ea6;
    11'b00000010000: data <= 32'hb16a4032;
    11'b00000010001: data <= 32'h383c3cae;
    11'b00000010010: data <= 32'h3c07398b;
    11'b00000010011: data <= 32'h1ee63bfc;
    11'b00000010100: data <= 32'hbdc03a92;
    11'b00000010101: data <= 32'hbc51b381;
    11'b00000010110: data <= 32'h3ca8bbee;
    11'b00000010111: data <= 32'h4186b9e2;
    11'b00000011000: data <= 32'h4006b531;
    11'b00000011001: data <= 32'h3475b7ff;
    11'b00000011010: data <= 32'hb432b835;
    11'b00000011011: data <= 32'h344434d0;
    11'b00000011100: data <= 32'h300b3b2c;
    11'b00000011101: data <= 32'hbc1ab24c;
    11'b00000011110: data <= 32'hbebfc056;
    11'b00000011111: data <= 32'hbc1ec121;
    11'b00000100000: data <= 32'hae5db9d3;
    11'b00000100001: data <= 32'h2bb43c9c;
    11'b00000100010: data <= 32'had1b3ca1;
    11'b00000100011: data <= 32'h30f1336f;
    11'b00000100100: data <= 32'h2f49368e;
    11'b00000100101: data <= 32'hbb9d3e51;
    11'b00000100110: data <= 32'hbff23f46;
    11'b00000100111: data <= 32'hbce73815;
    11'b00000101000: data <= 32'h3bd9ba1a;
    11'b00000101001: data <= 32'h407ab998;
    11'b00000101010: data <= 32'h3daf276d;
    11'b00000101011: data <= 32'h33a834f3;
    11'b00000101100: data <= 32'h387135c4;
    11'b00000101101: data <= 32'h3e393a22;
    11'b00000101110: data <= 32'h3c9e3abb;
    11'b00000101111: data <= 32'hb92eb657;
    11'b00000110000: data <= 32'hbec7c03d;
    11'b00000110001: data <= 32'hbaf2c0b7;
    11'b00000110010: data <= 32'h3779bb2a;
    11'b00000110011: data <= 32'h39c83377;
    11'b00000110100: data <= 32'h31acb3e1;
    11'b00000110101: data <= 32'hb117bb5a;
    11'b00000110110: data <= 32'hb71f262d;
    11'b00000110111: data <= 32'hbd433f25;
    11'b00000111000: data <= 32'hc0354005;
    11'b00000111001: data <= 32'hbe083500;
    11'b00000111010: data <= 32'h2fecbc87;
    11'b00000111011: data <= 32'h3b84b9cf;
    11'b00000111100: data <= 32'h357f389b;
    11'b00000111101: data <= 32'ha6813c90;
    11'b00000111110: data <= 32'h3c303bf9;
    11'b00000111111: data <= 32'h405e3c35;
    11'b00001000000: data <= 32'h3d8f3c64;
    11'b00001000001: data <= 32'hb9ce33dc;
    11'b00001000010: data <= 32'hbe48bc70;
    11'b00001000011: data <= 32'hb2d2be20;
    11'b00001000100: data <= 32'h3db5baca;
    11'b00001000101: data <= 32'h3dddb861;
    11'b00001000110: data <= 32'h3744bd1b;
    11'b00001000111: data <= 32'hadafbe39;
    11'b00001001000: data <= 32'hb096b017;
    11'b00001001001: data <= 32'hb99b3e96;
    11'b00001001010: data <= 32'hbe773dc3;
    11'b00001001011: data <= 32'hbedab8aa;
    11'b00001001100: data <= 32'hbb13bf4e;
    11'b00001001101: data <= 32'hb5c0bae4;
    11'b00001001110: data <= 32'hb8723a78;
    11'b00001001111: data <= 32'hb4a23d08;
    11'b00001010000: data <= 32'h3c203a62;
    11'b00001010001: data <= 32'h3f8f3b0a;
    11'b00001010010: data <= 32'h3a0b3df9;
    11'b00001010011: data <= 32'hbcf23d76;
    11'b00001010100: data <= 32'hbe0a347a;
    11'b00001010101: data <= 32'h3565b889;
    11'b00001010110: data <= 32'h3fd6b90f;
    11'b00001010111: data <= 32'h3e8eba33;
    11'b00001011000: data <= 32'h37d6bd85;
    11'b00001011001: data <= 32'h3589bd42;
    11'b00001011010: data <= 32'h3b5e2f59;
    11'b00001011011: data <= 32'h38d13da0;
    11'b00001011100: data <= 32'hba263958;
    11'b00001011101: data <= 32'hbec9bdad;
    11'b00001011110: data <= 32'hbdc3c086;
    11'b00001011111: data <= 32'hbb27bbc1;
    11'b00001100000: data <= 32'hb9d53822;
    11'b00001100001: data <= 32'hb50d3710;
    11'b00001100010: data <= 32'h3973b42e;
    11'b00001100011: data <= 32'h3c393432;
    11'b00001100100: data <= 32'hb2043f00;
    11'b00001100101: data <= 32'hbf1a408c;
    11'b00001100110: data <= 32'hbe3f3cd1;
    11'b00001100111: data <= 32'h353fac3e;
    11'b00001101000: data <= 32'h3e30b709;
    11'b00001101001: data <= 32'h3b88b704;
    11'b00001101010: data <= 32'h305eb946;
    11'b00001101011: data <= 32'h3ab8b79b;
    11'b00001101100: data <= 32'h40383895;
    11'b00001101101: data <= 32'h3f423d2e;
    11'b00001101110: data <= 32'had533567;
    11'b00001101111: data <= 32'hbe04bddf;
    11'b00001110000: data <= 32'hbd20bfe5;
    11'b00001110001: data <= 32'hb713bad2;
    11'b00001110010: data <= 32'hb0d4ade0;
    11'b00001110011: data <= 32'hacc1badc;
    11'b00001110100: data <= 32'h3582be65;
    11'b00001110101: data <= 32'h3688b74d;
    11'b00001110110: data <= 32'hb9193edf;
    11'b00001110111: data <= 32'hbf5540e7;
    11'b00001111000: data <= 32'hbe653c94;
    11'b00001111001: data <= 32'hb3adb4f1;
    11'b00001111010: data <= 32'h35a6b6e0;
    11'b00001111011: data <= 32'hb51d2f17;
    11'b00001111100: data <= 32'hb7a73317;
    11'b00001111101: data <= 32'h3c40335e;
    11'b00001111110: data <= 32'h416a3a9c;
    11'b00001111111: data <= 32'h406b3d67;
    11'b00010000000: data <= 32'h219339be;
    11'b00010000001: data <= 32'hbd40b885;
    11'b00010000010: data <= 32'hb912bbc7;
    11'b00010000011: data <= 32'h383eb731;
    11'b00010000100: data <= 32'h3920b8a9;
    11'b00010000101: data <= 32'h3219bf64;
    11'b00010000110: data <= 32'h3428c0d5;
    11'b00010000111: data <= 32'h37b1ba9e;
    11'b00010001000: data <= 32'hb02a3de6;
    11'b00010001001: data <= 32'hbcc33f8f;
    11'b00010001010: data <= 32'hbdd2344d;
    11'b00010001011: data <= 32'hbb93bc18;
    11'b00010001100: data <= 32'hbb2eb883;
    11'b00010001101: data <= 32'hbdae374c;
    11'b00010001110: data <= 32'hbc063841;
    11'b00010001111: data <= 32'h3b3e307a;
    11'b00010010000: data <= 32'h40d73835;
    11'b00010010001: data <= 32'h3e823dad;
    11'b00010010010: data <= 32'hb7d03e24;
    11'b00010010011: data <= 32'hbd003a27;
    11'b00010010100: data <= 32'h9ce432ab;
    11'b00010010101: data <= 32'h3ce22c8e;
    11'b00010010110: data <= 32'h3b5bb90a;
    11'b00010010111: data <= 32'h3027bfd2;
    11'b00010011000: data <= 32'h3668c086;
    11'b00010011001: data <= 32'h3d00b917;
    11'b00010011010: data <= 32'h3c6f3ce4;
    11'b00010011011: data <= 32'hafd63c42;
    11'b00010011100: data <= 32'hbc68b98b;
    11'b00010011101: data <= 32'hbd27be40;
    11'b00010011110: data <= 32'hbdbcb8d8;
    11'b00010011111: data <= 32'hbee036b7;
    11'b00010100000: data <= 32'hbc879e5a;
    11'b00010100001: data <= 32'h3831bac7;
    11'b00010100010: data <= 32'h3e37b4e8;
    11'b00010100011: data <= 32'h38b63d4a;
    11'b00010100100: data <= 32'hbc7b4067;
    11'b00010100101: data <= 32'hbd0d3ec5;
    11'b00010100110: data <= 32'h327b3af8;
    11'b00010100111: data <= 32'h3c4536b0;
    11'b00010101000: data <= 32'h34dbb384;
    11'b00010101001: data <= 32'hb6c3bcde;
    11'b00010101010: data <= 32'h3850bd74;
    11'b00010101011: data <= 32'h405bae61;
    11'b00010101100: data <= 32'h40a13c5f;
    11'b00010101101: data <= 32'h3a0f386e;
    11'b00010101110: data <= 32'hb99dbbda;
    11'b00010101111: data <= 32'hbc25bd75;
    11'b00010110000: data <= 32'hbbceb502;
    11'b00010110001: data <= 32'hbc7b30fe;
    11'b00010110010: data <= 32'hbab4bc25;
    11'b00010110011: data <= 32'h31c7c059;
    11'b00010110100: data <= 32'h3a14bcfa;
    11'b00010110101: data <= 32'had153c24;
    11'b00010110110: data <= 32'hbd21407f;
    11'b00010110111: data <= 32'hbc9d3e89;
    11'b00010111000: data <= 32'ha8f7393a;
    11'b00010111001: data <= 32'h30a1369b;
    11'b00010111010: data <= 32'hbb8c3520;
    11'b00010111011: data <= 32'hbd17b30e;
    11'b00010111100: data <= 32'h377fb761;
    11'b00010111101: data <= 32'h413c344c;
    11'b00010111110: data <= 32'h41703c25;
    11'b00010111111: data <= 32'h3b603910;
    11'b00011000000: data <= 32'hb7a4b594;
    11'b00011000001: data <= 32'hb5f0b62f;
    11'b00011000010: data <= 32'h2d7f354e;
    11'b00011000011: data <= 32'hb11da334;
    11'b00011000100: data <= 32'hb742bf5f;
    11'b00011000101: data <= 32'h246dc205;
    11'b00011000110: data <= 32'h387cbeed;
    11'b00011000111: data <= 32'h311939a7;
    11'b00011001000: data <= 32'hb9703e9b;
    11'b00011001001: data <= 32'hba303987;
    11'b00011001010: data <= 32'hb689b250;
    11'b00011001011: data <= 32'hbb3b3150;
    11'b00011001100: data <= 32'hc02439bc;
    11'b00011001101: data <= 32'hbfd83548;
    11'b00011001110: data <= 32'h3189b49a;
    11'b00011001111: data <= 32'h408a27a9;
    11'b00011010000: data <= 32'h402e3b18;
    11'b00011010001: data <= 32'h35363c6d;
    11'b00011010010: data <= 32'hb8143a23;
    11'b00011010011: data <= 32'h34ad3a9d;
    11'b00011010100: data <= 32'h3be43c35;
    11'b00011010101: data <= 32'h35fe3011;
    11'b00011010110: data <= 32'hb6e3bf78;
    11'b00011010111: data <= 32'ha817c1a9;
    11'b00011011000: data <= 32'h3bf3bdf3;
    11'b00011011001: data <= 32'h3cab3829;
    11'b00011011010: data <= 32'h36b93a63;
    11'b00011011011: data <= 32'hb212b745;
    11'b00011011100: data <= 32'hb81fbbd6;
    11'b00011011101: data <= 32'hbd57256a;
    11'b00011011110: data <= 32'hc0bb3ab5;
    11'b00011011111: data <= 32'hc02b2f59;
    11'b00011100000: data <= 32'hb1c3bc21;
    11'b00011100001: data <= 32'h3d80ba97;
    11'b00011100010: data <= 32'h3b243857;
    11'b00011100011: data <= 32'hb8473e01;
    11'b00011100100: data <= 32'hb91b3e42;
    11'b00011100101: data <= 32'h39043e0b;
    11'b00011100110: data <= 32'h3c8d3dd0;
    11'b00011100111: data <= 32'h20bb3852;
    11'b00011101000: data <= 32'hbbe4bc61;
    11'b00011101001: data <= 32'hb090bf31;
    11'b00011101010: data <= 32'h3e7fb9f7;
    11'b00011101011: data <= 32'h40743819;
    11'b00011101100: data <= 32'h3d5d31f4;
    11'b00011101101: data <= 32'h351ebc1f;
    11'b00011101110: data <= 32'hb236bc29;
    11'b00011101111: data <= 32'hbaaa34b7;
    11'b00011110000: data <= 32'hbea93a85;
    11'b00011110001: data <= 32'hbe79b8d5;
    11'b00011110010: data <= 32'hb681c065;
    11'b00011110011: data <= 32'h3801bf43;
    11'b00011110100: data <= 32'ha9e02e35;
    11'b00011110101: data <= 32'hbbb53db7;
    11'b00011110110: data <= 32'hb8973dcc;
    11'b00011110111: data <= 32'h38df3ce3;
    11'b00011111000: data <= 32'h38433d48;
    11'b00011111001: data <= 32'hbc3e3bf6;
    11'b00011111010: data <= 32'hbf96a843;
    11'b00011111011: data <= 32'hb68fb927;
    11'b00011111100: data <= 32'h3f96aeb6;
    11'b00011111101: data <= 32'h41203837;
    11'b00011111110: data <= 32'h3ddf2c0e;
    11'b00011111111: data <= 32'h3782b9be;
    11'b00100000000: data <= 32'h3668b417;
    11'b00100000001: data <= 32'h348f3bfc;
    11'b00100000010: data <= 32'hb79e3af3;
    11'b00100000011: data <= 32'hbbb6bcd3;
    11'b00100000100: data <= 32'hb795c1e7;
    11'b00100000101: data <= 32'h2ff6c098;
    11'b00100000110: data <= 32'hb016b2db;
    11'b00100000111: data <= 32'hb8963ae6;
    11'b00100001000: data <= 32'hb0b13741;
    11'b00100001001: data <= 32'h37ab3175;
    11'b00100001010: data <= 32'hb4813a89;
    11'b00100001011: data <= 32'hc0323d1f;
    11'b00100001100: data <= 32'hc139395b;
    11'b00100001101: data <= 32'hb9f6b0e6;
    11'b00100001110: data <= 32'h3e26aee5;
    11'b00100001111: data <= 32'h3f8435a0;
    11'b00100010000: data <= 32'h399f34ad;
    11'b00100010001: data <= 32'h32a33076;
    11'b00100010010: data <= 32'h3b983ad9;
    11'b00100010011: data <= 32'h3d443f18;
    11'b00100010100: data <= 32'h35ea3c69;
    11'b00100010101: data <= 32'hb977bcb5;
    11'b00100010110: data <= 32'hb829c170;
    11'b00100010111: data <= 32'h3513bfaf;
    11'b00100011000: data <= 32'h38ceb2ab;
    11'b00100011001: data <= 32'h368a2f56;
    11'b00100011010: data <= 32'h3817ba77;
    11'b00100011011: data <= 32'h381dbb4e;
    11'b00100011100: data <= 32'hb8f43660;
    11'b00100011101: data <= 32'hc0ae3d79;
    11'b00100011110: data <= 32'hc1493973;
    11'b00100011111: data <= 32'hbb9db8d1;
    11'b00100100000: data <= 32'h39d6ba93;
    11'b00100100001: data <= 32'h389bacad;
    11'b00100100010: data <= 32'hb722380b;
    11'b00100100011: data <= 32'hb27f3a73;
    11'b00100100100: data <= 32'h3ce63df5;
    11'b00100100101: data <= 32'h3eb74040;
    11'b00100100110: data <= 32'h34ff3db1;
    11'b00100100111: data <= 32'hbc4bb77a;
    11'b00100101000: data <= 32'hb9a4be5c;
    11'b00100101001: data <= 32'h39ecbb47;
    11'b00100101010: data <= 32'h3dfd2c28;
    11'b00100101011: data <= 32'h3d1db6b9;
    11'b00100101100: data <= 32'h3c11be52;
    11'b00100101101: data <= 32'h3a66bd2b;
    11'b00100101110: data <= 32'hb0d237a6;
    11'b00100101111: data <= 32'hbe383d9c;
    11'b00100110000: data <= 32'hbfbe31e6;
    11'b00100110001: data <= 32'hbb45be4c;
    11'b00100110010: data <= 32'hab4cbf08;
    11'b00100110011: data <= 32'hb862b86c;
    11'b00100110100: data <= 32'hbcd03694;
    11'b00100110101: data <= 32'hb5c73988;
    11'b00100110110: data <= 32'h3cf83c86;
    11'b00100110111: data <= 32'h3d363f2a;
    11'b00100111000: data <= 32'hb84d3e89;
    11'b00100111001: data <= 32'hbfaa3807;
    11'b00100111010: data <= 32'hbc22b434;
    11'b00100111011: data <= 32'h3b832c3f;
    11'b00100111100: data <= 32'h3f313548;
    11'b00100111101: data <= 32'h3d66b86f;
    11'b00100111110: data <= 32'h3c0cbdff;
    11'b00100111111: data <= 32'h3cc2ba04;
    11'b00101000000: data <= 32'h3b0f3c62;
    11'b00101000001: data <= 32'hb29a3e22;
    11'b00101000010: data <= 32'hbb93b4d5;
    11'b00101000011: data <= 32'hb9a0c087;
    11'b00101000100: data <= 32'hb6b8c064;
    11'b00101000101: data <= 32'hbae3ba11;
    11'b00101000110: data <= 32'hbc56120a;
    11'b00101000111: data <= 32'ha988b37a;
    11'b00101001000: data <= 32'h3cc8ac27;
    11'b00101001001: data <= 32'h39183bba;
    11'b00101001010: data <= 32'hbdee3e89;
    11'b00101001011: data <= 32'hc1323caf;
    11'b00101001100: data <= 32'hbd3f3756;
    11'b00101001101: data <= 32'h397935cc;
    11'b00101001110: data <= 32'h3caa34bc;
    11'b00101001111: data <= 32'h374eb675;
    11'b00101010000: data <= 32'h3737ba89;
    11'b00101010001: data <= 32'h3dd233b6;
    11'b00101010010: data <= 32'h3f743f61;
    11'b00101010011: data <= 32'h3aed3f05;
    11'b00101010100: data <= 32'hb577b53a;
    11'b00101010101: data <= 32'hb893c01f;
    11'b00101010110: data <= 32'hb4acbed7;
    11'b00101010111: data <= 32'hb545b7cf;
    11'b00101011000: data <= 32'hb400b7af;
    11'b00101011001: data <= 32'h38b2bdc0;
    11'b00101011010: data <= 32'h3d05bd7a;
    11'b00101011011: data <= 32'h34ae3286;
    11'b00101011100: data <= 32'hbef53e09;
    11'b00101011101: data <= 32'hc1163ce9;
    11'b00101011110: data <= 32'hbd2e3322;
    11'b00101011111: data <= 32'h2f6cb16f;
    11'b00101100000: data <= 32'had12adc2;
    11'b00101100001: data <= 32'hbb3db3cc;
    11'b00101100010: data <= 32'hb501b206;
    11'b00101100011: data <= 32'h3df53af5;
    11'b00101100100: data <= 32'h40804046;
    11'b00101100101: data <= 32'h3c233f99;
    11'b00101100110: data <= 32'hb81b31b0;
    11'b00101100111: data <= 32'hb98ebbe4;
    11'b00101101000: data <= 32'h2be1b7f3;
    11'b00101101001: data <= 32'h37d43074;
    11'b00101101010: data <= 32'h38c1ba08;
    11'b00101101011: data <= 32'h3c3bc070;
    11'b00101101100: data <= 32'h3dadbff1;
    11'b00101101101: data <= 32'h38c4272c;
    11'b00101101110: data <= 32'hbc023dcc;
    11'b00101101111: data <= 32'hbe9b3a71;
    11'b00101110000: data <= 32'hbb45b918;
    11'b00101110001: data <= 32'hb66cbc38;
    11'b00101110010: data <= 32'hbcceb86a;
    11'b00101110011: data <= 32'hbfa4b445;
    11'b00101110100: data <= 32'hba18b1c4;
    11'b00101110101: data <= 32'h3d843871;
    11'b00101110110: data <= 32'h3fc73e94;
    11'b00101110111: data <= 32'h35343f2b;
    11'b00101111000: data <= 32'hbd1b3b0c;
    11'b00101111001: data <= 32'hbc0c354d;
    11'b00101111010: data <= 32'h349b39e3;
    11'b00101111011: data <= 32'h3af439d3;
    11'b00101111100: data <= 32'h39a1b9ce;
    11'b00101111101: data <= 32'h3b69c067;
    11'b00101111110: data <= 32'h3e1bbe74;
    11'b00101111111: data <= 32'h3d7e3845;
    11'b00110000000: data <= 32'h35493e42;
    11'b00110000001: data <= 32'hb6713530;
    11'b00110000010: data <= 32'hb5a8bd76;
    11'b00110000011: data <= 32'hb88fbe18;
    11'b00110000100: data <= 32'hbe49b952;
    11'b00110000101: data <= 32'hbff2b70d;
    11'b00110000110: data <= 32'hb8c2bafc;
    11'b00110000111: data <= 32'h3d36b8f4;
    11'b00110001000: data <= 32'h3d3b3888;
    11'b00110001001: data <= 32'hb8f93db5;
    11'b00110001010: data <= 32'hbfe93d4f;
    11'b00110001011: data <= 32'hbce93c69;
    11'b00110001100: data <= 32'h330e3d06;
    11'b00110001101: data <= 32'h370a3b1c;
    11'b00110001110: data <= 32'hb139b832;
    11'b00110001111: data <= 32'h302abe42;
    11'b00110010000: data <= 32'h3db5b937;
    11'b00110010001: data <= 32'h403b3d27;
    11'b00110010010: data <= 32'h3dc73f00;
    11'b00110010011: data <= 32'h37403117;
    11'b00110010100: data <= 32'h251bbd56;
    11'b00110010101: data <= 32'hb5ccbc46;
    11'b00110010110: data <= 32'hbc62b1e6;
    11'b00110010111: data <= 32'hbce1b894;
    11'b00110011000: data <= 32'h2572bf54;
    11'b00110011001: data <= 32'h3d61bfd6;
    11'b00110011010: data <= 32'h3aedb775;
    11'b00110011011: data <= 32'hbc143c10;
    11'b00110011100: data <= 32'hbfd73d16;
    11'b00110011101: data <= 32'hbc213b72;
    11'b00110011110: data <= 32'ha65f3aa4;
    11'b00110011111: data <= 32'hb8843860;
    11'b00110100000: data <= 32'hbe39b5b2;
    11'b00110100001: data <= 32'hbb55bb01;
    11'b00110100010: data <= 32'h3c8e2dba;
    11'b00110100011: data <= 32'h40b73e80;
    11'b00110100100: data <= 32'h3eba3f02;
    11'b00110100101: data <= 32'h36d935fe;
    11'b00110100110: data <= 32'ha4b2b7d6;
    11'b00110100111: data <= 32'h1aee316f;
    11'b00110101000: data <= 32'hb40039d4;
    11'b00110101001: data <= 32'hb4b5b802;
    11'b00110101010: data <= 32'h3853c0e2;
    11'b00110101011: data <= 32'h3d9dc14b;
    11'b00110101100: data <= 32'h3b58ba9f;
    11'b00110101101: data <= 32'hb8023a99;
    11'b00110101110: data <= 32'hbc353a92;
    11'b00110101111: data <= 32'hb5e22c6f;
    11'b00110110000: data <= 32'hb1f0ae85;
    11'b00110110001: data <= 32'hbdfd2911;
    11'b00110110010: data <= 32'hc145b4f2;
    11'b00110110011: data <= 32'hbe5bb945;
    11'b00110110100: data <= 32'h3ac9a55b;
    11'b00110110101: data <= 32'h40013c86;
    11'b00110110110: data <= 32'h3bed3d88;
    11'b00110110111: data <= 32'hb58139c4;
    11'b00110111000: data <= 32'hb5e03904;
    11'b00110111001: data <= 32'h345e3dec;
    11'b00110111010: data <= 32'h34c23e4d;
    11'b00110111011: data <= 32'h18b4b3db;
    11'b00110111100: data <= 32'h36d6c0b3;
    11'b00110111101: data <= 32'h3d1ec09e;
    11'b00110111110: data <= 32'h3d67b5aa;
    11'b00110111111: data <= 32'h38fe3b93;
    11'b00111000000: data <= 32'h346834fd;
    11'b00111000001: data <= 32'h3792ba4f;
    11'b00111000010: data <= 32'had66b9e7;
    11'b00111000011: data <= 32'hbf14af11;
    11'b00111000100: data <= 32'hc187b4a1;
    11'b00111000101: data <= 32'hbdfebc1d;
    11'b00111000110: data <= 32'h39f8bbe0;
    11'b00111000111: data <= 32'h3d5da513;
    11'b00111001000: data <= 32'hab0139bb;
    11'b00111001001: data <= 32'hbcc33ae6;
    11'b00111001010: data <= 32'hb9123d1f;
    11'b00111001011: data <= 32'h35c54026;
    11'b00111001100: data <= 32'h312f3f71;
    11'b00111001101: data <= 32'hb93b25d1;
    11'b00111001110: data <= 32'hb6dabebe;
    11'b00111001111: data <= 32'h3b02bd1d;
    11'b00111010000: data <= 32'h3f0e3829;
    11'b00111010001: data <= 32'h3e693cc2;
    11'b00111010010: data <= 32'h3ce426ce;
    11'b00111010011: data <= 32'h3c17bc14;
    11'b00111010100: data <= 32'h3396b7da;
    11'b00111010101: data <= 32'hbd0a3692;
    11'b00111010110: data <= 32'hbfd4b01a;
    11'b00111010111: data <= 32'hba5abe97;
    11'b00111011000: data <= 32'h3ac0c059;
    11'b00111011001: data <= 32'h3a75bca1;
    11'b00111011010: data <= 32'hb97a2d2a;
    11'b00111011011: data <= 32'hbd823924;
    11'b00111011100: data <= 32'hb6b93c3f;
    11'b00111011101: data <= 32'h362b3e8d;
    11'b00111011110: data <= 32'hb8073de2;
    11'b00111011111: data <= 32'hbf8a30ba;
    11'b00111100000: data <= 32'hbe58bb6d;
    11'b00111100001: data <= 32'h3535b554;
    11'b00111100010: data <= 32'h3f2f3c3a;
    11'b00111100011: data <= 32'h3f1c3cca;
    11'b00111100100: data <= 32'h3ce00677;
    11'b00111100101: data <= 32'h3be4b80b;
    11'b00111100110: data <= 32'h38aa38a0;
    11'b00111100111: data <= 32'hb5c33dbd;
    11'b00111101000: data <= 32'hbada336c;
    11'b00111101001: data <= 32'had30c004;
    11'b00111101010: data <= 32'h3b75c191;
    11'b00111101011: data <= 32'h3933be49;
    11'b00111101100: data <= 32'hb7bcb15a;
    11'b00111101101: data <= 32'hb92d31a6;
    11'b00111101110: data <= 32'h359430f1;
    11'b00111101111: data <= 32'h38383880;
    11'b00111110000: data <= 32'hbca33a48;
    11'b00111110001: data <= 32'hc1c130a4;
    11'b00111110010: data <= 32'hc0aeb846;
    11'b00111110011: data <= 32'had09b085;
    11'b00111110100: data <= 32'h3d853a06;
    11'b00111110101: data <= 32'h3c2a39ed;
    11'b00111110110: data <= 32'h35652941;
    11'b00111110111: data <= 32'h37c2350d;
    11'b00111111000: data <= 32'h3a5a3f2d;
    11'b00111111001: data <= 32'h355440c6;
    11'b00111111010: data <= 32'hb469393a;
    11'b00111111011: data <= 32'h200ebf41;
    11'b00111111100: data <= 32'h39f8c0cd;
    11'b00111111101: data <= 32'h3a49bc18;
    11'b00111111110: data <= 32'h35572c8f;
    11'b00111111111: data <= 32'h389bb473;
    11'b01000000000: data <= 32'h3d44ba97;
    11'b01000000001: data <= 32'h3abdb563;
    11'b01000000010: data <= 32'hbd2836c3;
    11'b01000000011: data <= 32'hc1ea324c;
    11'b01000000100: data <= 32'hc06db903;
    11'b01000000101: data <= 32'haf07ba51;
    11'b01000000110: data <= 32'h3a10b47c;
    11'b01000000111: data <= 32'haec9ac25;
    11'b01000001000: data <= 32'hb9ffac78;
    11'b01000001001: data <= 32'h18633a50;
    11'b01000001010: data <= 32'h3b1340ad;
    11'b01000001011: data <= 32'h3732415c;
    11'b01000001100: data <= 32'hb8eb3b38;
    11'b01000001101: data <= 32'hb9b2bca8;
    11'b01000001110: data <= 32'h3291bd1e;
    11'b01000001111: data <= 32'h3b592c40;
    11'b01000010000: data <= 32'h3c663833;
    11'b01000010001: data <= 32'h3de6b858;
    11'b01000010010: data <= 32'h3faabd20;
    11'b01000010011: data <= 32'h3cceb678;
    11'b01000010100: data <= 32'hba1c3a4e;
    11'b01000010101: data <= 32'hc02437b4;
    11'b01000010110: data <= 32'hbd4abb9c;
    11'b01000010111: data <= 32'h31efbef6;
    11'b01000011000: data <= 32'h3428bd78;
    11'b01000011001: data <= 32'hbb81ba52;
    11'b01000011010: data <= 32'hbcfdb62c;
    11'b01000011011: data <= 32'h290a382b;
    11'b01000011100: data <= 32'h3c0a3f58;
    11'b01000011101: data <= 32'h2d124048;
    11'b01000011110: data <= 32'hbe583ad5;
    11'b01000011111: data <= 32'hbf40b728;
    11'b01000100000: data <= 32'hb776b0df;
    11'b01000100001: data <= 32'h3a653b45;
    11'b01000100010: data <= 32'h3cc339d5;
    11'b01000100011: data <= 32'h3dacb928;
    11'b01000100100: data <= 32'h3f1bbc38;
    11'b01000100101: data <= 32'h3da5363e;
    11'b01000100110: data <= 32'h2e433efa;
    11'b01000100111: data <= 32'hba763bdb;
    11'b01000101000: data <= 32'hb501bc76;
    11'b01000101001: data <= 32'h37ccc077;
    11'b01000101010: data <= 32'h2aeebef6;
    11'b01000101011: data <= 32'hbc0fbbe3;
    11'b01000101100: data <= 32'hba71ba1d;
    11'b01000101101: data <= 32'h39cab5c1;
    11'b01000101110: data <= 32'h3d3438ee;
    11'b01000101111: data <= 32'hb58b3cb2;
    11'b01000110000: data <= 32'hc0dd3906;
    11'b01000110001: data <= 32'hc111a7f3;
    11'b01000110010: data <= 32'hbaf434e3;
    11'b01000110011: data <= 32'h36a93b41;
    11'b01000110100: data <= 32'h37603611;
    11'b01000110101: data <= 32'h3695b9ff;
    11'b01000110110: data <= 32'h3c15b7ca;
    11'b01000110111: data <= 32'h3d993dbc;
    11'b01000111000: data <= 32'h3a574159;
    11'b01000111001: data <= 32'h269a3dcc;
    11'b01000111010: data <= 32'h2de6bb2e;
    11'b01000111011: data <= 32'h36f8bf52;
    11'b01000111100: data <= 32'h2b2cbc59;
    11'b01000111101: data <= 32'hb779b83c;
    11'b01000111110: data <= 32'h332ebc0c;
    11'b01000111111: data <= 32'h3eb1bd4e;
    11'b01001000000: data <= 32'h3eceb829;
    11'b01001000001: data <= 32'hb66737c6;
    11'b01001000010: data <= 32'hc0f1381d;
    11'b01001000011: data <= 32'hc0a6a0c4;
    11'b01001000100: data <= 32'hb9cfac12;
    11'b01001000101: data <= 32'ha7362dcd;
    11'b01001000110: data <= 32'hb95fb677;
    11'b01001000111: data <= 32'hbb2dbbd6;
    11'b01001001000: data <= 32'h32afb056;
    11'b01001001001: data <= 32'h3d303faa;
    11'b01001001010: data <= 32'h3bfc41cf;
    11'b01001001011: data <= 32'ha7c13e4b;
    11'b01001001100: data <= 32'hb626b632;
    11'b01001001101: data <= 32'hac67b9c2;
    11'b01001001110: data <= 32'h2a2f32a6;
    11'b01001001111: data <= 32'h305e33ea;
    11'b01001010000: data <= 32'h3c2abc44;
    11'b01001010001: data <= 32'h4079bf65;
    11'b01001010010: data <= 32'h3ff6baf8;
    11'b01001010011: data <= 32'h279338a6;
    11'b01001010100: data <= 32'hbe5939e8;
    11'b01001010101: data <= 32'hbcfdb1f0;
    11'b01001010110: data <= 32'hafe7ba8a;
    11'b01001010111: data <= 32'hb4f2bb24;
    11'b01001011000: data <= 32'hbe34bc76;
    11'b01001011001: data <= 32'hbeb3bd1f;
    11'b01001011010: data <= 32'haa3ab5b0;
    11'b01001011011: data <= 32'h3d553da1;
    11'b01001011100: data <= 32'h3a2d4069;
    11'b01001011101: data <= 32'hba3b3cfa;
    11'b01001011110: data <= 32'hbd6e2f6a;
    11'b01001011111: data <= 32'hb9ec3716;
    11'b01001100000: data <= 32'haed33d51;
    11'b01001100001: data <= 32'h333b3a25;
    11'b01001100010: data <= 32'h3bc0bc2f;
    11'b01001100011: data <= 32'h3fdebf06;
    11'b01001100100: data <= 32'h3fd4b51a;
    11'b01001100101: data <= 32'h39893d88;
    11'b01001100110: data <= 32'hb4b73cf7;
    11'b01001100111: data <= 32'h28d4b461;
    11'b01001101000: data <= 32'h381abd0c;
    11'b01001101001: data <= 32'hb5d2bcf5;
    11'b01001101010: data <= 32'hbefdbcde;
    11'b01001101011: data <= 32'hbdf8bddc;
    11'b01001101100: data <= 32'h373dbc3f;
    11'b01001101101: data <= 32'h3e79314d;
    11'b01001101110: data <= 32'h37383bc7;
    11'b01001101111: data <= 32'hbe243962;
    11'b01001110000: data <= 32'hc01535b3;
    11'b01001110001: data <= 32'hbc543c08;
    11'b01001110010: data <= 32'hb59d3e69;
    11'b01001110011: data <= 32'hb5d03912;
    11'b01001110100: data <= 32'hab2dbc85;
    11'b01001110101: data <= 32'h3bb6bd3d;
    11'b01001110110: data <= 32'h3e6a38d2;
    11'b01001110111: data <= 32'h3cc54086;
    11'b01001111000: data <= 32'h39113eb6;
    11'b01001111001: data <= 32'h39e0b070;
    11'b01001111010: data <= 32'h39b4bbb1;
    11'b01001111011: data <= 32'hb514b890;
    11'b01001111100: data <= 32'hbd54b853;
    11'b01001111101: data <= 32'hb8eebd8d;
    11'b01001111110: data <= 32'h3d57bf50;
    11'b01001111111: data <= 32'h4006bc38;
    11'b01010000000: data <= 32'h35d3a545;
    11'b01010000001: data <= 32'hbe8c3458;
    11'b01010000010: data <= 32'hbf4334dc;
    11'b01010000011: data <= 32'hba083a34;
    11'b01010000100: data <= 32'hb8033bc4;
    11'b01010000101: data <= 32'hbd33abd7;
    11'b01010000110: data <= 32'hbdc1bd79;
    11'b01010000111: data <= 32'hb10dbbc2;
    11'b01010001000: data <= 32'h3cba3c71;
    11'b01010001001: data <= 32'h3d2b40f5;
    11'b01010001010: data <= 32'h39b53e9f;
    11'b01010001011: data <= 32'h37942f97;
    11'b01010001100: data <= 32'h353aa7f4;
    11'b01010001101: data <= 32'hb5663a56;
    11'b01010001110: data <= 32'hba373859;
    11'b01010001111: data <= 32'h3226bc69;
    11'b01010010000: data <= 32'h3f8ec06e;
    11'b01010010001: data <= 32'h4063be26;
    11'b01010010010: data <= 32'h38b3b180;
    11'b01010010011: data <= 32'hbb4c356c;
    11'b01010010100: data <= 32'hb96d303b;
    11'b01010010101: data <= 32'h30ab2e5f;
    11'b01010010110: data <= 32'hb6f827ad;
    11'b01010010111: data <= 32'hc00dba1a;
    11'b01010011000: data <= 32'hc0b1be68;
    11'b01010011001: data <= 32'hb986bc21;
    11'b01010011010: data <= 32'h3c1339e8;
    11'b01010011011: data <= 32'h3c353eeb;
    11'b01010011100: data <= 32'h2c1f3c31;
    11'b01010011101: data <= 32'hb6bc3478;
    11'b01010011110: data <= 32'hb53b3bbe;
    11'b01010011111: data <= 32'hb75b4014;
    11'b01010100000: data <= 32'hb8a33d75;
    11'b01010100001: data <= 32'h336fbabc;
    11'b01010100010: data <= 32'h3e55c02b;
    11'b01010100011: data <= 32'h3fa7bc65;
    11'b01010100100: data <= 32'h3b64381e;
    11'b01010100101: data <= 32'h32ce3a73;
    11'b01010100110: data <= 32'h39da288e;
    11'b01010100111: data <= 32'h3c69b680;
    11'b01010101000: data <= 32'hb2cfb674;
    11'b01010101001: data <= 32'hc051bac2;
    11'b01010101010: data <= 32'hc093be51;
    11'b01010101011: data <= 32'hb578bdc3;
    11'b01010101100: data <= 32'h3cf7b56b;
    11'b01010101101: data <= 32'h39e03607;
    11'b01010101110: data <= 32'hb9b43096;
    11'b01010101111: data <= 32'hbca732c5;
    11'b01010110000: data <= 32'hb9513dca;
    11'b01010110001: data <= 32'hb85640e6;
    11'b01010110010: data <= 32'hbb443db0;
    11'b01010110011: data <= 32'hb912baa1;
    11'b01010110100: data <= 32'h378abe93;
    11'b01010110101: data <= 32'h3ce5b211;
    11'b01010110110: data <= 32'h3c613db1;
    11'b01010110111: data <= 32'h3c273cfd;
    11'b01010111000: data <= 32'h3e4e2ac1;
    11'b01010111001: data <= 32'h3e25b52b;
    11'b01010111010: data <= 32'ha7752f8a;
    11'b01010111011: data <= 32'hbef7aceb;
    11'b01010111100: data <= 32'hbdcdbcb9;
    11'b01010111101: data <= 32'h3852bf79;
    11'b01010111110: data <= 32'h3e90bdc4;
    11'b01010111111: data <= 32'h388aba32;
    11'b01011000000: data <= 32'hbbebb843;
    11'b01011000001: data <= 32'hbc4ba59a;
    11'b01011000010: data <= 32'hb43d3cce;
    11'b01011000011: data <= 32'hb65f3f89;
    11'b01011000100: data <= 32'hbe0d3a19;
    11'b01011000101: data <= 32'hbf8fbc43;
    11'b01011000110: data <= 32'hba83bd02;
    11'b01011000111: data <= 32'h37e33747;
    11'b01011001000: data <= 32'h3bc23f0e;
    11'b01011001001: data <= 32'h3c5c3cb3;
    11'b01011001010: data <= 32'h3da32a65;
    11'b01011001011: data <= 32'h3ce934aa;
    11'b01011001100: data <= 32'ha81f3d65;
    11'b01011001101: data <= 32'hbca13cae;
    11'b01011001110: data <= 32'hb855b87e;
    11'b01011001111: data <= 32'h3cd0bff9;
    11'b01011010000: data <= 32'h3f2fbf85;
    11'b01011010001: data <= 32'h388ebc2e;
    11'b01011010010: data <= 32'hb873b8bb;
    11'b01011010011: data <= 32'hac63b3a5;
    11'b01011010100: data <= 32'h3a523816;
    11'b01011010101: data <= 32'h226e3b05;
    11'b01011010110: data <= 32'hbfcba833;
    11'b01011010111: data <= 32'hc179bd2e;
    11'b01011011000: data <= 32'hbdf6bc8a;
    11'b01011011001: data <= 32'h30df358b;
    11'b01011011010: data <= 32'h392b3c96;
    11'b01011011011: data <= 32'h36e336d6;
    11'b01011011100: data <= 32'h37beb03a;
    11'b01011011101: data <= 32'h38083be0;
    11'b01011011110: data <= 32'hb14b410e;
    11'b01011011111: data <= 32'hba90404f;
    11'b01011100000: data <= 32'hb441acc5;
    11'b01011100001: data <= 32'h3c23bef1;
    11'b01011100010: data <= 32'h3d96bdb7;
    11'b01011100011: data <= 32'h389cb5d2;
    11'b01011100100: data <= 32'h341dad99;
    11'b01011100101: data <= 32'h3d10b521;
    11'b01011100110: data <= 32'h3fb7ae5a;
    11'b01011100111: data <= 32'h380b33a4;
    11'b01011101000: data <= 32'hbfa8b413;
    11'b01011101001: data <= 32'hc153bcbb;
    11'b01011101010: data <= 32'hbcbabcf3;
    11'b01011101011: data <= 32'h35e9b6bb;
    11'b01011101100: data <= 32'h3557afe6;
    11'b01011101101: data <= 32'hb6c7b95f;
    11'b01011101110: data <= 32'hb6eab80b;
    11'b01011101111: data <= 32'h26b53d0c;
    11'b01011110000: data <= 32'hb21441d5;
    11'b01011110001: data <= 32'hbb024094;
    11'b01011110010: data <= 32'hbaa4a01a;
    11'b01011110011: data <= 32'h234dbd1d;
    11'b01011110100: data <= 32'h3819b763;
    11'b01011110101: data <= 32'h36a8397d;
    11'b01011110110: data <= 32'h3acc37c8;
    11'b01011110111: data <= 32'h402db553;
    11'b01011111000: data <= 32'h40f4b407;
    11'b01011111001: data <= 32'h3a5b378b;
    11'b01011111010: data <= 32'hbdd0368a;
    11'b01011111011: data <= 32'hbf1fb8cc;
    11'b01011111100: data <= 32'hb21bbd48;
    11'b01011111101: data <= 32'h3b19bd11;
    11'b01011111110: data <= 32'h310bbd01;
    11'b01011111111: data <= 32'hbb33bdfe;
    11'b01100000000: data <= 32'hb8e8bb31;
    11'b01100000001: data <= 32'h34ec3b85;
    11'b01100000010: data <= 32'h2f7640a2;
    11'b01100000011: data <= 32'hbc8d3e39;
    11'b01100000100: data <= 32'hbf40b573;
    11'b01100000101: data <= 32'hbcf9bb1e;
    11'b01100000110: data <= 32'hb66d359e;
    11'b01100000111: data <= 32'h2cf33d1f;
    11'b01100001000: data <= 32'h3a55385d;
    11'b01100001001: data <= 32'h3f97b783;
    11'b01100001010: data <= 32'h4045288b;
    11'b01100001011: data <= 32'h39d53daf;
    11'b01100001100: data <= 32'hbafc3e7b;
    11'b01100001101: data <= 32'hb9d53326;
    11'b01100001110: data <= 32'h39a9bcbe;
    11'b01100001111: data <= 32'h3cbdbe3e;
    11'b01100010000: data <= 32'h2b3cbe0a;
    11'b01100010001: data <= 32'hba2ebe4b;
    11'b01100010010: data <= 32'h2eeabc64;
    11'b01100010011: data <= 32'h3d4433df;
    11'b01100010100: data <= 32'h39ec3cc4;
    11'b01100010101: data <= 32'hbd1e385f;
    11'b01100010110: data <= 32'hc0f8b9c2;
    11'b01100010111: data <= 32'hbfaab997;
    11'b01100011000: data <= 32'hba783832;
    11'b01100011001: data <= 32'hb47f3b93;
    11'b01100011010: data <= 32'h2f2eb091;
    11'b01100011011: data <= 32'h3b04bae6;
    11'b01100011100: data <= 32'h3ce8369e;
    11'b01100011101: data <= 32'h372340cd;
    11'b01100011110: data <= 32'hb7d14138;
    11'b01100011111: data <= 32'hb2453a97;
    11'b01100100000: data <= 32'h3a95bab1;
    11'b01100100001: data <= 32'h3aebbc44;
    11'b01100100010: data <= 32'hb055ba07;
    11'b01100100011: data <= 32'hb489bb5c;
    11'b01100100100: data <= 32'h3ce8bc2b;
    11'b01100100101: data <= 32'h40edb642;
    11'b01100100110: data <= 32'h3d8c3522;
    11'b01100100111: data <= 32'hbc66293f;
    11'b01100101000: data <= 32'hc0aeb9ad;
    11'b01100101001: data <= 32'hbe36b8fd;
    11'b01100101010: data <= 32'hb7c92d60;
    11'b01100101011: data <= 32'hb7b9adf7;
    11'b01100101100: data <= 32'hba11bd00;
    11'b01100101101: data <= 32'hb3ddbdb1;
    11'b01100101110: data <= 32'h378437f6;
    11'b01100101111: data <= 32'h34b84164;
    11'b01100110000: data <= 32'hb64f416b;
    11'b01100110001: data <= 32'hb7063aae;
    11'b01100110010: data <= 32'h2a1ab73e;
    11'b01100110011: data <= 32'ha5dcad48;
    11'b01100110100: data <= 32'hb80c37a9;
    11'b01100110101: data <= 32'h2cdcad1a;
    11'b01100110110: data <= 32'h3fbcbb46;
    11'b01100110111: data <= 32'h4200b94d;
    11'b01100111000: data <= 32'h3eb233c7;
    11'b01100111001: data <= 32'hb955371a;
    11'b01100111010: data <= 32'hbdbdb077;
    11'b01100111011: data <= 32'hb674b7c6;
    11'b01100111100: data <= 32'h3471b7f5;
    11'b01100111101: data <= 32'hb80bbc59;
    11'b01100111110: data <= 32'hbd4ec02e;
    11'b01100111111: data <= 32'hb9c8bf7a;
    11'b01101000000: data <= 32'h37a030f3;
    11'b01101000001: data <= 32'h3884401f;
    11'b01101000010: data <= 32'hb7053f5e;
    11'b01101000011: data <= 32'hbc89348d;
    11'b01101000100: data <= 32'hbc3ab2d5;
    11'b01101000101: data <= 32'hbbbb3a6b;
    11'b01101000110: data <= 32'hbb9a3d69;
    11'b01101000111: data <= 32'haae83440;
    11'b01101001000: data <= 32'h3ec9bbd9;
    11'b01101001001: data <= 32'h411cb8a1;
    11'b01101001010: data <= 32'h3db73b21;
    11'b01101001011: data <= 32'hb31b3dee;
    11'b01101001100: data <= 32'hb52e39c7;
    11'b01101001101: data <= 32'h3a17b26b;
    11'b01101001110: data <= 32'h3af5b95e;
    11'b01101001111: data <= 32'hb81dbd26;
    11'b01101010000: data <= 32'hbd87c02f;
    11'b01101010001: data <= 32'hb4f2bfbe;
    11'b01101010010: data <= 32'h3d2bb6da;
    11'b01101010011: data <= 32'h3ce63b12;
    11'b01101010100: data <= 32'hb65938a9;
    11'b01101010101: data <= 32'hbe91b642;
    11'b01101010110: data <= 32'hbea2b06c;
    11'b01101010111: data <= 32'hbd5a3c8d;
    11'b01101011000: data <= 32'hbcef3d53;
    11'b01101011001: data <= 32'hb93fb2a1;
    11'b01101011010: data <= 32'h3908bd98;
    11'b01101011011: data <= 32'h3daab674;
    11'b01101011100: data <= 32'h3ad63eb0;
    11'b01101011101: data <= 32'h274440c6;
    11'b01101011110: data <= 32'h35a13d47;
    11'b01101011111: data <= 32'h3cc23043;
    11'b01101100000: data <= 32'h3a4eb2c5;
    11'b01101100001: data <= 32'hb9b3b7c7;
    11'b01101100010: data <= 32'hbc6abcf5;
    11'b01101100011: data <= 32'h38a8be6e;
    11'b01101100100: data <= 32'h40afbb61;
    11'b01101100101: data <= 32'h3f95af24;
    11'b01101100110: data <= 32'hb1a6b3a2;
    11'b01101100111: data <= 32'hbdf3b92a;
    11'b01101101000: data <= 32'hbd00ad3c;
    11'b01101101001: data <= 32'hbacf3b43;
    11'b01101101010: data <= 32'hbcc73853;
    11'b01101101011: data <= 32'hbd8bbcd0;
    11'b01101101100: data <= 32'hb8d3c001;
    11'b01101101101: data <= 32'h358db68b;
    11'b01101101110: data <= 32'h36a43fa8;
    11'b01101101111: data <= 32'h2cc040e1;
    11'b01101110000: data <= 32'h35043cd2;
    11'b01101110001: data <= 32'h397c3522;
    11'b01101110010: data <= 32'h282e392e;
    11'b01101110011: data <= 32'hbc8c3abe;
    11'b01101110100: data <= 32'hbafeae1c;
    11'b01101110101: data <= 32'h3ccdbcad;
    11'b01101110110: data <= 32'h41aabc77;
    11'b01101110111: data <= 32'h4032b623;
    11'b01101111000: data <= 32'h2f2ab00c;
    11'b01101111001: data <= 32'hb973b384;
    11'b01101111010: data <= 32'ha26a2ef2;
    11'b01101111011: data <= 32'h326c37cd;
    11'b01101111100: data <= 32'hbb43b54a;
    11'b01101111101: data <= 32'hbf6abffc;
    11'b01101111110: data <= 32'hbd0bc0d0;
    11'b01101111111: data <= 32'h29c3b949;
    11'b01110000000: data <= 32'h37e03d66;
    11'b01110000001: data <= 32'h2c743df9;
    11'b01110000010: data <= 32'hb2553640;
    11'b01110000011: data <= 32'hb43a3424;
    11'b01110000100: data <= 32'hbae63dac;
    11'b01110000101: data <= 32'hbe4f3f8c;
    11'b01110000110: data <= 32'hbbbe3895;
    11'b01110000111: data <= 32'h3c04bc0e;
    11'b01110001000: data <= 32'h40a2bc33;
    11'b01110001001: data <= 32'h3e7b2c68;
    11'b01110001010: data <= 32'h346939ce;
    11'b01110001011: data <= 32'h34fe388a;
    11'b01110001100: data <= 32'h3d4036c4;
    11'b01110001101: data <= 32'h3c80354b;
    11'b01110001110: data <= 32'hb943b855;
    11'b01110001111: data <= 32'hbf99bfc6;
    11'b01110010000: data <= 32'hbc31c090;
    11'b01110010001: data <= 32'h3927bbf5;
    11'b01110010010: data <= 32'h3c4b3492;
    11'b01110010011: data <= 32'h31242d32;
    11'b01110010100: data <= 32'hb924b8fc;
    11'b01110010101: data <= 32'hbac42a7a;
    11'b01110010110: data <= 32'hbcc53ee1;
    11'b01110010111: data <= 32'hbede4022;
    11'b01110011000: data <= 32'hbd723587;
    11'b01110011001: data <= 32'h2903bd4e;
    11'b01110011010: data <= 32'h3c25bb6f;
    11'b01110011011: data <= 32'h39af39fc;
    11'b01110011100: data <= 32'h33373e51;
    11'b01110011101: data <= 32'h3b783c8b;
    11'b01110011110: data <= 32'h3fc8394d;
    11'b01110011111: data <= 32'h3d46390d;
    11'b01110100000: data <= 32'hb9bf317d;
    11'b01110100001: data <= 32'hbeb1bbb7;
    11'b01110100010: data <= 32'hb494be87;
    11'b01110100011: data <= 32'h3e73bcb9;
    11'b01110100100: data <= 32'h3ee1b91e;
    11'b01110100101: data <= 32'h3551bb92;
    11'b01110100110: data <= 32'hb8c2bcbb;
    11'b01110100111: data <= 32'hb80eac47;
    11'b01110101000: data <= 32'hb8cc3e1f;
    11'b01110101001: data <= 32'hbd8b3db6;
    11'b01110101010: data <= 32'hbf2bb84f;
    11'b01110101011: data <= 32'hbc73bf9e;
    11'b01110101100: data <= 32'hb3b0bb64;
    11'b01110101101: data <= 32'habd53c31;
    11'b01110101110: data <= 32'h2ba83eba;
    11'b01110101111: data <= 32'h3b5d3b80;
    11'b01110110000: data <= 32'h3e7338c8;
    11'b01110110001: data <= 32'h39aa3cd8;
    11'b01110110010: data <= 32'hbc6d3daa;
    11'b01110110011: data <= 32'hbdd6361e;
    11'b01110110100: data <= 32'h358dbabd;
    11'b01110110101: data <= 32'h4043bc83;
    11'b01110110110: data <= 32'h3f72bb5a;
    11'b01110110111: data <= 32'h369fbc1a;
    11'b01110111000: data <= 32'ha890bba3;
    11'b01110111001: data <= 32'h392f2c66;
    11'b01110111010: data <= 32'h39273c95;
    11'b01110111011: data <= 32'hb9ec38a4;
    11'b01110111100: data <= 32'hbff1bd5f;
    11'b01110111101: data <= 32'hbf0ac089;
    11'b01110111110: data <= 32'hba00bc11;
    11'b01110111111: data <= 32'hb2b3398c;
    11'b01111000000: data <= 32'ha78a3a7e;
    11'b01111000001: data <= 32'h3743ab01;
    11'b01111000010: data <= 32'h39c531d9;
    11'b01111000011: data <= 32'hb1a83ec7;
    11'b01111000100: data <= 32'hbe1c40de;
    11'b01111000101: data <= 32'hbdc43d16;
    11'b01111000110: data <= 32'h3524b6b6;
    11'b01111000111: data <= 32'h3ec1bb84;
    11'b01111001000: data <= 32'h3ce7b818;
    11'b01111001001: data <= 32'h33c5b43d;
    11'b01111001010: data <= 32'h3958b214;
    11'b01111001011: data <= 32'h3fc235fc;
    11'b01111001100: data <= 32'h3f343b5c;
    11'b01111001101: data <= 32'hb1ef3399;
    11'b01111001110: data <= 32'hbf7bbd6f;
    11'b01111001111: data <= 32'hbe57c006;
    11'b01111010000: data <= 32'hb463bc2c;
    11'b01111010001: data <= 32'h34c8adb9;
    11'b01111010010: data <= 32'h2a9bb87e;
    11'b01111010011: data <= 32'ha5cabd3a;
    11'b01111010100: data <= 32'h2a03b5c5;
    11'b01111010101: data <= 32'hb8933f32;
    11'b01111010110: data <= 32'hbe47414a;
    11'b01111010111: data <= 32'hbe443cca;
    11'b01111011000: data <= 32'hb60eb8ef;
    11'b01111011001: data <= 32'h3738ba5d;
    11'b01111011010: data <= 32'h2cfc3185;
    11'b01111011011: data <= 32'hb13a3926;
    11'b01111011100: data <= 32'h3c4236f4;
    11'b01111011101: data <= 32'h41303864;
    11'b01111011110: data <= 32'h405a3bfb;
    11'b01111011111: data <= 32'had7439a8;
    11'b01111100000: data <= 32'hbe62b6db;
    11'b01111100001: data <= 32'hbaafbc8a;
    11'b01111100010: data <= 32'h39b4baec;
    11'b01111100011: data <= 32'h3be6ba26;
    11'b01111100100: data <= 32'h31f2be6f;
    11'b01111100101: data <= 32'hb0d3c028;
    11'b01111100110: data <= 32'h316db97c;
    11'b01111100111: data <= 32'ha89a3e21;
    11'b01111101000: data <= 32'hbc1e400e;
    11'b01111101001: data <= 32'hbe8c3545;
    11'b01111101010: data <= 32'hbd15bcdc;
    11'b01111101011: data <= 32'hbab9ba29;
    11'b01111101100: data <= 32'hbb7638d9;
    11'b01111101101: data <= 32'hb8ac3b76;
    11'b01111101110: data <= 32'h3b8a34d2;
    11'b01111101111: data <= 32'h409534e3;
    11'b01111110000: data <= 32'h3e793cf2;
    11'b01111110001: data <= 32'hb7783ec1;
    11'b01111110010: data <= 32'hbd7b3b6c;
    11'b01111110011: data <= 32'haeb5ad87;
    11'b01111110100: data <= 32'h3d8fb81d;
    11'b01111110101: data <= 32'h3cccbb40;
    11'b01111110110: data <= 32'h2feabee6;
    11'b01111110111: data <= 32'h2e3cbfc6;
    11'b01111111000: data <= 32'h3c44b8c1;
    11'b01111111001: data <= 32'h3cd73c89;
    11'b01111111010: data <= 32'haf773c73;
    11'b01111111011: data <= 32'hbdfeb8d5;
    11'b01111111100: data <= 32'hbefcbe9f;
    11'b01111111101: data <= 32'hbd93ba07;
    11'b01111111110: data <= 32'hbcdf3835;
    11'b01111111111: data <= 32'hba1b34f6;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    