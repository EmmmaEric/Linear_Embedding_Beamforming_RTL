
module memory_rom_7(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbe50b1d3;
    11'b00000000001: data <= 32'hba91abf7;
    11'b00000000010: data <= 32'h3bf331ed;
    11'b00000000011: data <= 32'h3e0f3c6c;
    11'b00000000100: data <= 32'hb1af3eeb;
    11'b00000000101: data <= 32'hbfff3d1a;
    11'b00000000110: data <= 32'hbebf387b;
    11'b00000000111: data <= 32'h30853878;
    11'b00000001000: data <= 32'h3ccc3917;
    11'b00000001001: data <= 32'h3b1fb467;
    11'b00000001010: data <= 32'h3958bdb2;
    11'b00000001011: data <= 32'h3d3bbbe9;
    11'b00000001100: data <= 32'h3edf3b66;
    11'b00000001101: data <= 32'h3bc33f96;
    11'b00000001110: data <= 32'hb01f37dc;
    11'b00000001111: data <= 32'hb7acbe7e;
    11'b00000010000: data <= 32'hb723c017;
    11'b00000010001: data <= 32'hbad9bb8c;
    11'b00000010010: data <= 32'hbca3b603;
    11'b00000010011: data <= 32'hb43abbc0;
    11'b00000010100: data <= 32'h3ca4bcc4;
    11'b00000010101: data <= 32'h3c4daafe;
    11'b00000010110: data <= 32'hbb003d36;
    11'b00000010111: data <= 32'hc0e33df8;
    11'b00000011000: data <= 32'hbf343b08;
    11'b00000011001: data <= 32'hae033874;
    11'b00000011010: data <= 32'h365336bc;
    11'b00000011011: data <= 32'hb5b6b351;
    11'b00000011100: data <= 32'hb5cdba97;
    11'b00000011101: data <= 32'h3c4caceb;
    11'b00000011110: data <= 32'h407f3e7a;
    11'b00000011111: data <= 32'h3ecc404a;
    11'b00000100000: data <= 32'h347a3901;
    11'b00000100001: data <= 32'hb649bc6e;
    11'b00000100010: data <= 32'hb40dbc74;
    11'b00000100011: data <= 32'hb2f4b142;
    11'b00000100100: data <= 32'hb318b61a;
    11'b00000100101: data <= 32'h37a2bf42;
    11'b00000100110: data <= 32'h3d8dc09b;
    11'b00000100111: data <= 32'h3c00ba65;
    11'b00000101000: data <= 32'hba0f3c27;
    11'b00000101001: data <= 32'hbfca3d36;
    11'b00000101010: data <= 32'hbd6035ca;
    11'b00000101011: data <= 32'hb4edb362;
    11'b00000101100: data <= 32'hb942b1dc;
    11'b00000101101: data <= 32'hbee5b4a7;
    11'b00000101110: data <= 32'hbd45b785;
    11'b00000101111: data <= 32'h3a3e32f7;
    11'b00000110000: data <= 32'h407b3e42;
    11'b00000110001: data <= 32'h3dea3fff;
    11'b00000110010: data <= 32'hb2f03bb7;
    11'b00000110011: data <= 32'hba09a5bf;
    11'b00000110100: data <= 32'had4334d9;
    11'b00000110101: data <= 32'h36bb3aa9;
    11'b00000110110: data <= 32'h36b7b20e;
    11'b00000110111: data <= 32'h3a10c03e;
    11'b00000111000: data <= 32'h3dc6c107;
    11'b00000111001: data <= 32'h3d5bb97e;
    11'b00000111010: data <= 32'h31cf3c8f;
    11'b00000111011: data <= 32'hb9923b8a;
    11'b00000111100: data <= 32'hb7c3b7aa;
    11'b00000111101: data <= 32'hb500bc65;
    11'b00000111110: data <= 32'hbd46b91f;
    11'b00000111111: data <= 32'hc0ceb613;
    11'b00001000000: data <= 32'hbe70b93d;
    11'b00001000001: data <= 32'h395ab6df;
    11'b00001000010: data <= 32'h3f4a3911;
    11'b00001000011: data <= 32'h38d83da4;
    11'b00001000100: data <= 32'hbc943cdc;
    11'b00001000101: data <= 32'hbcea3b97;
    11'b00001000110: data <= 32'ha9793d75;
    11'b00001000111: data <= 32'h38433dce;
    11'b00001001000: data <= 32'h314d2911;
    11'b00001001001: data <= 32'h32a7bf38;
    11'b00001001010: data <= 32'h3c9dbf48;
    11'b00001001011: data <= 32'h3f3e2ef4;
    11'b00001001100: data <= 32'h3d6d3e01;
    11'b00001001101: data <= 32'h38a6397f;
    11'b00001001110: data <= 32'h34bbbbae;
    11'b00001001111: data <= 32'hae83bd1c;
    11'b00001010000: data <= 32'hbcfab735;
    11'b00001010001: data <= 32'hc021b4ef;
    11'b00001010010: data <= 32'hbc78bcee;
    11'b00001010011: data <= 32'h3a97bea2;
    11'b00001010100: data <= 32'h3d68b964;
    11'b00001010101: data <= 32'hb26a394a;
    11'b00001010110: data <= 32'hbed43cb1;
    11'b00001010111: data <= 32'hbd483cde;
    11'b00001011000: data <= 32'haaa13ddf;
    11'b00001011001: data <= 32'h28563d62;
    11'b00001011010: data <= 32'hbb752fdf;
    11'b00001011011: data <= 32'hbbb7bcbf;
    11'b00001011100: data <= 32'h38a7baad;
    11'b00001011101: data <= 32'h40193b3b;
    11'b00001011110: data <= 32'h40093efd;
    11'b00001011111: data <= 32'h3c783916;
    11'b00001100000: data <= 32'h3855b9c2;
    11'b00001100001: data <= 32'h313cb7e8;
    11'b00001100010: data <= 32'hb8c13753;
    11'b00001100011: data <= 32'hbc572685;
    11'b00001100100: data <= 32'hb4bfbf11;
    11'b00001100101: data <= 32'h3c42c160;
    11'b00001100110: data <= 32'h3c84be44;
    11'b00001100111: data <= 32'hb54131f8;
    11'b00001101000: data <= 32'hbd6f3af3;
    11'b00001101001: data <= 32'hba04397f;
    11'b00001101010: data <= 32'h2c0c3964;
    11'b00001101011: data <= 32'hb996398a;
    11'b00001101100: data <= 32'hc06a293d;
    11'b00001101101: data <= 32'hc02ab9ca;
    11'b00001101110: data <= 32'h282fb534;
    11'b00001101111: data <= 32'h3f883bf9;
    11'b00001110000: data <= 32'h3f1c3e0e;
    11'b00001110001: data <= 32'h39313954;
    11'b00001110010: data <= 32'h317729de;
    11'b00001110011: data <= 32'h35213a98;
    11'b00001110100: data <= 32'h2fd53e86;
    11'b00001110101: data <= 32'hb42f3816;
    11'b00001110110: data <= 32'h3037bf7e;
    11'b00001110111: data <= 32'h3c41c1bd;
    11'b00001111000: data <= 32'h3cc2be10;
    11'b00001111001: data <= 32'h34c73402;
    11'b00001111010: data <= 32'hb2ce3806;
    11'b00001111011: data <= 32'h3498b2bf;
    11'b00001111100: data <= 32'h3614b580;
    11'b00001111101: data <= 32'hbc812df2;
    11'b00001111110: data <= 32'hc1b3a549;
    11'b00001111111: data <= 32'hc0f1b956;
    11'b00010000000: data <= 32'hb15bb963;
    11'b00010000001: data <= 32'h3db931d0;
    11'b00010000010: data <= 32'h3ae13a01;
    11'b00010000011: data <= 32'hb65338a1;
    11'b00010000100: data <= 32'hb6eb3a0f;
    11'b00010000101: data <= 32'h35d23f64;
    11'b00010000110: data <= 32'h370440c2;
    11'b00010000111: data <= 32'hb37c3b0e;
    11'b00010001000: data <= 32'hb4a4bdf5;
    11'b00010001001: data <= 32'h38eec048;
    11'b00010001010: data <= 32'h3d48b91a;
    11'b00010001011: data <= 32'h3cc839be;
    11'b00010001100: data <= 32'h3c18341c;
    11'b00010001101: data <= 32'h3cecbae3;
    11'b00010001110: data <= 32'h3a4aba46;
    11'b00010001111: data <= 32'hbb98308f;
    11'b00010010000: data <= 32'hc0f731c8;
    11'b00010010001: data <= 32'hbfbcbb50;
    11'b00010010010: data <= 32'h2c0bbe72;
    11'b00010010011: data <= 32'h3bc6bc4f;
    11'b00010010100: data <= 32'had91b1f7;
    11'b00010010101: data <= 32'hbcca34ac;
    11'b00010010110: data <= 32'hb9653b18;
    11'b00010010111: data <= 32'h37433fb8;
    11'b00010011000: data <= 32'h33f5408b;
    11'b00010011001: data <= 32'hbc263b70;
    11'b00010011010: data <= 32'hbd9dbb03;
    11'b00010011011: data <= 32'hb0fbbc25;
    11'b00010011100: data <= 32'h3d1a3606;
    11'b00010011101: data <= 32'h3ebc3c7b;
    11'b00010011110: data <= 32'h3e2f305e;
    11'b00010011111: data <= 32'h3e17bb3c;
    11'b00010100000: data <= 32'h3c44b4b2;
    11'b00010100001: data <= 32'hb4a13bd4;
    11'b00010100010: data <= 32'hbda239b9;
    11'b00010100011: data <= 32'hbb5cbc8c;
    11'b00010100100: data <= 32'h3760c0e1;
    11'b00010100101: data <= 32'h39a8bfd8;
    11'b00010100110: data <= 32'hb78fba09;
    11'b00010100111: data <= 32'hbc8ead61;
    11'b00010101000: data <= 32'hb239352f;
    11'b00010101001: data <= 32'h3a133c3c;
    11'b00010101010: data <= 32'hb1213dd5;
    11'b00010101011: data <= 32'hc02e3998;
    11'b00010101100: data <= 32'hc108b648;
    11'b00010101101: data <= 32'hbab9b4b9;
    11'b00010101110: data <= 32'h3bd63a0d;
    11'b00010101111: data <= 32'h3d863bf9;
    11'b00010110000: data <= 32'h3c139cd9;
    11'b00010110001: data <= 32'h3c21b76e;
    11'b00010110010: data <= 32'h3c623a4c;
    11'b00010110011: data <= 32'h36f5404a;
    11'b00010110100: data <= 32'hb60b3d7b;
    11'b00010110101: data <= 32'hb2aabc41;
    11'b00010110110: data <= 32'h38bcc110;
    11'b00010110111: data <= 32'h38f9bf7a;
    11'b00010111000: data <= 32'hb150b8f3;
    11'b00010111001: data <= 32'hb3d4b5ba;
    11'b00010111010: data <= 32'h3aadb8a1;
    11'b00010111011: data <= 32'h3d15b07b;
    11'b00010111100: data <= 32'hb5d838b0;
    11'b00010111101: data <= 32'hc13c37c7;
    11'b00010111110: data <= 32'hc1c3b308;
    11'b00010111111: data <= 32'hbc14b552;
    11'b00011000000: data <= 32'h38963297;
    11'b00011000001: data <= 32'h373c3413;
    11'b00011000010: data <= 32'hb1ddb4d2;
    11'b00011000011: data <= 32'h3194a125;
    11'b00011000100: data <= 32'h3bcf3eb1;
    11'b00011000101: data <= 32'h3ab341c8;
    11'b00011000110: data <= 32'haae83f19;
    11'b00011000111: data <= 32'hb5a1b968;
    11'b00011001000: data <= 32'h31fcbf1b;
    11'b00011001001: data <= 32'h3856badb;
    11'b00011001010: data <= 32'h37292ce0;
    11'b00011001011: data <= 32'h3aadb70e;
    11'b00011001100: data <= 32'h3f2bbd2a;
    11'b00011001101: data <= 32'h3f0cbae0;
    11'b00011001110: data <= 32'hb0413587;
    11'b00011001111: data <= 32'hc06b38f0;
    11'b00011010000: data <= 32'hc078b446;
    11'b00011010001: data <= 32'hb8c7bbc5;
    11'b00011010010: data <= 32'h343fbb02;
    11'b00011010011: data <= 32'hb857b9a8;
    11'b00011010100: data <= 32'hbcfdb9c1;
    11'b00011010101: data <= 32'hb5d62325;
    11'b00011010110: data <= 32'h3bbe3ecc;
    11'b00011010111: data <= 32'h3a9d4167;
    11'b00011011000: data <= 32'hb8663eb1;
    11'b00011011001: data <= 32'hbd11b21e;
    11'b00011011010: data <= 32'hb8e4b90e;
    11'b00011011011: data <= 32'h353c3672;
    11'b00011011100: data <= 32'h3a443a3b;
    11'b00011011101: data <= 32'h3d25b701;
    11'b00011011110: data <= 32'h4012bdf6;
    11'b00011011111: data <= 32'h3fc8b96d;
    11'b00011100000: data <= 32'h36e73bb2;
    11'b00011100001: data <= 32'hbc633cac;
    11'b00011100010: data <= 32'hbbf1b4c3;
    11'b00011100011: data <= 32'h2e2ebe6c;
    11'b00011100100: data <= 32'h3099beb2;
    11'b00011100101: data <= 32'hbc3fbd09;
    11'b00011100110: data <= 32'hbdfebc3b;
    11'b00011100111: data <= 32'hb00db7e8;
    11'b00011101000: data <= 32'h3d163a56;
    11'b00011101001: data <= 32'h38f73ebd;
    11'b00011101010: data <= 32'hbd833ca4;
    11'b00011101011: data <= 32'hc08e3072;
    11'b00011101100: data <= 32'hbd3a3329;
    11'b00011101101: data <= 32'h21573c5e;
    11'b00011101110: data <= 32'h37d53b5a;
    11'b00011101111: data <= 32'h39c6b86e;
    11'b00011110000: data <= 32'h3d7ebd03;
    11'b00011110001: data <= 32'h3ee130f5;
    11'b00011110010: data <= 32'h3c014005;
    11'b00011110011: data <= 32'h28233f6b;
    11'b00011110100: data <= 32'h2699b0d3;
    11'b00011110101: data <= 32'h381ebea4;
    11'b00011110110: data <= 32'h2f1bbe29;
    11'b00011110111: data <= 32'hbb9ebbe9;
    11'b00011111000: data <= 32'hbaf6bc78;
    11'b00011111001: data <= 32'h3a21bd03;
    11'b00011111010: data <= 32'h3f4db7e1;
    11'b00011111011: data <= 32'h3840381a;
    11'b00011111100: data <= 32'hbf4d3920;
    11'b00011111101: data <= 32'hc1313355;
    11'b00011111110: data <= 32'hbd9135f8;
    11'b00011111111: data <= 32'hb3663a9b;
    11'b00100000000: data <= 32'hb51b3567;
    11'b00100000001: data <= 32'hb873bb26;
    11'b00100000010: data <= 32'h3359bb95;
    11'b00100000011: data <= 32'h3d233b66;
    11'b00100000100: data <= 32'h3d2d416a;
    11'b00100000101: data <= 32'h383c4067;
    11'b00100000110: data <= 32'h31e63012;
    11'b00100000111: data <= 32'h34d0bbf5;
    11'b00100001000: data <= 32'h9969b758;
    11'b00100001001: data <= 32'hb817a786;
    11'b00100001010: data <= 32'h2bbdbb1d;
    11'b00100001011: data <= 32'h3eaebf5b;
    11'b00100001100: data <= 32'h4098bd7b;
    11'b00100001101: data <= 32'h39ada9a9;
    11'b00100001110: data <= 32'hbde53860;
    11'b00100001111: data <= 32'hbf8c3242;
    11'b00100010000: data <= 32'hb9dcacff;
    11'b00100010001: data <= 32'hb3deace1;
    11'b00100010010: data <= 32'hbcb8b87f;
    11'b00100010011: data <= 32'hbf12bd4f;
    11'b00100010100: data <= 32'hb916bb62;
    11'b00100010101: data <= 32'h3c123bca;
    11'b00100010110: data <= 32'h3d1440ed;
    11'b00100010111: data <= 32'h33423f9b;
    11'b00100011000: data <= 32'hb829358f;
    11'b00100011001: data <= 32'hb6b224f3;
    11'b00100011010: data <= 32'hb4193b83;
    11'b00100011011: data <= 32'hb32a3c05;
    11'b00100011100: data <= 32'h3806b8cd;
    11'b00100011101: data <= 32'h3f7cbffc;
    11'b00100011110: data <= 32'h40a6bd88;
    11'b00100011111: data <= 32'h3c313553;
    11'b00100100000: data <= 32'hb7b23bf3;
    11'b00100100001: data <= 32'hb82032db;
    11'b00100100010: data <= 32'h34aab8fc;
    11'b00100100011: data <= 32'hac08baa8;
    11'b00100100100: data <= 32'hbe89bc54;
    11'b00100100101: data <= 32'hc06bbe3a;
    11'b00100100110: data <= 32'hb951bd02;
    11'b00100100111: data <= 32'h3cbe3177;
    11'b00100101000: data <= 32'h3c713d51;
    11'b00100101001: data <= 32'hb7ae3c46;
    11'b00100101010: data <= 32'hbdd435d2;
    11'b00100101011: data <= 32'hbc5a3a57;
    11'b00100101100: data <= 32'hb8173f47;
    11'b00100101101: data <= 32'hb6423dc2;
    11'b00100101110: data <= 32'h25eab85b;
    11'b00100101111: data <= 32'h3c6ebf2d;
    11'b00100110000: data <= 32'h3f36b98d;
    11'b00100110001: data <= 32'h3d393d1a;
    11'b00100110010: data <= 32'h386e3e9c;
    11'b00100110011: data <= 32'h398e356f;
    11'b00100110100: data <= 32'h3c1fba02;
    11'b00100110101: data <= 32'h2f42ba17;
    11'b00100110110: data <= 32'hbe2cb9da;
    11'b00100110111: data <= 32'hbefabd6b;
    11'b00100111000: data <= 32'h2dbcbede;
    11'b00100111001: data <= 32'h3ecfbc0d;
    11'b00100111010: data <= 32'h3c1ea827;
    11'b00100111011: data <= 32'hbba33294;
    11'b00100111100: data <= 32'hbf4332ae;
    11'b00100111101: data <= 32'hbc733b88;
    11'b00100111110: data <= 32'hb8483eee;
    11'b00100111111: data <= 32'hbb7a3c20;
    11'b00101000000: data <= 32'hbc9ebaa4;
    11'b00101000001: data <= 32'hb2f2be11;
    11'b00101000010: data <= 32'h3c0c2c00;
    11'b00101000011: data <= 32'h3d4b3ff5;
    11'b00101000100: data <= 32'h3c1f3fd6;
    11'b00101000101: data <= 32'h3c303728;
    11'b00101000110: data <= 32'h3c1eb501;
    11'b00101000111: data <= 32'h2d293338;
    11'b00101001000: data <= 32'hbc903656;
    11'b00101001001: data <= 32'hbae5ba2f;
    11'b00101001010: data <= 32'h3be9c003;
    11'b00101001011: data <= 32'h404dbf6a;
    11'b00101001100: data <= 32'h3c56ba5f;
    11'b00101001101: data <= 32'hba4fb094;
    11'b00101001110: data <= 32'hbcc42b7f;
    11'b00101001111: data <= 32'hb4db383f;
    11'b00101010000: data <= 32'hb2c33b49;
    11'b00101010001: data <= 32'hbdf9312c;
    11'b00101010010: data <= 32'hc0a1bd02;
    11'b00101010011: data <= 32'hbd32bda6;
    11'b00101010100: data <= 32'h3736341c;
    11'b00101010101: data <= 32'h3c913f4c;
    11'b00101010110: data <= 32'h3a1a3e1f;
    11'b00101010111: data <= 32'h374535ae;
    11'b00101011000: data <= 32'h35f9367e;
    11'b00101011001: data <= 32'hb13c3e44;
    11'b00101011010: data <= 32'hba7f3e9d;
    11'b00101011011: data <= 32'hb504b109;
    11'b00101011100: data <= 32'h3d0cbfdf;
    11'b00101011101: data <= 32'h4028bf8e;
    11'b00101011110: data <= 32'h3c95b87c;
    11'b00101011111: data <= 32'hacd43268;
    11'b00101100000: data <= 32'h2fa62b64;
    11'b00101100001: data <= 32'h3b8fa67f;
    11'b00101100010: data <= 32'h35222dab;
    11'b00101100011: data <= 32'hbedfb6c1;
    11'b00101100100: data <= 32'hc18abda8;
    11'b00101100101: data <= 32'hbdfcbe07;
    11'b00101100110: data <= 32'h3785b49c;
    11'b00101100111: data <= 32'h3b863a05;
    11'b00101101000: data <= 32'h2c1d37a9;
    11'b00101101001: data <= 32'hb81620ed;
    11'b00101101010: data <= 32'hb58c3b68;
    11'b00101101011: data <= 32'hb61240e7;
    11'b00101101100: data <= 32'hba544090;
    11'b00101101101: data <= 32'hb87f2dfe;
    11'b00101101110: data <= 32'h3888bec5;
    11'b00101101111: data <= 32'h3d69bcdf;
    11'b00101110000: data <= 32'h3c2a3600;
    11'b00101110001: data <= 32'h39873b1b;
    11'b00101110010: data <= 32'h3d503143;
    11'b00101110011: data <= 32'h3f9db4bc;
    11'b00101110100: data <= 32'h39e9a94d;
    11'b00101110101: data <= 32'hbe15b0ab;
    11'b00101110110: data <= 32'hc0a7bc22;
    11'b00101110111: data <= 32'hba45be7e;
    11'b00101111000: data <= 32'h3be8bcc9;
    11'b00101111001: data <= 32'h3aceb8d3;
    11'b00101111010: data <= 32'hb81bb900;
    11'b00101111011: data <= 32'hbc27b6e5;
    11'b00101111100: data <= 32'hb7373b7a;
    11'b00101111101: data <= 32'hb42640c8;
    11'b00101111110: data <= 32'hbc0e3fcf;
    11'b00101111111: data <= 32'hbddeb116;
    11'b00110000000: data <= 32'hb9f5bd9f;
    11'b00110000001: data <= 32'h34efb63e;
    11'b00110000010: data <= 32'h39e33ce8;
    11'b00110000011: data <= 32'h3bf63d1c;
    11'b00110000100: data <= 32'h3ed93136;
    11'b00110000101: data <= 32'h400bb08e;
    11'b00110000110: data <= 32'h3a423975;
    11'b00110000111: data <= 32'hbc643bac;
    11'b00110001000: data <= 32'hbd97b254;
    11'b00110001001: data <= 32'h3327be42;
    11'b00110001010: data <= 32'h3e12bf58;
    11'b00110001011: data <= 32'h3a9fbd9b;
    11'b00110001100: data <= 32'hb8bfbc8a;
    11'b00110001101: data <= 32'hb94cb9a8;
    11'b00110001110: data <= 32'h353137c0;
    11'b00110001111: data <= 32'h34ec3e2d;
    11'b00110010000: data <= 32'hbcdb3c07;
    11'b00110010001: data <= 32'hc0cfb93c;
    11'b00110010010: data <= 32'hbf73bd00;
    11'b00110010011: data <= 32'hb74122e7;
    11'b00110010100: data <= 32'h35fe3d2d;
    11'b00110010101: data <= 32'h394b3b2b;
    11'b00110010110: data <= 32'h3c74b0dc;
    11'b00110010111: data <= 32'h3d50331a;
    11'b00110011000: data <= 32'h37b33f28;
    11'b00110011001: data <= 32'hb9ea4080;
    11'b00110011010: data <= 32'hb9673935;
    11'b00110011011: data <= 32'h39b5bd2e;
    11'b00110011100: data <= 32'h3e09bf1b;
    11'b00110011101: data <= 32'h398ebcb4;
    11'b00110011110: data <= 32'hb312ba65;
    11'b00110011111: data <= 32'h368db972;
    11'b00110100000: data <= 32'h3e6cadd3;
    11'b00110100001: data <= 32'h3c6238a4;
    11'b00110100010: data <= 32'hbcaa3327;
    11'b00110100011: data <= 32'hc179bb2a;
    11'b00110100100: data <= 32'hc02bbcbb;
    11'b00110100101: data <= 32'hb7d9b2c3;
    11'b00110100110: data <= 32'h311b376b;
    11'b00110100111: data <= 32'hab41b1d5;
    11'b00110101000: data <= 32'h28c0ba21;
    11'b00110101001: data <= 32'h36e336fe;
    11'b00110101010: data <= 32'h318a410e;
    11'b00110101011: data <= 32'hb8be41d6;
    11'b00110101100: data <= 32'hb9083c07;
    11'b00110101101: data <= 32'h3430bbaa;
    11'b00110101110: data <= 32'h3a28bc4d;
    11'b00110101111: data <= 32'h351eb103;
    11'b00110110000: data <= 32'h330128bd;
    11'b00110110001: data <= 32'h3dd2b7a8;
    11'b00110110010: data <= 32'h413db745;
    11'b00110110011: data <= 32'h3eac31e2;
    11'b00110110100: data <= 32'hbad93416;
    11'b00110110101: data <= 32'hc07eb830;
    11'b00110110110: data <= 32'hbd41bc29;
    11'b00110110111: data <= 32'h307bba40;
    11'b00110111000: data <= 32'h30fdb9b5;
    11'b00110111001: data <= 32'hb99ebd69;
    11'b00110111010: data <= 32'hb9d1bda0;
    11'b00110111011: data <= 32'h2d5d348a;
    11'b00110111100: data <= 32'h342840ce;
    11'b00110111101: data <= 32'hb8a2411d;
    11'b00110111110: data <= 32'hbcc6397b;
    11'b00110111111: data <= 32'hbaddb9e3;
    11'b00111000000: data <= 32'hb590b234;
    11'b00111000001: data <= 32'hb3203b3c;
    11'b00111000010: data <= 32'h350b394c;
    11'b00111000011: data <= 32'h3f09b6c2;
    11'b00111000100: data <= 32'h4177b80e;
    11'b00111000101: data <= 32'h3ec3389b;
    11'b00111000110: data <= 32'hb7803c9f;
    11'b00111000111: data <= 32'hbd15361a;
    11'b00111001000: data <= 32'hafdcb9c0;
    11'b00111001001: data <= 32'h3b2abcb1;
    11'b00111001010: data <= 32'h32babdab;
    11'b00111001011: data <= 32'hbba8bf8f;
    11'b00111001100: data <= 32'hb95bbede;
    11'b00111001101: data <= 32'h3924b16e;
    11'b00111001110: data <= 32'h3b0e3e0c;
    11'b00111001111: data <= 32'hb80b3dd2;
    11'b00111010000: data <= 32'hbf6aa4d6;
    11'b00111010001: data <= 32'hbf77b95d;
    11'b00111010010: data <= 32'hbca835b2;
    11'b00111010011: data <= 32'hb96a3d1a;
    11'b00111010100: data <= 32'hac413812;
    11'b00111010101: data <= 32'h3c74ba2c;
    11'b00111010110: data <= 32'h3fa7b69f;
    11'b00111010111: data <= 32'h3cd43d8a;
    11'b00111011000: data <= 32'hb27d40a5;
    11'b00111011001: data <= 32'hb6d13d3a;
    11'b00111011010: data <= 32'h393fb4d2;
    11'b00111011011: data <= 32'h3c80bc12;
    11'b00111011100: data <= 32'h2c4dbc90;
    11'b00111011101: data <= 32'hbac0bddc;
    11'b00111011110: data <= 32'h2dfcbe2f;
    11'b00111011111: data <= 32'h3f25b946;
    11'b00111100000: data <= 32'h3f0b3720;
    11'b00111100001: data <= 32'hb439365f;
    11'b00111100010: data <= 32'hc016b815;
    11'b00111100011: data <= 32'hc010b8f9;
    11'b00111100100: data <= 32'hbc9b35f8;
    11'b00111100101: data <= 32'hba623a13;
    11'b00111100110: data <= 32'hb9c1b6af;
    11'b00111100111: data <= 32'haa63bded;
    11'b00111101000: data <= 32'h3a1ab6d0;
    11'b00111101001: data <= 32'h39273fc6;
    11'b00111101010: data <= 32'hae7f41dc;
    11'b00111101011: data <= 32'hb1183e9c;
    11'b00111101100: data <= 32'h38309893;
    11'b00111101101: data <= 32'h3873b59c;
    11'b00111101110: data <= 32'hb660a9c7;
    11'b00111101111: data <= 32'hb93bb66c;
    11'b00111110000: data <= 32'h3b6dbc61;
    11'b00111110001: data <= 32'h4177bba5;
    11'b00111110010: data <= 32'h40b8b0c1;
    11'b00111110011: data <= 32'h2c3e2eed;
    11'b00111110100: data <= 32'hbe34b54e;
    11'b00111110101: data <= 32'hbcc3b66f;
    11'b00111110110: data <= 32'hb5372c2c;
    11'b00111110111: data <= 32'hb891b1cd;
    11'b00111111000: data <= 32'hbd24be12;
    11'b00111111001: data <= 32'hbbeac05e;
    11'b00111111010: data <= 32'h2e1cb93e;
    11'b00111111011: data <= 32'h38183f1d;
    11'b00111111100: data <= 32'ha8994101;
    11'b00111111101: data <= 32'hb7573cb0;
    11'b00111111110: data <= 32'hb5652539;
    11'b00111111111: data <= 32'hb7b0373b;
    11'b01000000000: data <= 32'hbc1f3cb1;
    11'b01000000001: data <= 32'hb97b384f;
    11'b01000000010: data <= 32'h3ca1ba62;
    11'b01000000011: data <= 32'h4194bc1f;
    11'b01000000100: data <= 32'h4088a3ac;
    11'b01000000101: data <= 32'h34b839d4;
    11'b01000000110: data <= 32'hb926379e;
    11'b01000000111: data <= 32'h30932698;
    11'b01000001000: data <= 32'h39e0b0f2;
    11'b01000001001: data <= 32'hb42eba36;
    11'b01000001010: data <= 32'hbe24c004;
    11'b01000001011: data <= 32'hbcb6c0da;
    11'b01000001100: data <= 32'h35b9bbfd;
    11'b01000001101: data <= 32'h3c0e3b80;
    11'b01000001110: data <= 32'h30b43d15;
    11'b01000001111: data <= 32'hbb4e31b9;
    11'b01000010000: data <= 32'hbcd2b197;
    11'b01000010001: data <= 32'hbd093bcb;
    11'b01000010010: data <= 32'hbdde3f1c;
    11'b01000010011: data <= 32'hbc0b3992;
    11'b01000010100: data <= 32'h3852bbfd;
    11'b01000010101: data <= 32'h3f6ebc26;
    11'b01000010110: data <= 32'h3e123886;
    11'b01000010111: data <= 32'h34e13ee9;
    11'b01000011000: data <= 32'h31173d77;
    11'b01000011001: data <= 32'h3c953789;
    11'b01000011010: data <= 32'h3d2819c1;
    11'b01000011011: data <= 32'hb33eb807;
    11'b01000011100: data <= 32'hbe04bdf3;
    11'b01000011101: data <= 32'hb940c00d;
    11'b01000011110: data <= 32'h3d39bcff;
    11'b01000011111: data <= 32'h3f69ad06;
    11'b01000100000: data <= 32'h373e09a2;
    11'b01000100001: data <= 32'hbc30b92f;
    11'b01000100010: data <= 32'hbd63b553;
    11'b01000100011: data <= 32'hbcaf3c36;
    11'b01000100100: data <= 32'hbd9d3e0a;
    11'b01000100101: data <= 32'hbdd3a09e;
    11'b01000100110: data <= 32'hb893bea2;
    11'b01000100111: data <= 32'h3809bc8d;
    11'b01000101000: data <= 32'h38e93c16;
    11'b01000101001: data <= 32'h31874091;
    11'b01000101010: data <= 32'h37753ea1;
    11'b01000101011: data <= 32'h3d11391b;
    11'b01000101100: data <= 32'h3bbe3807;
    11'b01000101101: data <= 32'hb8fc3860;
    11'b01000101110: data <= 32'hbdabb39e;
    11'b01000101111: data <= 32'h2915bcf3;
    11'b01000110000: data <= 32'h405bbd2c;
    11'b01000110001: data <= 32'h40d4b987;
    11'b01000110010: data <= 32'h39a1b860;
    11'b01000110011: data <= 32'hb961b9fb;
    11'b01000110100: data <= 32'hb850b2b1;
    11'b01000110101: data <= 32'hb1c13ad1;
    11'b01000110110: data <= 32'hbade39e8;
    11'b01000110111: data <= 32'hbf0ebc0b;
    11'b01000111000: data <= 32'hbe0cc0ad;
    11'b01000111001: data <= 32'hb6bfbd5a;
    11'b01000111010: data <= 32'h31903b69;
    11'b01000111011: data <= 32'h2efe3f80;
    11'b01000111100: data <= 32'h344a3c22;
    11'b01000111101: data <= 32'h38cf35f6;
    11'b01000111110: data <= 32'h2aec3c39;
    11'b01000111111: data <= 32'hbcf73f04;
    11'b01001000000: data <= 32'hbdd93bab;
    11'b01001000001: data <= 32'h34a7b8dd;
    11'b01001000010: data <= 32'h407bbcd0;
    11'b01001000011: data <= 32'h4069b92c;
    11'b01001000100: data <= 32'h3978b09d;
    11'b01001000101: data <= 32'h1cfbae01;
    11'b01001000110: data <= 32'h3a3c3287;
    11'b01001000111: data <= 32'h3c863976;
    11'b01001001000: data <= 32'hb2623142;
    11'b01001001001: data <= 32'hbf43bdfc;
    11'b01001001010: data <= 32'hbf18c0fd;
    11'b01001001011: data <= 32'hb655bdea;
    11'b01001001100: data <= 32'h37c33498;
    11'b01001001101: data <= 32'h34373945;
    11'b01001001110: data <= 32'haf0ab26f;
    11'b01001001111: data <= 32'hb293b1b6;
    11'b01001010000: data <= 32'hb9a63d6e;
    11'b01001010001: data <= 32'hbe7e40d5;
    11'b01001010010: data <= 32'hbe8d3d7a;
    11'b01001010011: data <= 32'hb10db8a4;
    11'b01001010100: data <= 32'h3d4abca0;
    11'b01001010101: data <= 32'h3cecb101;
    11'b01001010110: data <= 32'h35793a0c;
    11'b01001010111: data <= 32'h38983a15;
    11'b01001011000: data <= 32'h3f5138f9;
    11'b01001011001: data <= 32'h3fd039f2;
    11'b01001011010: data <= 32'h2e7d34e8;
    11'b01001011011: data <= 32'hbecebbef;
    11'b01001011100: data <= 32'hbd62bf92;
    11'b01001011101: data <= 32'h36bbbd95;
    11'b01001011110: data <= 32'h3d0fb7df;
    11'b01001011111: data <= 32'h3879b937;
    11'b01001100000: data <= 32'hb4aabd3c;
    11'b01001100001: data <= 32'hb701b91b;
    11'b01001100010: data <= 32'hb9173d48;
    11'b01001100011: data <= 32'hbd92407c;
    11'b01001100100: data <= 32'hbf1d3a99;
    11'b01001100101: data <= 32'hbc27bc9b;
    11'b01001100110: data <= 32'hac0dbd03;
    11'b01001100111: data <= 32'h28c234eb;
    11'b01001101000: data <= 32'hafd43d74;
    11'b01001101001: data <= 32'h39e03c47;
    11'b01001101010: data <= 32'h40153948;
    11'b01001101011: data <= 32'h3f4c3bdb;
    11'b01001101100: data <= 32'hb1843c90;
    11'b01001101101: data <= 32'hbe6b3488;
    11'b01001101110: data <= 32'hb963ba89;
    11'b01001101111: data <= 32'h3d3cbc57;
    11'b01001110000: data <= 32'h3f5ebb72;
    11'b01001110001: data <= 32'h39bfbd28;
    11'b01001110010: data <= 32'hb031be88;
    11'b01001110011: data <= 32'h31a4b96c;
    11'b01001110100: data <= 32'h35f63c63;
    11'b01001110101: data <= 32'hb8943e11;
    11'b01001110110: data <= 32'hbee5b119;
    11'b01001110111: data <= 32'hbf23bf5a;
    11'b01001111000: data <= 32'hbc4ebd93;
    11'b01001111001: data <= 32'hb946360a;
    11'b01001111010: data <= 32'hb6513c7e;
    11'b01001111011: data <= 32'h37e136fe;
    11'b01001111100: data <= 32'h3dc3308b;
    11'b01001111101: data <= 32'h3bb33cb7;
    11'b01001111110: data <= 32'hba4a4048;
    11'b01001111111: data <= 32'hbe783e41;
    11'b01010000000: data <= 32'hb4d12e37;
    11'b01010000001: data <= 32'h3e0eb9ea;
    11'b01010000010: data <= 32'h3e89ba85;
    11'b01010000011: data <= 32'h37a0bbb9;
    11'b01010000100: data <= 32'h32cbbc47;
    11'b01010000101: data <= 32'h3d26b4a8;
    11'b01010000110: data <= 32'h3f0e3b4d;
    11'b01010000111: data <= 32'h363b3ae6;
    11'b01010001000: data <= 32'hbdecba16;
    11'b01010001001: data <= 32'hbfc8c004;
    11'b01010001010: data <= 32'hbc91bd66;
    11'b01010001011: data <= 32'hb7b12981;
    11'b01010001100: data <= 32'hb4cd2ef3;
    11'b01010001101: data <= 32'h2ed9baf9;
    11'b01010001110: data <= 32'h38b9b9c4;
    11'b01010001111: data <= 32'h2f283c9f;
    11'b01010010000: data <= 32'hbcc6415b;
    11'b01010010001: data <= 32'hbe974025;
    11'b01010010010: data <= 32'hb7ae34d1;
    11'b01010010011: data <= 32'h3a4fb8bb;
    11'b01010010100: data <= 32'h38c1b501;
    11'b01010010101: data <= 32'hb19aaad1;
    11'b01010010110: data <= 32'h3706b0f5;
    11'b01010010111: data <= 32'h4062311a;
    11'b01010011000: data <= 32'h41633af1;
    11'b01010011001: data <= 32'h3b453a30;
    11'b01010011010: data <= 32'hbcdeb70f;
    11'b01010011011: data <= 32'hbdf7bd6e;
    11'b01010011100: data <= 32'hb56fbbbf;
    11'b01010011101: data <= 32'h352fb633;
    11'b01010011110: data <= 32'h2660bc2f;
    11'b01010011111: data <= 32'hb0a6c031;
    11'b01010100000: data <= 32'h3157bdc0;
    11'b01010100001: data <= 32'h1f7c3b63;
    11'b01010100010: data <= 32'hbb7b40eb;
    11'b01010100011: data <= 32'hbe0f3e45;
    11'b01010100100: data <= 32'hbc11b415;
    11'b01010100101: data <= 32'hb6ecb99c;
    11'b01010100110: data <= 32'hb9c6324f;
    11'b01010100111: data <= 32'hbb7139a6;
    11'b01010101000: data <= 32'h35c83509;
    11'b01010101001: data <= 32'h40af322b;
    11'b01010101010: data <= 32'h41403af2;
    11'b01010101011: data <= 32'h398d3d1d;
    11'b01010101100: data <= 32'hbc6f394d;
    11'b01010101101: data <= 32'hba49b11d;
    11'b01010101110: data <= 32'h3954b57b;
    11'b01010101111: data <= 32'h3c2db868;
    11'b01010110000: data <= 32'h3266be6b;
    11'b01010110001: data <= 32'hb1d9c103;
    11'b01010110010: data <= 32'h379dbe56;
    11'b01010110011: data <= 32'h3abb393a;
    11'b01010110100: data <= 32'h99593ed3;
    11'b01010110101: data <= 32'hbc8937f1;
    11'b01010110110: data <= 32'hbdd5bc42;
    11'b01010110111: data <= 32'hbd6abafa;
    11'b01010111000: data <= 32'hbe1e36d5;
    11'b01010111001: data <= 32'hbd7339f1;
    11'b01010111010: data <= 32'h2828b07c;
    11'b01010111011: data <= 32'h3edab6b3;
    11'b01010111100: data <= 32'h3ed439f2;
    11'b01010111101: data <= 32'ha4573fd5;
    11'b01010111110: data <= 32'hbca13f5a;
    11'b01010111111: data <= 32'hb4993b17;
    11'b01011000000: data <= 32'h3c7a32e2;
    11'b01011000001: data <= 32'h3c0fb4da;
    11'b01011000010: data <= 32'haf24bcff;
    11'b01011000011: data <= 32'hb09fbfae;
    11'b01011000100: data <= 32'h3d0abc8a;
    11'b01011000101: data <= 32'h403b3807;
    11'b01011000110: data <= 32'h3c6c3b9f;
    11'b01011000111: data <= 32'hb910b539;
    11'b01011001000: data <= 32'hbdc4bda9;
    11'b01011001001: data <= 32'hbd84ba46;
    11'b01011001010: data <= 32'hbd7635f3;
    11'b01011001011: data <= 32'hbd002a85;
    11'b01011001100: data <= 32'hb551bd4b;
    11'b01011001101: data <= 32'h3a48bdbb;
    11'b01011001110: data <= 32'h394c36dd;
    11'b01011001111: data <= 32'hb8d3408e;
    11'b01011010000: data <= 32'hbcb0409a;
    11'b01011010001: data <= 32'hb2ed3c91;
    11'b01011010010: data <= 32'h39aa3661;
    11'b01011010011: data <= 32'h2f073288;
    11'b01011010100: data <= 32'hbb4db468;
    11'b01011010101: data <= 32'hb359babb;
    11'b01011010110: data <= 32'h3fabb81b;
    11'b01011010111: data <= 32'h41fb377b;
    11'b01011011000: data <= 32'h3ed9392a;
    11'b01011011001: data <= 32'hb46fb4f7;
    11'b01011011010: data <= 32'hbb94bb49;
    11'b01011011011: data <= 32'hb835b43e;
    11'b01011011100: data <= 32'hb6e33432;
    11'b01011011101: data <= 32'hba2bbaac;
    11'b01011011110: data <= 32'hb876c0fa;
    11'b01011011111: data <= 32'h31a2c08a;
    11'b01011100000: data <= 32'h34442a3f;
    11'b01011100001: data <= 32'hb80e3feb;
    11'b01011100010: data <= 32'hbb623efe;
    11'b01011100011: data <= 32'hb6f237e7;
    11'b01011100100: data <= 32'hb3533140;
    11'b01011100101: data <= 32'hbc933973;
    11'b01011100110: data <= 32'hbf433920;
    11'b01011100111: data <= 32'hb80cae35;
    11'b01011101000: data <= 32'h3fcdb4d3;
    11'b01011101001: data <= 32'h41c33618;
    11'b01011101010: data <= 32'h3dc93ac0;
    11'b01011101011: data <= 32'hb40b37fa;
    11'b01011101100: data <= 32'hb44b32e7;
    11'b01011101101: data <= 32'h38e63838;
    11'b01011101110: data <= 32'h385c3575;
    11'b01011101111: data <= 32'hb682bcf7;
    11'b01011110000: data <= 32'hb935c1ba;
    11'b01011110001: data <= 32'h325dc0d2;
    11'b01011110010: data <= 32'h3a63b1e9;
    11'b01011110011: data <= 32'h356d3cf1;
    11'b01011110100: data <= 32'hb5e03880;
    11'b01011110101: data <= 32'hb8cab862;
    11'b01011110110: data <= 32'hbbc0b259;
    11'b01011110111: data <= 32'hbfb23b82;
    11'b01011111000: data <= 32'hc0943b83;
    11'b01011111001: data <= 32'hbad0b3e7;
    11'b01011111010: data <= 32'h3d3cba73;
    11'b01011111011: data <= 32'h3f762d9b;
    11'b01011111100: data <= 32'h383e3ce6;
    11'b01011111101: data <= 32'hb7cc3ddd;
    11'b01011111110: data <= 32'h33963cf6;
    11'b01011111111: data <= 32'h3d373cb1;
    11'b01100000000: data <= 32'h3a90394d;
    11'b01100000001: data <= 32'hb8b6bac8;
    11'b01100000010: data <= 32'hba1bc065;
    11'b01100000011: data <= 32'h3968bf2a;
    11'b01100000100: data <= 32'h3f5fb150;
    11'b01100000101: data <= 32'h3db437cc;
    11'b01100000110: data <= 32'h3430b7a6;
    11'b01100000111: data <= 32'hb73fbcce;
    11'b01100001000: data <= 32'hbb6cb434;
    11'b01100001001: data <= 32'hbeca3c0a;
    11'b01100001010: data <= 32'hc019386c;
    11'b01100001011: data <= 32'hbc4ebcbb;
    11'b01100001100: data <= 32'h3640bf2c;
    11'b01100001101: data <= 32'h38f8b623;
    11'b01100001110: data <= 32'hb5b13d76;
    11'b01100001111: data <= 32'hb9653f55;
    11'b01100010000: data <= 32'h368b3dd1;
    11'b01100010001: data <= 32'h3cc53d21;
    11'b01100010010: data <= 32'h31b43c49;
    11'b01100010011: data <= 32'hbd672f9e;
    11'b01100010100: data <= 32'hbc16bb86;
    11'b01100010101: data <= 32'h3c75bb07;
    11'b01100010110: data <= 32'h4132a29c;
    11'b01100010111: data <= 32'h40042ebd;
    11'b01100011000: data <= 32'h38caba07;
    11'b01100011001: data <= 32'h9f4fbbcf;
    11'b01100011010: data <= 32'hac81325d;
    11'b01100011011: data <= 32'hb8dc3c50;
    11'b01100011100: data <= 32'hbd34ad6d;
    11'b01100011101: data <= 32'hbc6cc069;
    11'b01100011110: data <= 32'hb453c13e;
    11'b01100011111: data <= 32'hab29ba62;
    11'b01100100000: data <= 32'hb8723c3f;
    11'b01100100001: data <= 32'hb8103d0a;
    11'b01100100010: data <= 32'h35d43966;
    11'b01100100011: data <= 32'h382e3a7c;
    11'b01100100100: data <= 32'hbb4b3d6e;
    11'b01100100101: data <= 32'hc0833c46;
    11'b01100100110: data <= 32'hbd842cc2;
    11'b01100100111: data <= 32'h3c5cb5ae;
    11'b01100101000: data <= 32'h40e622d4;
    11'b01100101001: data <= 32'h3e8d309e;
    11'b01100101010: data <= 32'h36d8b343;
    11'b01100101011: data <= 32'h3804a873;
    11'b01100101100: data <= 32'h3c5d3bff;
    11'b01100101101: data <= 32'h38fd3d1c;
    11'b01100101110: data <= 32'hb8edb63b;
    11'b01100101111: data <= 32'hbc38c10d;
    11'b01100110000: data <= 32'hb62fc15f;
    11'b01100110001: data <= 32'h31debb14;
    11'b01100110010: data <= 32'h2d23374d;
    11'b01100110011: data <= 32'h2a712ad6;
    11'b01100110100: data <= 32'h3598b8d9;
    11'b01100110101: data <= 32'hac9d300a;
    11'b01100110110: data <= 32'hbe7f3dca;
    11'b01100110111: data <= 32'hc15e3def;
    11'b01100111000: data <= 32'hbe87331e;
    11'b01100111001: data <= 32'h3864b8f9;
    11'b01100111010: data <= 32'h3da3b440;
    11'b01100111011: data <= 32'h380435b7;
    11'b01100111100: data <= 32'haf9d3878;
    11'b01100111101: data <= 32'h3a9d3b43;
    11'b01100111110: data <= 32'h3f853e85;
    11'b01100111111: data <= 32'h3ccc3e41;
    11'b01101000000: data <= 32'hb841aadc;
    11'b01101000001: data <= 32'hbc82bf55;
    11'b01101000010: data <= 32'had46bf7c;
    11'b01101000011: data <= 32'h3c10b898;
    11'b01101000100: data <= 32'h3c44aef3;
    11'b01101000101: data <= 32'h3981bc48;
    11'b01101000110: data <= 32'h381fbe3f;
    11'b01101000111: data <= 32'ha9d7b35a;
    11'b01101001000: data <= 32'hbd7b3dcc;
    11'b01101001001: data <= 32'hc0913d10;
    11'b01101001010: data <= 32'hbe63b7a3;
    11'b01101001011: data <= 32'hb22abdf1;
    11'b01101001100: data <= 32'h2de2ba12;
    11'b01101001101: data <= 32'hb97b36e2;
    11'b01101001110: data <= 32'hb8f53b2c;
    11'b01101001111: data <= 32'h3b323c5d;
    11'b01101010000: data <= 32'h3fb63e77;
    11'b01101010001: data <= 32'h3a823f06;
    11'b01101010010: data <= 32'hbc933a08;
    11'b01101010011: data <= 32'hbda2b815;
    11'b01101010100: data <= 32'h3409b94d;
    11'b01101010101: data <= 32'h3eccadda;
    11'b01101010110: data <= 32'h3e75b5d7;
    11'b01101010111: data <= 32'h3b8bbdfb;
    11'b01101011000: data <= 32'h3a63be73;
    11'b01101011001: data <= 32'h396d2a95;
    11'b01101011010: data <= 32'hb3253e21;
    11'b01101011011: data <= 32'hbd033a0d;
    11'b01101011100: data <= 32'hbd2abd93;
    11'b01101011101: data <= 32'hb9a8c08b;
    11'b01101011110: data <= 32'hb9cfbc83;
    11'b01101011111: data <= 32'hbcba3374;
    11'b01101100000: data <= 32'hb95936cc;
    11'b01101100001: data <= 32'h3ad13436;
    11'b01101100010: data <= 32'h3d9d3b1b;
    11'b01101100011: data <= 32'hb0703edd;
    11'b01101100100: data <= 32'hbfff3e2d;
    11'b01101100101: data <= 32'hbf023917;
    11'b01101100110: data <= 32'h3480319e;
    11'b01101100111: data <= 32'h3e7931fd;
    11'b01101101000: data <= 32'h3ccfb4cc;
    11'b01101101001: data <= 32'h3865bc80;
    11'b01101101010: data <= 32'h3c05bab6;
    11'b01101101011: data <= 32'h3eb73a4d;
    11'b01101101100: data <= 32'h3c853ef7;
    11'b01101101101: data <= 32'hb3af3725;
    11'b01101101110: data <= 32'hbb9fbefe;
    11'b01101101111: data <= 32'hba27c09b;
    11'b01101110000: data <= 32'hb933bc21;
    11'b01101110001: data <= 32'hb9faaec9;
    11'b01101110010: data <= 32'hb253b908;
    11'b01101110011: data <= 32'h3ae5bc87;
    11'b01101110100: data <= 32'h3ac2b00f;
    11'b01101110101: data <= 32'hbad63df7;
    11'b01101110110: data <= 32'hc0ce3f82;
    11'b01101110111: data <= 32'hbf773b99;
    11'b01101111000: data <= 32'ha8b730a3;
    11'b01101111001: data <= 32'h39bb274e;
    11'b01101111010: data <= 32'ha8e3af4f;
    11'b01101111011: data <= 32'hb525b692;
    11'b01101111100: data <= 32'h3c012ce5;
    11'b01101111101: data <= 32'h40ba3d9c;
    11'b01101111110: data <= 32'h3f7d3fba;
    11'b01101111111: data <= 32'h2f3c38d8;
    11'b01110000000: data <= 32'hbaebbcb3;
    11'b01110000001: data <= 32'hb7babd95;
    11'b01110000010: data <= 32'h2d52b69d;
    11'b01110000011: data <= 32'h31bbb572;
    11'b01110000100: data <= 32'h36d3be8a;
    11'b01110000101: data <= 32'h3bcbc082;
    11'b01110000110: data <= 32'h39f0ba41;
    11'b01110000111: data <= 32'hb9a03d2a;
    11'b01110001000: data <= 32'hbfb43ea3;
    11'b01110001001: data <= 32'hbe3235f0;
    11'b01110001010: data <= 32'hb753b8fc;
    11'b01110001011: data <= 32'hb7a4b715;
    11'b01110001100: data <= 32'hbd92a59e;
    11'b01110001101: data <= 32'hbc962037;
    11'b01110001110: data <= 32'h3aa9357f;
    11'b01110001111: data <= 32'h40c83d56;
    11'b01110010000: data <= 32'h3e803f85;
    11'b01110010001: data <= 32'hb5d73c73;
    11'b01110010010: data <= 32'hbc6b25a5;
    11'b01110010011: data <= 32'hb0d4a58e;
    11'b01110010100: data <= 32'h3a70369a;
    11'b01110010101: data <= 32'h3a50b52b;
    11'b01110010110: data <= 32'h3931c00b;
    11'b01110010111: data <= 32'h3c3bc0eb;
    11'b01110011000: data <= 32'h3cc9b965;
    11'b01110011001: data <= 32'h351f3d38;
    11'b01110011010: data <= 32'hb9e73ca6;
    11'b01110011011: data <= 32'hbb21b85e;
    11'b01110011100: data <= 32'hb962bdca;
    11'b01110011101: data <= 32'hbcf7ba61;
    11'b01110011110: data <= 32'hc01fac4d;
    11'b01110011111: data <= 32'hbda5b36e;
    11'b01110100000: data <= 32'h3974b5d7;
    11'b01110100001: data <= 32'h3f853770;
    11'b01110100010: data <= 32'h39a03dfa;
    11'b01110100011: data <= 32'hbced3e5b;
    11'b01110100100: data <= 32'hbdc73c67;
    11'b01110100101: data <= 32'ha2ba3c04;
    11'b01110100110: data <= 32'h3b503b9d;
    11'b01110100111: data <= 32'h37d7af5b;
    11'b01110101000: data <= 32'h3064bea5;
    11'b01110101001: data <= 32'h3b83befc;
    11'b01110101010: data <= 32'h3f86296e;
    11'b01110101011: data <= 32'h3e623e0d;
    11'b01110101100: data <= 32'h37963a3e;
    11'b01110101101: data <= 32'hb408bc36;
    11'b01110101110: data <= 32'hb867be56;
    11'b01110101111: data <= 32'hbcacb8e0;
    11'b01110110000: data <= 32'hbedfaf2e;
    11'b01110110001: data <= 32'hbbfbbbd6;
    11'b01110110010: data <= 32'h3976beb3;
    11'b01110110011: data <= 32'h3d1cba08;
    11'b01110110100: data <= 32'hb0263b7e;
    11'b01110110101: data <= 32'hbeef3eca;
    11'b01110110110: data <= 32'hbdf93da1;
    11'b01110110111: data <= 32'hacd33c64;
    11'b01110111000: data <= 32'h34ca3b29;
    11'b01110111001: data <= 32'hb94a2e48;
    11'b01110111010: data <= 32'hbb78bb65;
    11'b01110111011: data <= 32'h38abb9fc;
    11'b01110111100: data <= 32'h409f39f7;
    11'b01110111101: data <= 32'h40a43ea9;
    11'b01110111110: data <= 32'h3bdb39ca;
    11'b01110111111: data <= 32'ha146b9f4;
    11'b01111000000: data <= 32'hb2a3ba28;
    11'b01111000001: data <= 32'hb6d33258;
    11'b01111000010: data <= 32'hb9f520d6;
    11'b01111000011: data <= 32'hb4cebed8;
    11'b01111000100: data <= 32'h3a3cc18b;
    11'b01111000101: data <= 32'h3c01be5d;
    11'b01111000110: data <= 32'hb2fd383f;
    11'b01111000111: data <= 32'hbd6c3d8c;
    11'b01111001000: data <= 32'hbc073a9f;
    11'b01111001001: data <= 32'hb0b93520;
    11'b01111001010: data <= 32'hb8e23606;
    11'b01111001011: data <= 32'hbff23220;
    11'b01111001100: data <= 32'hbfdcb5ec;
    11'b01111001101: data <= 32'h3132b444;
    11'b01111001110: data <= 32'h40693a48;
    11'b01111001111: data <= 32'h40263de2;
    11'b01111010000: data <= 32'h38443b34;
    11'b01111010001: data <= 32'hb4303155;
    11'b01111010010: data <= 32'h2ff43890;
    11'b01111010011: data <= 32'h36593cfd;
    11'b01111010100: data <= 32'h2a90351e;
    11'b01111010101: data <= 32'h28bbbfba;
    11'b01111010110: data <= 32'h3a0cc1f6;
    11'b01111010111: data <= 32'h3c9cbe36;
    11'b01111011000: data <= 32'h382b3817;
    11'b01111011001: data <= 32'hb2b63b09;
    11'b01111011010: data <= 32'haf7db146;
    11'b01111011011: data <= 32'ha8e9b948;
    11'b01111011100: data <= 32'hbcb7ae0d;
    11'b01111011101: data <= 32'hc1533307;
    11'b01111011110: data <= 32'hc0aeb577;
    11'b01111011111: data <= 32'hac87b997;
    11'b01111100000: data <= 32'h3ea9a780;
    11'b01111100001: data <= 32'h3c633adc;
    11'b01111100010: data <= 32'hb7513c20;
    11'b01111100011: data <= 32'hb9b03c1b;
    11'b01111100100: data <= 32'h34eb3e6f;
    11'b01111100101: data <= 32'h39e83fc2;
    11'b01111100110: data <= 32'h246f394e;
    11'b01111100111: data <= 32'hb674be10;
    11'b01111101000: data <= 32'h36d1c074;
    11'b01111101001: data <= 32'h3df1b9f8;
    11'b01111101010: data <= 32'h3e3c3a80;
    11'b01111101011: data <= 32'h3c113785;
    11'b01111101100: data <= 32'h39b6baf7;
    11'b01111101101: data <= 32'h345dbc31;
    11'b01111101110: data <= 32'hbc161cf2;
    11'b01111101111: data <= 32'hc09735bf;
    11'b01111110000: data <= 32'hbf82b9f8;
    11'b01111110001: data <= 32'h95f7bf09;
    11'b01111110010: data <= 32'h3c2ebd09;
    11'b01111110011: data <= 32'h2df62cfb;
    11'b01111110100: data <= 32'hbcc93b39;
    11'b01111110101: data <= 32'hbae93ce2;
    11'b01111110110: data <= 32'h36623eca;
    11'b01111110111: data <= 32'h37323f87;
    11'b01111111000: data <= 32'hbb063ac0;
    11'b01111111001: data <= 32'hbde9ba19;
    11'b01111111010: data <= 32'hb16abc57;
    11'b01111111011: data <= 32'h3e8c31a9;
    11'b01111111100: data <= 32'h404a3c54;
    11'b01111111101: data <= 32'h3e2634a9;
    11'b01111111110: data <= 32'h3c07baf0;
    11'b01111111111: data <= 32'h390ab7e3;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    