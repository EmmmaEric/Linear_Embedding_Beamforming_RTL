
    module interp_rom_0(
    CLK, rst,
    Addr, CEB, Q
    );

    input CLK, rst;
    input [9:0] Addr;
    input CEB;		
    output [20:0] Q;

    (*rom_style = "block" *) reg [20:0] data;

    always @(posedge CLK) begin
    if (rst) begin
        data <= 20'd0;
    end else begin
    if (CEB)
    case(Addr)
        10'b00000000: data <= 20'b11000011001100000010;
        10'b00000001: data <= 20'b11001011011100100001;
        10'b00000010: data <= 20'b01001100100100101001;
        10'b00000011: data <= 20'b01001000010100010110;
        10'b00000100: data <= 20'b01000110110100000001;
        10'b00000101: data <= 20'b01000001110011111100;
        10'b00000110: data <= 20'b10111010110100010001;
        10'b00000111: data <= 20'b11001100101100101111;
        10'b00001000: data <= 20'b01000000111100100111;
        10'b00001001: data <= 20'b01001011001100100111;
        10'b00001010: data <= 20'b01001000100100001100;
        10'b00001011: data <= 20'b01000011100100001010;
        10'b00001100: data <= 20'b00111110100100010001;
        10'b00001101: data <= 20'b10101111100100011010;
        10'b00001110: data <= 20'b11000000110100111111;
        10'b00001111: data <= 20'b01001000111100011011;
        10'b00010000: data <= 20'b01000101101100010000;
        10'b00010001: data <= 20'b01000101111011111110;
        10'b00010010: data <= 20'b00111001110011100001;
        10'b00010011: data <= 20'b11000101110100011000;
        10'b00010100: data <= 20'b10111100010100100011;
        10'b00010101: data <= 20'b00110111000100110001;
        10'b00010110: data <= 20'b01001010111011111100;
        10'b00010111: data <= 20'b01000100111011101101;
        10'b00011000: data <= 20'b00111101000011010101;
        10'b00011001: data <= 20'b11001001001100011101;
        10'b00011010: data <= 20'b00110101111100110100;
        10'b00011011: data <= 20'b11001001000101000011;
        10'b00011100: data <= 20'b00110000010100110011;
        10'b00011101: data <= 20'b01001100000100010000;
        10'b00011110: data <= 20'b01000100110011100011;
        10'b00011111: data <= 20'b00111000100100000000;
        10'b00100000: data <= 20'b11001010110100100101;
        10'b00100001: data <= 20'b01001011011100011011;
        10'b00100010: data <= 20'b01001010001100011000;
        10'b00100011: data <= 20'b01010001010100100010;
        10'b00100100: data <= 20'b01001101110100100010;
        10'b00100101: data <= 20'b01000100000011111010;
        10'b00100110: data <= 20'b10110011000100000110;
        10'b00100111: data <= 20'b11001000010100100000;
        10'b00101000: data <= 20'b01001100111011101111;
        10'b00101001: data <= 20'b01001000001011110001;
        10'b00101010: data <= 20'b01000110011011110111;
        10'b00101011: data <= 20'b01000100011100000101;
        10'b00101100: data <= 20'b00100101010100010011;
        10'b00101101: data <= 20'b11000001110100001011;
        10'b00101110: data <= 20'b11001000110100010100;
        10'b00101111: data <= 20'b01001111110011100100;
        10'b00110000: data <= 20'b01000111100011001100;
        10'b00110001: data <= 20'b01000010110011101110;
        10'b00110010: data <= 20'b10111000000100010111;
        10'b00110011: data <= 20'b01001000100100100110;
        10'b00110100: data <= 20'b11001110100100111101;
        10'b00110101: data <= 20'b11001011001100001011;
        10'b00110110: data <= 20'b01001010001101000011;
        10'b00110111: data <= 20'b01000111110010010011;
        10'b00111000: data <= 20'b01000000110011110101;
        10'b00111001: data <= 20'b11000010110100010101;
        10'b00111010: data <= 20'b01001001010100101000;
        10'b00111011: data <= 20'b01001010110100011000;
        10'b00111100: data <= 20'b01001010101100110000;
        10'b00111101: data <= 20'b01000001011100100011;
        10'b00111110: data <= 20'b01000110011100000011;
        10'b00111111: data <= 20'b00111100100011101101;
        10'b01000000: data <= 20'b11000101010100000010;
        10'b01000001: data <= 20'b01001011010100111000;
        10'b01000010: data <= 20'b01001001000100010011;
        10'b01000011: data <= 20'b01001000110011111000;
        10'b01000100: data <= 20'b01000100101011111011;
        10'b01000101: data <= 20'b00111110010011011101;
        10'b01000110: data <= 20'b11000001110010100011;
        10'b01000111: data <= 20'b11000110011100001000;
        10'b01001000: data <= 20'b11010000011101010100;
        10'b01001001: data <= 20'b01001001110100010000;
        10'b01001010: data <= 20'b01000110010100000110;
        10'b01001011: data <= 20'b01000011100100000100;
        10'b01001100: data <= 20'b00111110100100010000;
        10'b01001101: data <= 20'b11000101000100100110;
        10'b01001110: data <= 20'b11000000101100101110;
        10'b01001111: data <= 20'b01000010001100101000;
        10'b01010000: data <= 20'b01001010011100000011;
        10'b01010001: data <= 20'b01000100110100000000;
        10'b01010010: data <= 20'b00110110000100001101;
        10'b01010011: data <= 20'b00111100010100011101;
        10'b01010100: data <= 20'b00111101100100100110;
        10'b01010101: data <= 20'b01001111001100011011;
        10'b01010110: data <= 20'b01000110001100010100;
        10'b01010111: data <= 20'b01000100101100001011;
        10'b01011000: data <= 20'b01000001111011011000;
        10'b01011001: data <= 20'b11000010101011010001;
        10'b01011010: data <= 20'b11000110010100101100;
        10'b01011011: data <= 20'b01000010000100101000;
        10'b01011100: data <= 20'b01001011100100101000;
        10'b01011101: data <= 20'b01000111011011110111;
        10'b01011110: data <= 20'b01000001101010100111;
        10'b01011111: data <= 20'b11000001010011110001;
        10'b01100000: data <= 20'b11000001111100100111;
        10'b01100001: data <= 20'b10110111111100111010;
        10'b01100010: data <= 20'b01001010000100110101;
        10'b01100011: data <= 20'b01001000110100101000;
        10'b01100100: data <= 20'b01000111110011110110;
        10'b01100101: data <= 20'b01000000110011111011;
        10'b01100110: data <= 20'b11000000110100010001;
        10'b01100111: data <= 20'b01010000101101000111;
        10'b01101000: data <= 20'b01001000101100011010;
        10'b01101001: data <= 20'b01001010001100011010;
        10'b01101010: data <= 20'b01001010100100100001;
        10'b01101011: data <= 20'b01000110010100001111;
        10'b01101100: data <= 20'b00111101010100001001;
        10'b01101101: data <= 20'b11000001000100010100;
        10'b01101110: data <= 20'b11000000000101001011;
        10'b01101111: data <= 20'b01001001001100000011;
        10'b01110000: data <= 20'b01000101111011110110;
        10'b01110001: data <= 20'b01000011101011110001;
        10'b01110010: data <= 20'b11001010111011010000;
        10'b01110011: data <= 20'b11000101000100011100;
        10'b01110100: data <= 20'b11000101000100011000;
        10'b01110101: data <= 20'b11001100110100110110;
        10'b01110110: data <= 20'b01001010001011101100;
        10'b01110111: data <= 20'b01000100100011010001;
        10'b01111000: data <= 20'b00111000100011111011;
        10'b01111001: data <= 20'b01000111000100111010;
        10'b01111010: data <= 20'b01001101110100001010;
        10'b01111011: data <= 20'b11010000110100101000;
        10'b01111100: data <= 20'b11001110111011110111;
        10'b01111101: data <= 20'b01001011111100001100;
        10'b01111110: data <= 20'b01000100010011101001;
        10'b01111111: data <= 20'b10110101010100000001;
        10'b10000000: data <= 20'b11000111010100110100;
        10'b10000001: data <= 20'b01001010110100001101;
        10'b10000010: data <= 20'b01001010111011010011;
        10'b10000011: data <= 20'b01000101111100101101;
        10'b10000100: data <= 20'b01000101101100100000;
        10'b10000101: data <= 20'b01000010010011100010;
        10'b10000110: data <= 20'b10111110010011111010;
        10'b10000111: data <= 20'b11001011100100100000;
        10'b10001000: data <= 20'b01001011110100010011;
        10'b10001001: data <= 20'b01001000000011111101;
        10'b10001010: data <= 20'b01000110101001100101;
        10'b10001011: data <= 20'b01000001100011011111;
        10'b10001100: data <= 20'b10111011000100001100;
        10'b10001101: data <= 20'b11000101011011011010;
        10'b10001110: data <= 20'b11001010001100010100;
        10'b10001111: data <= 20'b01001110001011110010;
        10'b10010000: data <= 20'b01000111010011111110;
        10'b10010001: data <= 20'b01000011000100000001;
        10'b10010010: data <= 20'b01000000000100010100;
        10'b10010011: data <= 20'b01000000010100100000;
        10'b10010100: data <= 20'b11010011000100111010;
        10'b10010101: data <= 20'b10111100101100101000;
        10'b10010110: data <= 20'b01000111111100101000;
        10'b10010111: data <= 20'b01000111010011011010;
        10'b10011000: data <= 20'b00111110110011111011;
        10'b10011001: data <= 20'b11000001010100011100;
        10'b10011010: data <= 20'b01000011110100100100;
        10'b10011011: data <= 20'b01001001000100101011;
        10'b10011100: data <= 20'b01001001011100011101;
        10'b10011101: data <= 20'b01000100001100001111;
        10'b10011110: data <= 20'b01000011011011111111;
        10'b10011111: data <= 20'b10110011101011011000;
        10'b10100000: data <= 20'b11001000110010110011;
        10'b10100001: data <= 20'b01000110000100110011;
        10'b10100010: data <= 20'b01001000000100100011;
        10'b10100011: data <= 20'b01001001110011111110;
        10'b10100100: data <= 20'b01000100011011011000;
        10'b10100101: data <= 20'b00111010000011110101;
        10'b10100110: data <= 20'b11001000011100001010;
        10'b10100111: data <= 20'b11000000011100100111;
        10'b10101000: data <= 20'b01001111011101000001;
        10'b10101001: data <= 20'b01001001100100100001;
        10'b10101010: data <= 20'b01000111110100010100;
        10'b10101011: data <= 20'b01000100000100000000;
        10'b10101100: data <= 20'b00111000110100001011;
        10'b10101101: data <= 20'b11001000100100100111;
        10'b10101110: data <= 20'b01001001011100100111;
        10'b10101111: data <= 20'b01000111011100011010;
        10'b10110000: data <= 20'b01001010001100000011;
        10'b10110001: data <= 20'b01000101010100001110;
        10'b10110010: data <= 20'b00111100110100010000;
        10'b10110011: data <= 20'b10110101010100010101;
        10'b10110100: data <= 20'b11000100010100100110;
        10'b10110101: data <= 20'b01001101011100001101;
        10'b10110110: data <= 20'b01000110101100000001;
        10'b10110111: data <= 20'b01000011101011110011;
        10'b10111000: data <= 20'b10111011011011110110;
        10'b10111001: data <= 20'b11001010011100011111;
        10'b10111010: data <= 20'b11000110010100100101;
        10'b10111011: data <= 20'b11000101100100100111;
        10'b10111100: data <= 20'b01001111010100101001;
        10'b10111101: data <= 20'b01000110111011011001;
        10'b10111110: data <= 20'b01000000110011101001;
        10'b10111111: data <= 20'b11000101000100010001;
        10'b11000000: data <= 20'b01001101111100100000;
        10'b11000001: data <= 20'b01001110001100100111;
        10'b11000010: data <= 20'b11001111000101000000;
        10'b11000011: data <= 20'b01010011110101010011;
        10'b11000100: data <= 20'b01000111010011001111;
        10'b11000101: data <= 20'b00111111000011111001;
        10'b11000110: data <= 20'b11000100010100010010;
        10'b11000111: data <= 20'b01001111000100100000;
        10'b11001000: data <= 20'b01001001101011101001;
        10'b11001001: data <= 20'b01001001111100001110;
        10'b11001010: data <= 20'b01000101001100110000;
        10'b11001011: data <= 20'b01000110001011101111;
        10'b11001100: data <= 20'b00110100110011111110;
        10'b11001101: data <= 20'b11000101000100001001;
        10'b11001110: data <= 20'b01010001100101001011;
        10'b11001111: data <= 20'b01001001000011101001;
        10'b11010000: data <= 20'b01000110000011100011;
        10'b11010001: data <= 20'b01000010110011110000;
        10'b11010010: data <= 20'b01000001000100010011;
        10'b11010011: data <= 20'b11000110010100010100;
        10'b11010100: data <= 20'b11001000001011000000;
        10'b11010101: data <= 20'b11010000011100111100;
        10'b11010110: data <= 20'b01001001100011010011;
        10'b11010111: data <= 20'b01000100100011110100;
        10'b11011000: data <= 20'b00111000000100001010;
        10'b11011001: data <= 20'b01000011100100100010;
        10'b11011010: data <= 20'b01001000010100101011;
        10'b11011011: data <= 20'b11001000001100111100;
        10'b11011100: data <= 20'b10111010011100101010;
        10'b11011101: data <= 20'b01001001001100010011;
        10'b11011110: data <= 20'b01000011010011101101;
        10'b11011111: data <= 20'b10111110010100000010;
        10'b11100000: data <= 20'b00110011000100110000;
        10'b11100001: data <= 20'b01001000100100100010;
        10'b11100010: data <= 20'b01001100000100001100;
        10'b11100011: data <= 20'b01000101111100010101;
        10'b11100100: data <= 20'b01000010101100000111;
        10'b11100101: data <= 20'b00111101101011010111;
        10'b11100110: data <= 20'b11000010101011100011;
        10'b11100111: data <= 20'b11001111000100100010;
        10'b11101000: data <= 20'b01001010000100100010;
        10'b11101001: data <= 20'b01001000100100010100;
        10'b11101010: data <= 20'b01000110110011010100;
        10'b11101011: data <= 20'b01000001000011110010;
        10'b11101100: data <= 20'b11000001010100001100;
        10'b11101101: data <= 20'b11000110001100100001;
        10'b11101110: data <= 20'b11000000111100101101;
        10'b11101111: data <= 20'b01001101100011010110;
        10'b11110000: data <= 20'b01000111100100010000;
        10'b11110001: data <= 20'b01000100010100001001;
        10'b11110010: data <= 20'b01000000000100001110;
        10'b11110011: data <= 20'b10111010000100011011;
        10'b11110100: data <= 20'b01011000111101101010;
        10'b11110101: data <= 20'b01000110101100011111;
        10'b11110110: data <= 20'b01000111001100011000;
        10'b11110111: data <= 20'b01000111010011101001;
        10'b11111000: data <= 20'b00111011010100000001;
        10'b11111001: data <= 20'b10111100110100011011;
        10'b11111010: data <= 20'b10110101110100100001;
        10'b11111011: data <= 20'b01000110110100111000;
        10'b11111100: data <= 20'b01001000111100001011;
        10'b11111101: data <= 20'b01000100011011111001;
        10'b11111110: data <= 20'b00111101111011101000;
        10'b11111111: data <= 20'b11000010101100010011;
        10'b100000000: data <= 20'b11001101011100011101;
        10'b100000001: data <= 20'b11000000100100101111;
        10'b100000010: data <= 20'b01000001110100110010;
        10'b100000011: data <= 20'b01001010000011010011;
        10'b100000100: data <= 20'b01000100000011010101;
        10'b100000101: data <= 20'b10101101110011111111;
        10'b100000110: data <= 20'b11010001111100011010;
        10'b100000111: data <= 20'b01001001111100100100;
        10'b100001000: data <= 20'b01001111001100101100;
        10'b100001001: data <= 20'b01001000000100111011;
        10'b100001010: data <= 20'b01001011010100010000;
        10'b100001011: data <= 20'b01000011010011111000;
        10'b100001100: data <= 20'b10111000010100000111;
        10'b100001101: data <= 20'b11001011000100110000;
        10'b100001110: data <= 20'b01001011001100000111;
        10'b100001111: data <= 20'b01001000001100000010;
        10'b100010000: data <= 20'b01001001011100010001;
        10'b100010001: data <= 20'b01001100011100001101;
        10'b100010010: data <= 20'b00111110000100000110;
        10'b100010011: data <= 20'b11000000000100001011;
        10'b100010100: data <= 20'b11001001110100100001;
        10'b100010101: data <= 20'b01001100011011010110;
        10'b100010110: data <= 20'b01000110111010110100;
        10'b100010111: data <= 20'b01000011000011100000;
        10'b100011000: data <= 20'b00111011100100011100;
        10'b100011001: data <= 20'b01000110100100110010;
        10'b100011010: data <= 20'b11001000110100010011;
        10'b100011011: data <= 20'b11001011000011111010;
        10'b100011100: data <= 20'b01001111001100011111;
        10'b100011101: data <= 20'b01000110100011011110;
        10'b100011110: data <= 20'b01000000000011111000;
        10'b100011111: data <= 20'b11000010010100100001;
        10'b100100000: data <= 20'b01001001110100100011;
        10'b100100001: data <= 20'b01001110000100011110;
        10'b100100010: data <= 20'b11000110001100110011;
        10'b100100011: data <= 20'b01000100111100101111;
        10'b100100100: data <= 20'b01000110011011011000;
        10'b100100101: data <= 20'b00111011100011110101;
        10'b100100110: data <= 20'b11000110100100010101;
        10'b100100111: data <= 20'b01001010110100101000;
        10'b100101000: data <= 20'b01001001010100010001;
        10'b100101001: data <= 20'b01001001101100000100;
        10'b100101010: data <= 20'b01000011011100001100;
        10'b100101011: data <= 20'b01000000101011101110;
        10'b100101100: data <= 20'b10111101000011001110;
        10'b100101101: data <= 20'b11001000001011100110;
        10'b100101110: data <= 20'b01010000110100111001;
        10'b100101111: data <= 20'b01001000110100001111;
        10'b100110000: data <= 20'b01000110100100000011;
        10'b100110001: data <= 20'b01000011100011110110;
        10'b100110010: data <= 20'b00111100100100001101;
        10'b100110011: data <= 20'b11001001110100001010;
        10'b100110100: data <= 20'b11000101001100100011;
        10'b100110101: data <= 20'b01000101011100110110;
        10'b100110110: data <= 20'b01001001100011111100;
        10'b100110111: data <= 20'b01000100100100000011;
        10'b100111000: data <= 20'b00111101110100010001;
        10'b100111001: data <= 20'b00111110010100011010;
        10'b100111010: data <= 20'b00110110110100101101;
        10'b100111011: data <= 20'b01001001101100101110;
        10'b100111100: data <= 20'b01000100111100011011;
        10'b100111101: data <= 20'b01000111011100001110;
        10'b100111110: data <= 20'b01000010000011101100;
        10'b100111111: data <= 20'b11000010110100000101;
        10'b101000000: data <= 20'b10101101110100100110;
        10'b101000001: data <= 20'b01000010110100101000;
        10'b101000010: data <= 20'b01001100110100001010;
        10'b101000011: data <= 20'b01000101111100000010;
        10'b101000100: data <= 20'b01000001011011101011;
        10'b101000101: data <= 20'b10111111101011110101;
        10'b101000110: data <= 20'b11000100111100011011;
        10'b101000111: data <= 20'b11010011010100111010;
        10'b101001000: data <= 20'b01000110010100101101;
        10'b101001001: data <= 20'b01001010000100100011;
        10'b101001010: data <= 20'b01000110100011010011;
        10'b101001011: data <= 20'b01000000000011110111;
        10'b101001100: data <= 20'b11000100110100010001;
        10'b101001101: data <= 20'b01001000011100110011;
        10'b101001110: data <= 20'b01001000011100100101;
        10'b101001111: data <= 20'b01001110010011110110;
        10'b101010000: data <= 20'b01001000110100100011;
        10'b101010001: data <= 20'b01000101110100000101;
        10'b101010010: data <= 20'b00111101010100000111;
        10'b101010011: data <= 20'b11000010100100011000;
        10'b101010100: data <= 20'b01010001111100001010;
        10'b101010101: data <= 20'b01001000011100001011;
        10'b101010110: data <= 20'b01000110101100000110;
        10'b101010111: data <= 20'b01001000011011001100;
        10'b101011000: data <= 20'b10110100100100001110;
        10'b101011001: data <= 20'b10111101010100010011;
        10'b101011010: data <= 20'b11000100010100011001;
        10'b101011011: data <= 20'b01001000110101001100;
        10'b101011100: data <= 20'b01001000101011110010;
        10'b101011101: data <= 20'b01000100011010110101;
        10'b101011110: data <= 20'b00100001010011111001;
        10'b101011111: data <= 20'b01010000110100110100;
        10'b101100000: data <= 20'b11001010110101011001;
        10'b101100001: data <= 20'b11001010000100100000;
        10'b101100010: data <= 20'b11010000110100110101;
        10'b101100011: data <= 20'b01001001101011101000;
        10'b101100100: data <= 20'b01000011010011101011;
        10'b101100101: data <= 20'b10111100000100000101;
        10'b101100110: data <= 20'b01001001110100111011;
        10'b101100111: data <= 20'b01001011010011111101;
        10'b101101000: data <= 20'b01001110011100100100;
        10'b101101001: data <= 20'b11001000001100110110;
        10'b101101010: data <= 20'b01001001101100010110;
        10'b101101011: data <= 20'b01000001110011110000;
        10'b101101100: data <= 20'b10111111110100000010;
        10'b101101101: data <= 20'b11001011000100111011;
        10'b101101110: data <= 20'b01001010010100001000;
        10'b101101111: data <= 20'b01001000100011101101;
        10'b101110000: data <= 20'b01000110111100001011;
        10'b101110001: data <= 20'b01000001011011111000;
        10'b101110010: data <= 20'b10101110010011110101;
        10'b101110011: data <= 20'b11000100000011100110;
        10'b101110100: data <= 20'b11001101011011100010;
        10'b101110101: data <= 20'b01001011110100000110;
        10'b101110110: data <= 20'b01000110110011111100;
        10'b101110111: data <= 20'b01000011110011111111;
        10'b101111000: data <= 20'b01000001000100010000;
        10'b101111001: data <= 20'b00110010100100100010;
        10'b101111010: data <= 20'b11001010111100011011;
        10'b101111011: data <= 20'b11000110011100101000;
        10'b101111100: data <= 20'b01001100001100100001;
        10'b101111101: data <= 20'b01000110010011110101;
        10'b101111110: data <= 20'b00111110010100000010;
        10'b101111111: data <= 20'b00110010000100100000;
        10'b110000000: data <= 20'b01000100000100100011;
        10'b110000001: data <= 20'b01001110010100110011;
        10'b110000010: data <= 20'b01000101101100100010;
        10'b110000011: data <= 20'b01000100101100011000;
        10'b110000100: data <= 20'b01000101001011101000;
        10'b110000101: data <= 20'b10110011000011100110;
        10'b110000110: data <= 20'b11001000100100011101;
        10'b110000111: data <= 20'b01000110010100101001;
        10'b110001000: data <= 20'b01001000110100100011;
        10'b110001001: data <= 20'b01001001001100000000;
        10'b110001010: data <= 20'b01000011101011110011;
        10'b110001011: data <= 20'b00110110110011001100;
        10'b110001100: data <= 20'b11000011101100001100;
        10'b110001101: data <= 20'b11001000011100100100;
        10'b110001110: data <= 20'b01001110100100111001;
        10'b110001111: data <= 20'b01001000100100100000;
        10'b110010000: data <= 20'b01001000010100001011;
        10'b110010001: data <= 20'b01000011010011110110;
        10'b110010010: data <= 20'b10011111100100001011;
        10'b110010011: data <= 20'b11001110100100001100;
        10'b110010100: data <= 20'b01000101111100100110;
        10'b110010101: data <= 20'b01001000111100100101;
        10'b110010110: data <= 20'b01001010010100010000;
        10'b110010111: data <= 20'b01000101010100010001;
        10'b110011000: data <= 20'b01000000100100001101;
        10'b110011001: data <= 20'b10110010100100010100;
        10'b110011010: data <= 20'b11000110100100110000;
        10'b110011011: data <= 20'b01001010101100011001;
        10'b110011100: data <= 20'b01000110001100001001;
        10'b110011101: data <= 20'b01000101011100000010;
        10'b110011110: data <= 20'b00111110110011010100;
        10'b110011111: data <= 20'b11000110010100010010;
        10'b110100000: data <= 20'b11000000110100011111;
        10'b110100001: data <= 20'b11000100110100101011;
        10'b110100010: data <= 20'b01001100111010100011;
        10'b110100011: data <= 20'b01000101111011100111;
        10'b110100100: data <= 20'b01000000010011011100;
        10'b110100101: data <= 20'b11001001010100000110;
        10'b110100110: data <= 20'b01001011101100110011;
        10'b110100111: data <= 20'b11010010100101010010;
        10'b110101000: data <= 20'b11001000110100110001;
        10'b110101001: data <= 20'b01001111100100100011;
        10'b110101010: data <= 20'b01000101110011011000;
        10'b110101011: data <= 20'b00111101100011111010;
        10'b110101100: data <= 20'b11000110110100011011;
        10'b110101101: data <= 20'b01001101001011110011;
        10'b110101110: data <= 20'b01001010001100000111;
        10'b110101111: data <= 20'b01001110101100110001;
        10'b110110000: data <= 20'b01001110001101000101;
        10'b110110001: data <= 20'b01000101100011100010;
        10'b110110010: data <= 20'b00110110000100000000;
        10'b110110011: data <= 20'b11000110010100010011;
        10'b110110100: data <= 20'b01001110110100011011;
        10'b110110101: data <= 20'b01001000100011000011;
        10'b110110110: data <= 20'b01000110101011011100;
        10'b110110111: data <= 20'b01000011101011111011;
        10'b110111000: data <= 20'b00111110110100001001;
        10'b110111001: data <= 20'b11000001110100000011;
        10'b110111010: data <= 20'b11001000000011111111;
        10'b110111011: data <= 20'b01010110101100100011;
        10'b110111100: data <= 20'b01001000100011101000;
        10'b110111101: data <= 20'b01000100010011110011;
        10'b110111110: data <= 20'b00111011100100010000;
        10'b110111111: data <= 20'b01000100100100100001;
        10'b111000000: data <= 20'b10111101000100111011;
        10'b111000001: data <= 20'b11001001111100100001;
        10'b111000010: data <= 20'b11000010111100110101;
        10'b111000011: data <= 20'b01001000111011101101;
        10'b111000100: data <= 20'b01000010100011110100;
        10'b111000101: data <= 20'b10111111100100001110;
        10'b111000110: data <= 20'b01000101000100101010;
        10'b111000111: data <= 20'b01001001000100100010;
        10'b111001000: data <= 20'b01001100111100100010;
        10'b111001001: data <= 20'b01000011101100011101;
        10'b111001010: data <= 20'b01000101011100010000;
        10'b111001011: data <= 20'b00111111100011011000;
        10'b111001100: data <= 20'b11000011110011110000;
        10'b111001101: data <= 20'b11000010100100111101;
        10'b111001110: data <= 20'b01001001000100011111;
        10'b111001111: data <= 20'b01001001010100001110;
        10'b111010000: data <= 20'b01000101111011110111;
        10'b111010001: data <= 20'b01000000000011010001;
        10'b111010010: data <= 20'b11000010010011100010;
        10'b111010011: data <= 20'b11000101001100010011;
        10'b111010100: data <= 20'b11001011111100111010;
        10'b111010101: data <= 20'b01001011010100011010;
        10'b111010110: data <= 20'b01000111010100010000;
        10'b111010111: data <= 20'b01000100110100000011;
        10'b111011000: data <= 20'b00111111100100001001;
        10'b111011001: data <= 20'b11000001010100011110;
        10'b111011010: data <= 20'b00110011001100110111;
        10'b111011011: data <= 20'b01000100101100100100;
        10'b111011100: data <= 20'b01001010011100011001;
        10'b111011101: data <= 20'b01000110010100000100;
        10'b111011110: data <= 20'b00111101110100001010;
        10'b111011111: data <= 20'b00111001000100011000;
        10'b111100000: data <= 20'b10110110100100100010;
        10'b111100001: data <= 20'b01010000100100110101;
        10'b111100010: data <= 20'b01000111101100010010;
        10'b111100011: data <= 20'b01000100101100000101;
        10'b111100100: data <= 20'b01000010101011110010;
        10'b111100101: data <= 20'b11000001001011110110;
        10'b111100110: data <= 20'b11001000110100100101;
        10'b111100111: data <= 20'b10110111000100101000;
        10'b111101000: data <= 20'b01001000100100110100;
        10'b111101001: data <= 20'b01001000101011110011;
        10'b111101010: data <= 20'b01000011001010100101;
        10'b111101011: data <= 20'b10111100000011111000;
        10'b111101100: data <= 20'b11000100111100110101;
        10'b111101101: data <= 20'b01001000001100110011;
        10'b111101110: data <= 20'b01001010010101000101;
        10'b111101111: data <= 20'b01000110010100110100;
        10'b111110000: data <= 20'b01001001010011111000;
        10'b111110001: data <= 20'b01000010010011110101;
        10'b111110010: data <= 20'b10111100110100001001;
        10'b111110011: data <= 20'b11010001000101010011;
        10'b111110100: data <= 20'b01001001111100010010;
        10'b111110101: data <= 20'b01001001011100010011;
        10'b111110110: data <= 20'b01001111010100001111;
        10'b111110111: data <= 20'b01001010000100001011;
        10'b111111000: data <= 20'b01000000000100000011;
        10'b111111001: data <= 20'b10111111110100001110;
        10'b111111010: data <= 20'b11001100000100110011;
        10'b111111011: data <= 20'b01001010011011110100;
        10'b111111100: data <= 20'b01000110101011100101;
        10'b111111101: data <= 20'b01000100001011011111;
        10'b111111110: data <= 20'b01000000110100011010;
        10'b111111111: data <= 20'b11000100100100100000;
        10'b1000000000: data <= 20'b11000101010100010000;
        10'b1000000001: data <= 20'b11001100010100011100;
        10'b1000000010: data <= 20'b01001100001011110000;
        10'b1000000011: data <= 20'b01000101110011011110;
        10'b1000000100: data <= 20'b00111110110011111001;
        10'b1000000101: data <= 20'b10110000100100101001;
        10'b1000000110: data <= 20'b01001011000100100011;
        10'b1000000111: data <= 20'b11010111100100110010;
        10'b1000001000: data <= 20'b11001011101100100100;
        10'b1000001001: data <= 20'b01001100011100101010;
        10'b1000001010: data <= 20'b01000101010011100000;
        10'b1000001011: data <= 20'b00111000110011111011;
        10'b1000001100: data <= 20'b11000110110100100101;
        10'b1000001101: data <= 20'b01001010010100100000;
        10'b1000001110: data <= 20'b01001010100100001011;
        10'b1000001111: data <= 20'b01001000011100100100;
        10'b1000010000: data <= 20'b01000010111100011001;
        10'b1000010001: data <= 20'b01000011101011100010;
        10'b1000010010: data <= 20'b10111011000011101100;
        10'b1000010011: data <= 20'b11001001010100000111;
        10'b1000010100: data <= 20'b01001100100100100110;
        10'b1000010101: data <= 20'b01001000100100001011;
        10'b1000010110: data <= 20'b01000111100011101111;
        10'b1000010111: data <= 20'b01000010110011000111;
        10'b1000011000: data <= 20'b00110010000100000110;
        10'b1000011001: data <= 20'b11000110001011110110;
        10'b1000011010: data <= 20'b11001000001100011011;
        10'b1000011011: data <= 20'b01010000101100110010;
        10'b1000011100: data <= 20'b01001000100100000110;
        10'b1000011101: data <= 20'b01000100100100000100;
        10'b1000011110: data <= 20'b01000000110100001111;
        10'b1000011111: data <= 20'b00111101100100011001;
        10'b1000100000: data <= 20'b11001001000100111001;
        10'b1000100001: data <= 20'b01000001011100101010;
        10'b1000100010: data <= 20'b01000101011100100100;
        10'b1000100011: data <= 20'b01001000101011101000;
        10'b1000100100: data <= 20'b01000001100011111011;
        10'b1000100101: data <= 20'b11000000010100010100;
        10'b1000100110: data <= 20'b00111110010100100010;
        10'b1000100111: data <= 20'b01000100100100101100;
        10'b1000101000: data <= 20'b01001011101100010111;
        10'b1000101001: data <= 20'b01000101001100001010;
        10'b1000101010: data <= 20'b01000010011100000000;
        10'b1000101011: data <= 20'b00110001101011110000;
        10'b1000101100: data <= 20'b11000111011100000011;
        10'b1000101101: data <= 20'b10111111110100110101;
        10'b1000101110: data <= 20'b01000101110100101001;
        10'b1000101111: data <= 20'b01001011000100010101;
        10'b1000110000: data <= 20'b01000101011011011011;
        10'b1000110001: data <= 20'b00111110000011110000;
        10'b1000110010: data <= 20'b11001000010011110111;
        10'b1000110011: data <= 20'b00111110111100101011;
        10'b1000110100: data <= 20'b01001010011100110111;
        10'b1000110101: data <= 20'b01001011000100101101;
        10'b1000110110: data <= 20'b01001000110100100000;
        10'b1000110111: data <= 20'b01000101010011111011;
        10'b1000111000: data <= 20'b00111100010100000101;
        10'b1000111001: data <= 20'b11000101100100011101;
        10'b1000111010: data <= 20'b01001100111100101000;
        10'b1000111011: data <= 20'b01001000001100010011;
        10'b1000111100: data <= 20'b01001001001100010001;
        10'b1000111101: data <= 20'b01001000010100010110;
        10'b1000111110: data <= 20'b01000001000100001110;
        10'b1000111111: data <= 20'b10110011100100010001;
        10'b1001000000: data <= 20'b11000100100100011110;
        10'b1001000001: data <= 20'b01010000100100011000;
        10'b1001000010: data <= 20'b01001000001011111001;
        10'b1001000011: data <= 20'b01000100011011100111;
        10'b1001000100: data <= 20'b10110100110011100010;
        10'b1001000101: data <= 20'b11010000001101001011;
        10'b1001000110: data <= 20'b11001000010100100011;
        10'b1001000111: data <= 20'b11000111100100100000;
        10'b1001001000: data <= 20'b01001110110101010011;
        10'b1001001001: data <= 20'b01001000011011011001;
        10'b1001001010: data <= 20'b01000010100011101000;
        10'b1001001011: data <= 20'b11000000000100001011;
        10'b1001001100: data <= 20'b01001110000100101000;
        10'b1001001101: data <= 20'b01001101001011101010;
        10'b1001001110: data <= 20'b11010100001100110001;
        10'b1001001111: data <= 20'b11010000101101000000;
        10'b1001010000: data <= 20'b01001000111011110010;
        10'b1001010001: data <= 20'b01000001000011110011;
        10'b1001010010: data <= 20'b11000001010100001001;
        10'b1001010011: data <= 20'b01001100010100111110;
        10'b1001010100: data <= 20'b01001001110011111101;
        10'b1001010101: data <= 20'b01001001101011110011;
        10'b1001010110: data <= 20'b01000100111100100001;
        10'b1001010111: data <= 20'b01000100111100001101;
        10'b1001011000: data <= 20'b00111010110011110011;
        10'b1001011001: data <= 20'b11000100000011111100;
        10'b1001011010: data <= 20'b11010000110101000000;
        10'b1001011011: data <= 20'b01001010000100000011;
        10'b1001011100: data <= 20'b01000110110011110111;
        10'b1001011101: data <= 20'b01000100010011101111;
        10'b1001011110: data <= 20'b01000000100100001000;
        10'b1001011111: data <= 20'b11000100100100011010;
        10'b1001100000: data <= 20'b11000111101100000100;
        10'b1001100001: data <= 20'b11001011011100101101;
        10'b1001100010: data <= 20'b01001011101011010111;
        10'b1001100011: data <= 20'b01000101100011111010;
        10'b1001100100: data <= 20'b00111110100100000110;
        10'b1001100101: data <= 20'b01000000000100011101;
        10'b1001100110: data <= 20'b01000011110100100110;
        10'b1001100111: data <= 20'b01001100001101001101;
        10'b1001101000: data <= 20'b00111111101100100101;
        10'b1001101001: data <= 20'b01001000001100011110;
        10'b1001101010: data <= 20'b01000100110011100011;
        10'b1001101011: data <= 20'b10110111100011111011;
        10'b1001101100: data <= 20'b11000011000100101000;
        10'b1001101101: data <= 20'b01000110010100100101;
        10'b1001101110: data <= 20'b01001011010100100010;
        10'b1001101111: data <= 20'b01000111101100010010;
        10'b1001110000: data <= 20'b01000010111100000011;
        10'b1001110001: data <= 20'b00111101101011101100;
        10'b1001110010: data <= 20'b11000001001011111001;
        10'b1001110011: data <= 20'b11001100101100000101;
        10'b1001110100: data <= 20'b01001001100100101101;
        10'b1001110101: data <= 20'b01001000100100011111;
        10'b1001110110: data <= 20'b01001000000011101110;
        10'b1001110111: data <= 20'b01000010010011101001;
        10'b1001111000: data <= 20'b10111100010100001000;
        10'b1001111001: data <= 20'b11001001001100101001;
        10'b1001111010: data <= 20'b00111110001100101010;
        10'b1001111011: data <= 20'b01001110011100100101;
        10'b1001111100: data <= 20'b01001000100100011000;
        10'b1001111101: data <= 20'b01000101110100001111;
        10'b1001111110: data <= 20'b01000001000100001000;
        10'b1001111111: data <= 20'b10111000010100010100;
        10'b1010000000: data <= 20'b11001101000101000011;
        10'b1010000001: data <= 20'b01001000101100011101;
        10'b1010000010: data <= 20'b01000110101100010011;
        10'b1010000011: data <= 20'b01001000011011101110;
        10'b1010000100: data <= 20'b01000000010100000010;
        10'b1010000101: data <= 20'b10111100100100010110;
        10'b1010000110: data <= 20'b10111101010100011100;
        10'b1010000111: data <= 20'b11000100000100110010;
        10'b1010001000: data <= 20'b01001010101100000111;
        10'b1010001001: data <= 20'b01000101011011110100;
        10'b1010001010: data <= 20'b01000000001011010001;
        10'b1010001011: data <= 20'b11000111101100011011;
        10'b1010001100: data <= 20'b11001100001100111000;
        10'b1010001101: data <= 20'b11000111110100101101;
        10'b1010001110: data <= 20'b11000101110100110001;
        10'b1010001111: data <= 20'b01001100010011110101;
        10'b1010010000: data <= 20'b01000101000011010000;
        10'b1010010001: data <= 20'b00111011000011111001;
        10'b1010010010: data <= 20'b11001011000100100111;
        10'b1010010011: data <= 20'b01001100001100010110;
        10'b1010010100: data <= 20'b01001100111100100001;
        10'b1010010101: data <= 20'b11010000100101010001;
        10'b1010010110: data <= 20'b01001111110011011110;
        10'b1010010111: data <= 20'b01000100110011101110;
        10'b1010011000: data <= 20'b00110001010100000010;
        10'b1010011001: data <= 20'b11001000100100100000;
        10'b1010011010: data <= 20'b01001100100011100100;
        10'b1010011011: data <= 20'b01001000101011101011;
        10'b1010011100: data <= 20'b01001000101100001001;
        10'b1010011101: data <= 20'b01000100011100011111;
        10'b1010011110: data <= 20'b01000001000011111010;
        10'b1010011111: data <= 20'b10111110110100000011;
        10'b1010100000: data <= 20'b11001000100100010001;
        10'b1010100001: data <= 20'b01001110110100001000;
        10'b1010100010: data <= 20'b01000111110011100011;
        10'b1010100011: data <= 20'b01000100010011101101;
        10'b1010100100: data <= 20'b00111111100100001111;
        10'b1010100101: data <= 20'b01000011100100100010;
        10'b1010100110: data <= 20'b11001010010100010100;
        10'b1010100111: data <= 20'b11001001101100000111;
        10'b1010101000: data <= 20'b01001101101101000010;
        10'b1010101001: data <= 20'b01001000000011011110;
        10'b1010101010: data <= 20'b01000001110011110111;
        10'b1010101011: data <= 20'b10111110110100010110;
        10'b1010101100: data <= 20'b01000110110100100101;
        10'b1010101101: data <= 20'b01001011010100101001;
        10'b1010101110: data <= 20'b01000010011100110011;
        10'b1010101111: data <= 20'b01000001011100100101;
        10'b1010110000: data <= 20'b01000111011100000000;
        10'b1010110001: data <= 20'b00111111000011101111;
        10'b1010110010: data <= 20'b11000100110100001001;
        10'b1010110011: data <= 20'b01001000000100110001;
        10'b1010110100: data <= 20'b01001001000100011100;
        10'b1010110101: data <= 20'b01001010010011001111;
        10'b1010110110: data <= 20'b01000100101100001000;
        10'b1010110111: data <= 20'b01000000011011110000;
        10'b1010111000: data <= 20'b10111100011011011011;
        10'b1010111001: data <= 20'b11000110001100000010;
        10'b1010111010: data <= 20'b11010011000101100100;
        10'b1010111011: data <= 20'b01001001010100011001;
        10'b1010111100: data <= 20'b01000111100100001101;
        10'b1010111101: data <= 20'b01000100110011110011;
        10'b1010111110: data <= 20'b00111110000100000101;
        10'b1010111111: data <= 20'b11000111100100011010;
        10'b1011000000: data <= 20'b11000001111100101000;
        10'b1011000001: data <= 20'b01000010011100101110;
        10'b1011000010: data <= 20'b01001011010011101101;
        10'b1011000011: data <= 20'b01000101110100001001;
        10'b1011000100: data <= 20'b01000000110100001101;
        10'b1011000101: data <= 20'b00111100110100010101;
        10'b1011000110: data <= 20'b10111101000100100100;
        10'b1011000111: data <= 20'b01001101111100110001;
        10'b1011001000: data <= 20'b01000110001100010111;
        10'b1011001001: data <= 20'b01000110001100010000;
        10'b1011001010: data <= 20'b01000100010011100010;
        10'b1011001011: data <= 20'b11000000110011111001;
        10'b1011001100: data <= 20'b11000000000100100011;
        10'b1011001101: data <= 20'b00110010100100100110;
        10'b1011001110: data <= 20'b01001101010100101110;
        10'b1011001111: data <= 20'b01000111011100000000;
        10'b1011010000: data <= 20'b01000010011011100100;
        10'b1011010001: data <= 20'b10111110111010011111;
        10'b1011010010: data <= 20'b11000011001100100100;
        10'b1011010011: data <= 20'b11010001001101000000;
        10'b1011010100: data <= 20'b00111100110100110010;
        10'b1011010101: data <= 20'b01001001010100110001;
        10'b1011010110: data <= 20'b01001000000011010010;
        10'b1011010111: data <= 20'b01000001010011110010;
        10'b1011011000: data <= 20'b11000000110100001100;
        10'b1011011001: data <= 20'b01001111101101000010;
        10'b1011011010: data <= 20'b01001001011100011110;
        10'b1011011011: data <= 20'b01001101101100100000;
        10'b1011011100: data <= 20'b01001011010100110011;
        10'b1011011101: data <= 20'b01001000010100000011;
        10'b1011011110: data <= 20'b00111111110100000010;
        10'b1011011111: data <= 20'b11000000110100010001;
        10'b1011100000: data <= 20'b01000111110101010001;
        10'b1011100001: data <= 20'b01001001011100000001;
        10'b1011100010: data <= 20'b01000110111011111011;
        10'b1011100011: data <= 20'b01000111011100000111;
        10'b1011100100: data <= 20'b01000100100100001100;
        10'b1011100101: data <= 20'b10111100100100010000;
        10'b1011100110: data <= 20'b11000100000100010001;
        10'b1011100111: data <= 20'b11001110000100110110;
        10'b1011101000: data <= 20'b01001010001011100011;
        10'b1011101001: data <= 20'b01000101010011001110;
        10'b1011101010: data <= 20'b00111101110011111000;
        10'b1011101011: data <= 20'b01000101010100101100;
        10'b1011101100: data <= 20'b01001100100100111000;
        10'b1011101101: data <= 20'b11001011100100001110;
        10'b1011101110: data <= 20'b11001101111100001110;
        10'b1011101111: data <= 20'b01001011101100000111;
        10'b1011110000: data <= 20'b01000100100011101001;
        10'b1011110001: data <= 20'b00110000100100000001;
        10'b1011110010: data <= 20'b10111110010100110001;
        10'b1011110011: data <= 20'b01001010100100011001;
        10'b1011110100: data <= 20'b01001101011011011110;
        10'b1011110101: data <= 20'b00110100101100101110;
        10'b1011110110: data <= 20'b01000111001100100010;
        10'b1011110111: data <= 20'b01000011110011011000;
        10'b1011111000: data <= 20'b10111100000011111000;
        10'b1011111001: data <= 20'b11001010100100100110;
        10'b1011111010: data <= 20'b01001010110100011011;
        10'b1011111011: data <= 20'b01001000110100000110;
        10'b1011111100: data <= 20'b01001000001100000000;
        10'b1011111101: data <= 20'b01000001111011110100;
        10'b1011111110: data <= 20'b00101110110011101110;
        10'b1011111111: data <= 20'b11000011001011011110;
        10'b1100000000: data <= 20'b11001010101100010000;
        10'b1100000001: data <= 20'b01001101100100010101;
        10'b1100000010: data <= 20'b01000111110100000110;
        10'b1100000011: data <= 20'b01000100110100000010;
        10'b1100000100: data <= 20'b01000001100100001000;
        10'b1100000101: data <= 20'b00110111010100011001;
        10'b1100000110: data <= 20'b11001101101100011001;
        10'b1100000111: data <= 20'b11000000011100100111;
        10'b1100001000: data <= 20'b01001001111100101100;
        10'b1100001001: data <= 20'b01001000000011110111;
        10'b1100001010: data <= 20'b01000001000100000010;
        10'b1100001011: data <= 20'b00101011100100011000;
        10'b1100001100: data <= 20'b01000000000100100001;
        10'b1100001101: data <= 20'b01001000000100110101;
        10'b1100001110: data <= 20'b01001000101100100001;
        10'b1100001111: data <= 20'b01000100101100010011;
        10'b1100010000: data <= 20'b01000101011100000000;
        10'b1100010001: data <= 20'b00111001000011010001;
        10'b1100010010: data <= 20'b11001000000100001101;
        10'b1100010011: data <= 20'b01000000100100101011;
        10'b1100010100: data <= 20'b01000110100100101001;
        10'b1100010101: data <= 20'b01001010101011011001;
        10'b1100010110: data <= 20'b01000100101011110001;
        10'b1100010111: data <= 20'b00111100100011010110;
        10'b1100011000: data <= 20'b11000101101100001111;
        10'b1100011001: data <= 20'b11000100001100100111;
        10'b1100011010: data <= 20'b01010101000101010010;
        10'b1100011011: data <= 20'b01001000010100101000;
        10'b1100011100: data <= 20'b01001001010100010110;
        10'b1100011101: data <= 20'b01000100100011110001;
        10'b1100011110: data <= 20'b00111001100100000100;
        10'b1100011111: data <= 20'b11001010000100100001;
        10'b1100100000: data <= 20'b01001001001100100111;
        10'b1100100001: data <= 20'b01001000101100100000;
        10'b1100100010: data <= 20'b01001100010011111110;
        10'b1100100011: data <= 20'b01000111100100011001;
        10'b1100100100: data <= 20'b01000010100100001000;
        10'b1100100101: data <= 20'b00011111000100010000;
        10'b1100100110: data <= 20'b11000110000100100011;
        10'b1100100111: data <= 20'b01001101001100010100;
        10'b1100101000: data <= 20'b01000111001100000011;
        10'b1100101001: data <= 20'b01000101001011111101;
        10'b1100101010: data <= 20'b01000001101011000011;
        10'b1100101011: data <= 20'b11000111110100010000;
        10'b1100101100: data <= 20'b11000010100100011001;
        10'b1100101101: data <= 20'b11000110110100100010;
        10'b1100101110: data <= 20'b01010000000100011001;
        10'b1100101111: data <= 20'b01000111001011100001;
        10'b1100110000: data <= 20'b01000001110011100000;
        10'b1100110001: data <= 20'b11000100000100010010;
        10'b1100110010: data <= 20'b01001110111011101011;
        10'b1100110011: data <= 20'b01010111110101000011;
        10'b1100110100: data <= 20'b11001100100100100100;
        10'b1100110101: data <= 20'b01011010101011101111;
        10'b1100110110: data <= 20'b01000111101010011000;
        10'b1100110111: data <= 20'b01000000010011110101;
        10'b1100111000: data <= 20'b11000011110100010010;
        10'b1100111001: data <= 20'b01001101100100100101;
        10'b1100111010: data <= 20'b01001010010011010101;
        10'b1100111011: data <= 20'b01001100011100100011;
        10'b1100111100: data <= 20'b00111010011100110001;
        10'b1100111101: data <= 20'b01000111001011111010;
        10'b1100111110: data <= 20'b00111100000011110111;
        10'b1100111111: data <= 20'b11000100100100000111;
        10'b1101000000: data <= 20'b01001111010101000001;
        10'b1101000001: data <= 20'b01001001010011111100;
        10'b1101000010: data <= 20'b01000111010011100100;
        10'b1101000011: data <= 20'b01000100101011110011;
        10'b1101000100: data <= 20'b00111111100011111011;
        10'b1101000101: data <= 20'b11000010010011111111;
        10'b1101000110: data <= 20'b11000110111011010000;
        10'b1101000111: data <= 20'b11010010101101000010;
        10'b1101001000: data <= 20'b01001001100011110111;
        10'b1101001001: data <= 20'b01000101010011111010;
        10'b1101001010: data <= 20'b01000000000100001000;
        10'b1101001011: data <= 20'b01000001010100011010;
        10'b1101001100: data <= 20'b00111100010100101110;
        10'b1101001101: data <= 20'b11001000111100101101;
        10'b1101001110: data <= 20'b10111101111100101100;
        10'b1101001111: data <= 20'b01001010001100001100;
        10'b1101010000: data <= 20'b01000100010011110100;
        10'b1101010001: data <= 20'b10111001100100000110;
        10'b1101010010: data <= 20'b00111101110100100110;
        10'b1101010011: data <= 20'b01000110100100100101;
        10'b1101010100: data <= 20'b01001110000011101111;
        10'b1101010101: data <= 20'b01000101011100011001;
        10'b1101010110: data <= 20'b01000100001100010000;
        10'b1101010111: data <= 20'b01000001001011010001;
        10'b1101011000: data <= 20'b11000001100010101011;
        10'b1101011001: data <= 20'b11001011100100110001;
        10'b1101011010: data <= 20'b01001000010100100110;
        10'b1101011011: data <= 20'b01001001010100011100;
        10'b1101011100: data <= 20'b01000111011011110010;
        10'b1101011101: data <= 20'b01000001010011000000;
        10'b1101011110: data <= 20'b11000000100011111000;
        10'b1101011111: data <= 20'b11000100111100011100;
        10'b1101100000: data <= 20'b11000110001100110001;
        10'b1101100001: data <= 20'b01001101000100100100;
        10'b1101100010: data <= 20'b01001000000100011000;
        10'b1101100011: data <= 20'b01000110010100000101;
        10'b1101100100: data <= 20'b01000000110100000100;
        10'b1101100101: data <= 20'b10111110010100010101;
        10'b1101100110: data <= 20'b11001000011101001110;
        10'b1101100111: data <= 20'b01000110101100100001;
        10'b1101101000: data <= 20'b01001000111100011101;
        10'b1101101001: data <= 20'b01001000010100001000;
        10'b1101101010: data <= 20'b01000001010100001011;
        10'b1101101011: data <= 20'b00111001110100010011;
        10'b1101101100: data <= 20'b10111100100100011100;
        10'b1101101101: data <= 20'b01000010110101000001;
        10'b1101101110: data <= 20'b01001000111100010000;
        10'b1101101111: data <= 20'b01000101001100000001;
        10'b1101110000: data <= 20'b01000010001011110101;
        10'b1101110001: data <= 20'b11000000101100000110;
        10'b1101110010: data <= 20'b11001010010100011101;
        10'b1101110011: data <= 20'b11000010010100100100;
        10'b1101110100: data <= 20'b11000000010100110101;
        10'b1101110101: data <= 20'b01001010001011101101;
        10'b1101110110: data <= 20'b01000100011010011010;
        10'b1101110111: data <= 20'b00110100100011110111;
        10'b1101111000: data <= 20'b11010010111100101011;
        10'b1101111001: data <= 20'b01001011101100101001;
        10'b1101111010: data <= 20'b01010101010101011101;
        10'b1101111011: data <= 20'b11001000010100111011;
        10'b1101111100: data <= 20'b01001100000011110100;
        10'b1101111101: data <= 20'b01000100000011110000;
        10'b1101111110: data <= 20'b10110100010100000011;
        10'b1101111111: data <= 20'b11001011100100110001;
        10'b1110000000: data <= 20'b01001011011011111110;
        10'b1110000001: data <= 20'b01001001011100000101;
        10'b1110000010: data <= 20'b01001100101100101010;
        10'b1110000011: data <= 20'b01001100001100100111;
        10'b1110000100: data <= 20'b01000001110011111010;
        10'b1110000101: data <= 20'b10111101110100000101;
        10'b1110000110: data <= 20'b11001010000100100001;
        10'b1110000111: data <= 20'b01001100010011101011;
        10'b1110001000: data <= 20'b01000111010011000010;
        10'b1110001001: data <= 20'b01000100110010111001;
        10'b1110001010: data <= 20'b01000001010100000100;
        10'b1110001011: data <= 20'b10111010010100100000;
        10'b1110001100: data <= 20'b11000101110100000100;
        10'b1110001101: data <= 20'b11001010100011101001;
        10'b1110001110: data <= 20'b01001110101100001111;
        10'b1110001111: data <= 20'b01000110110011101000;
        10'b1110010000: data <= 20'b01000001010011111001;
        10'b1110010001: data <= 20'b10110011010100011110;
        10'b1110010010: data <= 20'b01000111010100100100;
        10'b1110010011: data <= 20'b01001111110101001101;
        10'b1110010100: data <= 20'b11000111111100101010;
        10'b1110010101: data <= 20'b01000111001100110001;
        10'b1110010110: data <= 20'b01000110111010101110;
        10'b1110010111: data <= 20'b00111101110011110110;
        10'b1110011000: data <= 20'b11000101000100011001;
        10'b1110011001: data <= 20'b01001000100100100111;
        10'b1110011010: data <= 20'b01001001110100011011;
        10'b1110011011: data <= 20'b01001010001100011100;
        10'b1110011100: data <= 20'b01000011011100010011;
        10'b1110011101: data <= 20'b01000011011011111101;
        10'b1110011110: data <= 20'b10110100000011001110;
        10'b1110011111: data <= 20'b11000111110011011000;
        10'b1110100000: data <= 20'b01001100100100110111;
        10'b1110100001: data <= 20'b01001000110100010110;
        10'b1110100010: data <= 20'b01001000010100000010;
        10'b1110100011: data <= 20'b01000100010010011000;
        10'b1110100100: data <= 20'b00111011010100000000;
        10'b1110100101: data <= 20'b11000111101011100101;
        10'b1110100110: data <= 20'b11000101011100100000;
        10'b1110100111: data <= 20'b01001001111101000000;
        10'b1110101000: data <= 20'b01001001100100010000;
        10'b1110101001: data <= 20'b01000101100100001010;
        10'b1110101010: data <= 20'b01000010000100001001;
        10'b1110101011: data <= 20'b00111100100100010011;
        10'b1110101100: data <= 20'b11000100110100101100;
        10'b1110101101: data <= 20'b01000111011100101110;
        10'b1110101110: data <= 20'b01000101011100011111;
        10'b1110101111: data <= 20'b01001000111100001001;
        10'b1110110000: data <= 20'b01000011110011111101;
        10'b1110110001: data <= 20'b10111101000100001111;
        10'b1110110010: data <= 20'b00110011000100011111;
        10'b1110110011: data <= 20'b00110111000100101000;
        10'b1110110100: data <= 20'b01001101101011111100;
        10'b1110110101: data <= 20'b01000110001100000111;
        10'b1110110110: data <= 20'b01000010101011111001;
        10'b1110110111: data <= 20'b00101001111011110110;
        10'b1110111000: data <= 20'b11000101111100010011;
        10'b1110111001: data <= 20'b11001001100100110011;
        10'b1110111010: data <= 20'b00111110010100101100;
        10'b1110111011: data <= 20'b01001100000100101000;
        10'b1110111100: data <= 20'b01000110111011011011;
        10'b1110111101: data <= 20'b01000000100011101011;
        10'b1110111110: data <= 20'b11000100110100001010;
        10'b1110111111: data <= 20'b01001000001100110010;
        10'b1111000000: data <= 20'b01001010001100101110;
        10'b1111000001: data <= 20'b01001101110100111010;
        10'b1111000010: data <= 20'b01001001110100101111;
        10'b1111000011: data <= 20'b01000111000011110111;
        10'b1111000100: data <= 20'b00111110110100000001;
        10'b1111000101: data <= 20'b11000011000100010100;
        10'b1111000110: data <= 20'b01010001001100011001;
        10'b1111000111: data <= 20'b01001000111100001011;
        10'b1111001000: data <= 20'b01001000011100001101;
        10'b1111001001: data <= 20'b01001100110100000011;
        10'b1111001010: data <= 20'b01000101010100001001;
        10'b1111001011: data <= 20'b00101100110100001010;
        10'b1111001100: data <= 20'b11000100000100010100;
        10'b1111001101: data <= 20'b01001110010101010001;
        10'b1111001110: data <= 20'b01001000111011101110;
        10'b1111001111: data <= 20'b01000101001011001101;
        10'b1111010000: data <= 20'b00111110000011110001;
        10'b1111010001: data <= 20'b01001000110100110000;
        10'b1111010010: data <= 20'b11001001010100101000;
        10'b1111010011: data <= 20'b11001000010100010010;
        10'b1111010100: data <= 20'b11010001100100101000;
        10'b1111010101: data <= 20'b01001001101011100010;
        10'b1111010110: data <= 20'b01000100000011101001;
        10'b1111010111: data <= 20'b10110110100100000101;
        10'b1111011000: data <= 20'b01001000000100110001;
        10'b1111011001: data <= 20'b01001100000100011000;
        10'b1111011010: data <= 20'b01000101001101010011;
        10'b1111011011: data <= 20'b11001000111100110001;
        10'b1111011100: data <= 20'b01001001111100010011;
        10'b1111011101: data <= 20'b01000010110011101100;
        10'b1111011110: data <= 20'b10111110000100000010;
        10'b1111011111: data <= 20'b11000100110100111000;
        10'b1111100000: data <= 20'b01001010000100010100;
        10'b1111100001: data <= 20'b01001001110011110110;
        10'b1111100010: data <= 20'b01000110011100011001;
        10'b1111100011: data <= 20'b01000010011100001011;
        10'b1111100100: data <= 20'b00111101010011011011;
        10'b1111100101: data <= 20'b11000010010011100100;
        10'b1111100110: data <= 20'b11001101110100010000;
        10'b1111100111: data <= 20'b01001011010100010100;
        10'b1111101000: data <= 20'b01000111100100000100;
        10'b1111101001: data <= 20'b01000101100011110100;
        10'b1111101010: data <= 20'b01000001000100000001;
        10'b1111101011: data <= 20'b10111111100100010111;
        10'b1111101100: data <= 20'b11001000001100010011;
        10'b1111101101: data <= 20'b11000111101100101000;
        10'b1111101110: data <= 20'b01001101001100010001;
        10'b1111101111: data <= 20'b01000110110100000001;
        10'b1111110000: data <= 20'b01000001010100000101;
        10'b1111110001: data <= 20'b00111110010100010111;
        10'b1111110010: data <= 20'b00111111000100100001;
        10'b1111110011: data <= 20'b01010100000101010011;
        10'b1111110100: data <= 20'b01000100101100100011;
        10'b1111110101: data <= 20'b01000110001100011101;
        10'b1111110110: data <= 20'b01000110001010101011;
        10'b1111110111: data <= 20'b00111000000011110101;
        10'b1111111000: data <= 20'b11000100100100100000;
        10'b1111111001: data <= 20'b01000010010100100110;
        10'b1111111010: data <= 20'b01001001000100101100;
        10'b1111111011: data <= 20'b01001001001100001111;
        10'b1111111100: data <= 20'b00111110001100000011;
    
    endcase
    end
    end

    assign Q = data;

    endmodule

        
