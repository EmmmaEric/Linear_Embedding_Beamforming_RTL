
module memory_rom_37(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbe3f3410;
    11'b00000000001: data <= 32'hbb00325c;
    11'b00000000010: data <= 32'h3b63af4d;
    11'b00000000011: data <= 32'h3f23388d;
    11'b00000000100: data <= 32'h36d93eb0;
    11'b00000000101: data <= 32'hbdf83f47;
    11'b00000000110: data <= 32'hbe0d3c3d;
    11'b00000000111: data <= 32'h32b9380e;
    11'b00000001000: data <= 32'h3d4b3488;
    11'b00000001001: data <= 32'h3a89b775;
    11'b00000001010: data <= 32'h3354be18;
    11'b00000001011: data <= 32'h3b4ebd81;
    11'b00000001100: data <= 32'h3f9034d9;
    11'b00000001101: data <= 32'h3e1e3e1f;
    11'b00000001110: data <= 32'h2d7e38c8;
    11'b00000001111: data <= 32'hbb3cbd62;
    11'b00000010000: data <= 32'hbc11bf70;
    11'b00000010001: data <= 32'hbc52b9c1;
    11'b00000010010: data <= 32'hbce6a507;
    11'b00000010011: data <= 32'hb8b3ba63;
    11'b00000010100: data <= 32'h39bcbdec;
    11'b00000010101: data <= 32'h3c30b72c;
    11'b00000010110: data <= 32'hb5fb3db5;
    11'b00000010111: data <= 32'hbf844048;
    11'b00000011000: data <= 32'hbe243da1;
    11'b00000011001: data <= 32'h1f7638ac;
    11'b00000011010: data <= 32'h382834cb;
    11'b00000011011: data <= 32'hb5cdad9d;
    11'b00000011100: data <= 32'hb8f4b95a;
    11'b00000011101: data <= 32'h3b46b6d1;
    11'b00000011110: data <= 32'h41283abe;
    11'b00000011111: data <= 32'h409e3e4d;
    11'b00000100000: data <= 32'h384338c5;
    11'b00000100001: data <= 32'hb963bb37;
    11'b00000100010: data <= 32'hb8a9bc1d;
    11'b00000100011: data <= 32'hb426b011;
    11'b00000100100: data <= 32'hb51bb402;
    11'b00000100101: data <= 32'hade5bf31;
    11'b00000100110: data <= 32'h3919c13e;
    11'b00000100111: data <= 32'h3a0dbca9;
    11'b00000101000: data <= 32'hb5bf3c85;
    11'b00000101001: data <= 32'hbde03f51;
    11'b00000101010: data <= 32'hbce63a5a;
    11'b00000101011: data <= 32'hb620af7b;
    11'b00000101100: data <= 32'hb9169d2f;
    11'b00000101101: data <= 32'hbecd3309;
    11'b00000101110: data <= 32'hbddcab4a;
    11'b00000101111: data <= 32'h3987a90d;
    11'b00000110000: data <= 32'h411f3a74;
    11'b00000110001: data <= 32'h40233df1;
    11'b00000110010: data <= 32'h30d23c1e;
    11'b00000110011: data <= 32'hb9df32eb;
    11'b00000110100: data <= 32'ha8ff34a1;
    11'b00000110101: data <= 32'h39143973;
    11'b00000110110: data <= 32'h35f1b300;
    11'b00000110111: data <= 32'h2efac056;
    11'b00000111000: data <= 32'h3904c1b5;
    11'b00000111001: data <= 32'h3c58bca1;
    11'b00000111010: data <= 32'h38603bd0;
    11'b00000111011: data <= 32'hb5dc3c99;
    11'b00000111100: data <= 32'hb8dab40e;
    11'b00000111101: data <= 32'hb8cbbbc1;
    11'b00000111110: data <= 32'hbd90b47b;
    11'b00000111111: data <= 32'hc0c73532;
    11'b00001000000: data <= 32'hbf3eb027;
    11'b00001000001: data <= 32'h3685b8d9;
    11'b00001000010: data <= 32'h3fa827b0;
    11'b00001000011: data <= 32'h3c473c8d;
    11'b00001000100: data <= 32'hb9823dfd;
    11'b00001000101: data <= 32'hbb8b3d14;
    11'b00001000110: data <= 32'h34a53d3d;
    11'b00001000111: data <= 32'h3b7d3d0d;
    11'b00001001000: data <= 32'h32ec2cdb;
    11'b00001001001: data <= 32'hb53cbee4;
    11'b00001001010: data <= 32'h3823c03a;
    11'b00001001011: data <= 32'h3eecb81a;
    11'b00001001100: data <= 32'h3f0d3c14;
    11'b00001001101: data <= 32'h3a6b3877;
    11'b00001001110: data <= 32'h2805bb99;
    11'b00001001111: data <= 32'hb6f9bce9;
    11'b00001010000: data <= 32'hbd17b014;
    11'b00001010001: data <= 32'hc01c351d;
    11'b00001010010: data <= 32'hbdf7ba52;
    11'b00001010011: data <= 32'h3381bf42;
    11'b00001010100: data <= 32'h3c70bc6e;
    11'b00001010101: data <= 32'h2ccf38ef;
    11'b00001010110: data <= 32'hbd123e65;
    11'b00001010111: data <= 32'hbbc53e39;
    11'b00001011000: data <= 32'h35333db0;
    11'b00001011001: data <= 32'h37553d32;
    11'b00001011010: data <= 32'hba603723;
    11'b00001011011: data <= 32'hbd2cba86;
    11'b00001011100: data <= 32'h32dcbc00;
    11'b00001011101: data <= 32'h405332bd;
    11'b00001011110: data <= 32'h40ef3c5e;
    11'b00001011111: data <= 32'h3d4335a2;
    11'b00001100000: data <= 32'h356aba89;
    11'b00001100001: data <= 32'h26c9b890;
    11'b00001100010: data <= 32'hb6833894;
    11'b00001100011: data <= 32'hbc10365e;
    11'b00001100100: data <= 32'hbaa1be07;
    11'b00001100101: data <= 32'h326dc1bd;
    11'b00001100110: data <= 32'h392cbfad;
    11'b00001100111: data <= 32'hb29231fb;
    11'b00001101000: data <= 32'hbc2b3cdc;
    11'b00001101001: data <= 32'hb8903b31;
    11'b00001101010: data <= 32'h33c638fd;
    11'b00001101011: data <= 32'hb6603ad6;
    11'b00001101100: data <= 32'hc015399b;
    11'b00001101101: data <= 32'hc084abd0;
    11'b00001101110: data <= 32'hb207b560;
    11'b00001101111: data <= 32'h400e35f2;
    11'b00001110000: data <= 32'h405d3b83;
    11'b00001110001: data <= 32'h3afd37cf;
    11'b00001110010: data <= 32'h31a99fbd;
    11'b00001110011: data <= 32'h382e3928;
    11'b00001110100: data <= 32'h38d63e12;
    11'b00001110101: data <= 32'hac6c3945;
    11'b00001110110: data <= 32'hb6babee4;
    11'b00001110111: data <= 32'h3108c21c;
    11'b00001111000: data <= 32'h399abf91;
    11'b00001111001: data <= 32'h362f2d8c;
    11'b00001111010: data <= 32'hab0a3887;
    11'b00001111011: data <= 32'h3232b3eb;
    11'b00001111100: data <= 32'h34a8b761;
    11'b00001111101: data <= 32'hbbb635e9;
    11'b00001111110: data <= 32'hc15e3a79;
    11'b00001111111: data <= 32'hc1402f78;
    11'b00010000000: data <= 32'hb78eb8b2;
    11'b00010000001: data <= 32'h3d8ab459;
    11'b00010000010: data <= 32'h3c63372a;
    11'b00010000011: data <= 32'hb1773956;
    11'b00010000100: data <= 32'hb3813a9d;
    11'b00010000101: data <= 32'h3aaa3e7b;
    11'b00010000110: data <= 32'h3c844054;
    11'b00010000111: data <= 32'h2da93c0a;
    11'b00010001000: data <= 32'hb99fbcfe;
    11'b00010001001: data <= 32'had1ac07b;
    11'b00010001010: data <= 32'h3c2cbc4b;
    11'b00010001011: data <= 32'h3d6f350b;
    11'b00010001100: data <= 32'h3c441dbb;
    11'b00010001101: data <= 32'h3b7cbc92;
    11'b00010001110: data <= 32'h388dbc1b;
    11'b00010001111: data <= 32'hba49358c;
    11'b00010010000: data <= 32'hc0923b41;
    11'b00010010001: data <= 32'hc058b3cd;
    11'b00010010010: data <= 32'hb7cbbe21;
    11'b00010010011: data <= 32'h38edbd6c;
    11'b00010010100: data <= 32'hacefb29e;
    11'b00010010101: data <= 32'hbc3338ce;
    11'b00010010110: data <= 32'hb7503c14;
    11'b00010010111: data <= 32'h3b8c3ebb;
    11'b00010011000: data <= 32'h3b894039;
    11'b00010011001: data <= 32'hb92d3d0c;
    11'b00010011010: data <= 32'hbe68b5f2;
    11'b00010011011: data <= 32'hb845bbb7;
    11'b00010011100: data <= 32'h3d0eabb3;
    11'b00010011101: data <= 32'h3fc038c6;
    11'b00010011110: data <= 32'h3e2db3f9;
    11'b00010011111: data <= 32'h3cd4bd27;
    11'b00010100000: data <= 32'h3bb1b947;
    11'b00010100001: data <= 32'h2c0b3bb2;
    11'b00010100010: data <= 32'hbc6c3c90;
    11'b00010100011: data <= 32'hbcf2b9be;
    11'b00010100100: data <= 32'hb4dec0dd;
    11'b00010100101: data <= 32'h3016c048;
    11'b00010100110: data <= 32'hb8fcb939;
    11'b00010100111: data <= 32'hbc823361;
    11'b00010101000: data <= 32'hb13b35c1;
    11'b00010101001: data <= 32'h3c0c3a1c;
    11'b00010101010: data <= 32'h35943db2;
    11'b00010101011: data <= 32'hbed93d36;
    11'b00010101100: data <= 32'hc1183637;
    11'b00010101101: data <= 32'hbbfeaa28;
    11'b00010101110: data <= 32'h3c5936ab;
    11'b00010101111: data <= 32'h3e8038a0;
    11'b00010110000: data <= 32'h3c02b3ff;
    11'b00010110001: data <= 32'h3ab9ba0b;
    11'b00010110010: data <= 32'h3d0d35b1;
    11'b00010110011: data <= 32'h3c463f91;
    11'b00010110100: data <= 32'h2d0f3e03;
    11'b00010110101: data <= 32'hb806bab7;
    11'b00010110110: data <= 32'hb1ddc123;
    11'b00010110111: data <= 32'h2c29c013;
    11'b00010111000: data <= 32'hb50eb8c3;
    11'b00010111001: data <= 32'hb5ccb415;
    11'b00010111010: data <= 32'h38a4ba38;
    11'b00010111011: data <= 32'h3cc3b855;
    11'b00010111100: data <= 32'had0938e6;
    11'b00010111101: data <= 32'hc0923ce2;
    11'b00010111110: data <= 32'hc1b93943;
    11'b00010111111: data <= 32'hbcb5a1d7;
    11'b00011000000: data <= 32'h38872560;
    11'b00011000001: data <= 32'h385a2fd5;
    11'b00011000010: data <= 32'hb3cdb30d;
    11'b00011000011: data <= 32'h2f27ae3b;
    11'b00011000100: data <= 32'h3d773cf8;
    11'b00011000101: data <= 32'h3ea54104;
    11'b00011000110: data <= 32'h38313f36;
    11'b00011000111: data <= 32'hb816b717;
    11'b00011001000: data <= 32'hb5c2befe;
    11'b00011001001: data <= 32'h340abc26;
    11'b00011001010: data <= 32'h372cac60;
    11'b00011001011: data <= 32'h3932b8d5;
    11'b00011001100: data <= 32'h3d42bee5;
    11'b00011001101: data <= 32'h3de2bd91;
    11'b00011001110: data <= 32'h2c7034a6;
    11'b00011001111: data <= 32'hbf7e3ce8;
    11'b00011010000: data <= 32'hc081372a;
    11'b00011010001: data <= 32'hbb62b9c9;
    11'b00011010010: data <= 32'h142cbb6e;
    11'b00011010011: data <= 32'hb95bb84d;
    11'b00011010100: data <= 32'hbd9eb56a;
    11'b00011010101: data <= 32'hb6e32cfe;
    11'b00011010110: data <= 32'h3d693d21;
    11'b00011010111: data <= 32'h3e7240ab;
    11'b00011011000: data <= 32'h293f3f4d;
    11'b00011011001: data <= 32'hbcfe33ec;
    11'b00011011010: data <= 32'hba91b707;
    11'b00011011011: data <= 32'h361b3406;
    11'b00011011100: data <= 32'h3bb83862;
    11'b00011011101: data <= 32'h3c62b9a9;
    11'b00011011110: data <= 32'h3dffbff8;
    11'b00011011111: data <= 32'h3ebebd2b;
    11'b00011100000: data <= 32'h3a1139b8;
    11'b00011100001: data <= 32'hb9503dd5;
    11'b00011100010: data <= 32'hbc362dd5;
    11'b00011100011: data <= 32'hb661be16;
    11'b00011100100: data <= 32'hb503beb0;
    11'b00011100101: data <= 32'hbd4ebb76;
    11'b00011100110: data <= 32'hbf0fb8b2;
    11'b00011100111: data <= 32'hb5c5b74c;
    11'b00011101000: data <= 32'h3d99356d;
    11'b00011101001: data <= 32'h3c9a3d9b;
    11'b00011101010: data <= 32'hbb1b3e1f;
    11'b00011101011: data <= 32'hc0463a8d;
    11'b00011101100: data <= 32'hbd0f389d;
    11'b00011101101: data <= 32'h34553c1b;
    11'b00011101110: data <= 32'h39e83a4c;
    11'b00011101111: data <= 32'h3844b94c;
    11'b00011110000: data <= 32'h3b5abe66;
    11'b00011110001: data <= 32'h3eaeb718;
    11'b00011110010: data <= 32'h3e473e48;
    11'b00011110011: data <= 32'h38e13f47;
    11'b00011110100: data <= 32'ha135a9ee;
    11'b00011110101: data <= 32'h23d7bed0;
    11'b00011110110: data <= 32'hb4d0be32;
    11'b00011110111: data <= 32'hbca6b994;
    11'b00011111000: data <= 32'hbcc7ba53;
    11'b00011111001: data <= 32'h3498bda1;
    11'b00011111010: data <= 32'h3e5dbc2f;
    11'b00011111011: data <= 32'h39ff346b;
    11'b00011111100: data <= 32'hbde23c81;
    11'b00011111101: data <= 32'hc0df3bdc;
    11'b00011111110: data <= 32'hbd373a0d;
    11'b00011111111: data <= 32'ha2293adc;
    11'b00100000000: data <= 32'hb18b3754;
    11'b00100000001: data <= 32'hba47b92e;
    11'b00100000010: data <= 32'hafa4bc02;
    11'b00100000011: data <= 32'h3dbb36ba;
    11'b00100000100: data <= 32'h400f4059;
    11'b00100000101: data <= 32'h3cc7400b;
    11'b00100000110: data <= 32'h33b03121;
    11'b00100000111: data <= 32'h1b9fbc1e;
    11'b00100001000: data <= 32'hafa3b7c6;
    11'b00100001001: data <= 32'hb7cc2ffe;
    11'b00100001010: data <= 32'hb3a4ba5c;
    11'b00100001011: data <= 32'h3c07c067;
    11'b00100001100: data <= 32'h3f40c010;
    11'b00100001101: data <= 32'h3a0fb550;
    11'b00100001110: data <= 32'hbcba3b65;
    11'b00100001111: data <= 32'hbf183a13;
    11'b00100010000: data <= 32'hba3a30ee;
    11'b00100010001: data <= 32'hb3b995d8;
    11'b00100010010: data <= 32'hbce9b1bb;
    11'b00100010011: data <= 32'hc027b9ec;
    11'b00100010100: data <= 32'hbbc6b9e2;
    11'b00100010101: data <= 32'h3caf387a;
    11'b00100010110: data <= 32'h3fc53fd8;
    11'b00100010111: data <= 32'h3aae3f38;
    11'b00100011000: data <= 32'hb5e73848;
    11'b00100011001: data <= 32'hb6a52f9a;
    11'b00100011010: data <= 32'h22083b77;
    11'b00100011011: data <= 32'h2cd23c46;
    11'b00100011100: data <= 32'h3480b8ea;
    11'b00100011101: data <= 32'h3caec0d1;
    11'b00100011110: data <= 32'h3f51c022;
    11'b00100011111: data <= 32'h3ca4acce;
    11'b00100100000: data <= 32'hb0233c56;
    11'b00100100001: data <= 32'hb7323694;
    11'b00100100010: data <= 32'h2d55b934;
    11'b00100100011: data <= 32'hb3d0ba54;
    11'b00100100100: data <= 32'hbf34b88b;
    11'b00100100101: data <= 32'hc12abab1;
    11'b00100100110: data <= 32'hbc6ebc16;
    11'b00100100111: data <= 32'h3c71b382;
    11'b00100101000: data <= 32'h3df43b53;
    11'b00100101001: data <= 32'hac5a3cb3;
    11'b00100101010: data <= 32'hbd1a3a38;
    11'b00100101011: data <= 32'hbae43c23;
    11'b00100101100: data <= 32'h20883f76;
    11'b00100101101: data <= 32'h2ad73e38;
    11'b00100101110: data <= 32'hb08cb6bd;
    11'b00100101111: data <= 32'h37f0c007;
    11'b00100110000: data <= 32'h3dfabd15;
    11'b00100110001: data <= 32'h3e8c3a21;
    11'b00100110010: data <= 32'h3c213dcb;
    11'b00100110011: data <= 32'h3a16327e;
    11'b00100110100: data <= 32'h3a45bbf2;
    11'b00100110101: data <= 32'ha94bba5b;
    11'b00100110110: data <= 32'hbe7fb42e;
    11'b00100110111: data <= 32'hc02fba01;
    11'b00100111000: data <= 32'hb816be95;
    11'b00100111001: data <= 32'h3d2ebdfe;
    11'b00100111010: data <= 32'h3c2eb61b;
    11'b00100111011: data <= 32'hba2f3735;
    11'b00100111100: data <= 32'hbebe39ac;
    11'b00100111101: data <= 32'hbad43cc0;
    11'b00100111110: data <= 32'ha58b3f35;
    11'b00100111111: data <= 32'hb8683d46;
    11'b00101000000: data <= 32'hbd57b61a;
    11'b00101000001: data <= 32'hb9b0bd93;
    11'b00101000010: data <= 32'h3b53b521;
    11'b00101000011: data <= 32'h3f513ddf;
    11'b00101000100: data <= 32'h3e4d3e81;
    11'b00101000101: data <= 32'h3c933258;
    11'b00101000110: data <= 32'h3b4fb8cf;
    11'b00101000111: data <= 32'h3239308f;
    11'b00101001000: data <= 32'hbb8039c2;
    11'b00101001001: data <= 32'hbc56b67e;
    11'b00101001010: data <= 32'h34a5c04b;
    11'b00101001011: data <= 32'h3e0cc0db;
    11'b00101001100: data <= 32'h3b0ebc96;
    11'b00101001101: data <= 32'hb9e32b1a;
    11'b00101001110: data <= 32'hbc9a364b;
    11'b00101001111: data <= 32'hb1ed38a2;
    11'b00101010000: data <= 32'h2de63b67;
    11'b00101010001: data <= 32'hbd3238fe;
    11'b00101010010: data <= 32'hc120b7b9;
    11'b00101010011: data <= 32'hbef6bbf6;
    11'b00101010100: data <= 32'h3696296b;
    11'b00101010101: data <= 32'h3e6d3d89;
    11'b00101010110: data <= 32'h3cd53d29;
    11'b00101010111: data <= 32'h386d33e7;
    11'b00101011000: data <= 32'h378e33a9;
    11'b00101011001: data <= 32'h35093df6;
    11'b00101011010: data <= 32'hb4713f6c;
    11'b00101011011: data <= 32'hb5ec2b88;
    11'b00101011100: data <= 32'h38b1c05b;
    11'b00101011101: data <= 32'h3dc1c0e7;
    11'b00101011110: data <= 32'h3be1bb8f;
    11'b00101011111: data <= 32'h22983239;
    11'b00101100000: data <= 32'h2e2729bd;
    11'b00101100001: data <= 32'h3b05b4b9;
    11'b00101100010: data <= 32'h367da6ab;
    11'b00101100011: data <= 32'hbea62e97;
    11'b00101100100: data <= 32'hc21ab82c;
    11'b00101100101: data <= 32'hbfe0bc0f;
    11'b00101100110: data <= 32'h347bb752;
    11'b00101100111: data <= 32'h3c8536ce;
    11'b00101101000: data <= 32'h340e3758;
    11'b00101101001: data <= 32'hb7b630d7;
    11'b00101101010: data <= 32'hae4c3b59;
    11'b00101101011: data <= 32'h357340cf;
    11'b00101101100: data <= 32'hac8a40f1;
    11'b00101101101: data <= 32'hb81a3602;
    11'b00101101110: data <= 32'h220ebeed;
    11'b00101101111: data <= 32'h3b55be77;
    11'b00101110000: data <= 32'h3c75a0d2;
    11'b00101110001: data <= 32'h3b553954;
    11'b00101110010: data <= 32'h3d27b185;
    11'b00101110011: data <= 32'h3ef9baa4;
    11'b00101110100: data <= 32'h3a48b4b0;
    11'b00101110101: data <= 32'hbd9a34b9;
    11'b00101110110: data <= 32'hc110b458;
    11'b00101110111: data <= 32'hbd41bd2f;
    11'b00101111000: data <= 32'h385fbdcc;
    11'b00101111001: data <= 32'h397dbace;
    11'b00101111010: data <= 32'hb8e6b75f;
    11'b00101111011: data <= 32'hbc8bb0a6;
    11'b00101111100: data <= 32'hb2fb3ba0;
    11'b00101111101: data <= 32'h371740a5;
    11'b00101111110: data <= 32'hb5974070;
    11'b00101111111: data <= 32'hbdb435e7;
    11'b00110000000: data <= 32'hbcaabc71;
    11'b00110000001: data <= 32'h2fd6b840;
    11'b00110000010: data <= 32'h3c233b56;
    11'b00110000011: data <= 32'h3d3d3bd9;
    11'b00110000100: data <= 32'h3ea9b475;
    11'b00110000101: data <= 32'h3fa0b9ec;
    11'b00110000110: data <= 32'h3c1435ce;
    11'b00110000111: data <= 32'hb9a23cf0;
    11'b00110001000: data <= 32'hbda634b7;
    11'b00110001001: data <= 32'hb4f7bdfa;
    11'b00110001010: data <= 32'h3b3ec067;
    11'b00110001011: data <= 32'h3737be7a;
    11'b00110001100: data <= 32'hbad0bb83;
    11'b00110001101: data <= 32'hbb0db81b;
    11'b00110001110: data <= 32'h36483515;
    11'b00110001111: data <= 32'h3a2e3d6e;
    11'b00110010000: data <= 32'hba343d68;
    11'b00110010001: data <= 32'hc0e73015;
    11'b00110010010: data <= 32'hc069b950;
    11'b00110010011: data <= 32'hb8192d4f;
    11'b00110010100: data <= 32'h399f3c73;
    11'b00110010101: data <= 32'h3b2339c7;
    11'b00110010110: data <= 32'h3c08b6e3;
    11'b00110010111: data <= 32'h3d51b34f;
    11'b00110011000: data <= 32'h3c0e3df8;
    11'b00110011001: data <= 32'ha3f040c5;
    11'b00110011010: data <= 32'hb78b3b6f;
    11'b00110011011: data <= 32'h3438bd72;
    11'b00110011100: data <= 32'h3b76c04b;
    11'b00110011101: data <= 32'h3604bd7d;
    11'b00110011110: data <= 32'hb6e2b9b2;
    11'b00110011111: data <= 32'h304cba1d;
    11'b00110100000: data <= 32'h3de1b89c;
    11'b00110100001: data <= 32'h3d25328c;
    11'b00110100010: data <= 32'hbb713878;
    11'b00110100011: data <= 32'hc1aea86c;
    11'b00110100100: data <= 32'hc0d2b847;
    11'b00110100101: data <= 32'hb8dcae28;
    11'b00110100110: data <= 32'h3489365e;
    11'b00110100111: data <= 32'had4eaf67;
    11'b00110101000: data <= 32'hb284b9f7;
    11'b00110101001: data <= 32'h38013293;
    11'b00110101010: data <= 32'h3b324092;
    11'b00110101011: data <= 32'h34f841ff;
    11'b00110101100: data <= 32'hb4df3d0e;
    11'b00110101101: data <= 32'haaa4bb67;
    11'b00110101110: data <= 32'h36b9bd22;
    11'b00110101111: data <= 32'h3471b490;
    11'b00110110000: data <= 32'h32639cfd;
    11'b00110110001: data <= 32'h3cc1baac;
    11'b00110110010: data <= 32'h40b6bcd0;
    11'b00110110011: data <= 32'h3ef3b5b5;
    11'b00110110100: data <= 32'hb90937a2;
    11'b00110110101: data <= 32'hc09031c6;
    11'b00110110110: data <= 32'hbe85b8be;
    11'b00110110111: data <= 32'hb065ba59;
    11'b00110111000: data <= 32'ha4e0b9c7;
    11'b00110111001: data <= 32'hbc16bc4a;
    11'b00110111010: data <= 32'hbc8bbca8;
    11'b00110111011: data <= 32'h2e2530de;
    11'b00110111100: data <= 32'h3b80404e;
    11'b00110111101: data <= 32'h33a6414d;
    11'b00110111110: data <= 32'hbb4a3c60;
    11'b00110111111: data <= 32'hbc38b6d9;
    11'b00111000000: data <= 32'hb6b4b064;
    11'b00111000001: data <= 32'h281b3b3a;
    11'b00111000010: data <= 32'h375338ce;
    11'b00111000011: data <= 32'h3e03baca;
    11'b00111000100: data <= 32'h40eabd31;
    11'b00111000101: data <= 32'h3f6fa297;
    11'b00111000110: data <= 32'ha7b13ce1;
    11'b00111000111: data <= 32'hbc6c3a4e;
    11'b00111001000: data <= 32'hb61eb8c1;
    11'b00111001001: data <= 32'h3819bd79;
    11'b00111001010: data <= 32'hb080bdac;
    11'b00111001011: data <= 32'hbdb2be1b;
    11'b00111001100: data <= 32'hbcc8bde8;
    11'b00111001101: data <= 32'h37d1b6bf;
    11'b00111001110: data <= 32'h3d2e3c8d;
    11'b00111001111: data <= 32'h26a43e3f;
    11'b00111010000: data <= 32'hbee83890;
    11'b00111010001: data <= 32'hc004af15;
    11'b00111010010: data <= 32'hbc4038f7;
    11'b00111010011: data <= 32'hb4d93da7;
    11'b00111010100: data <= 32'h2bba38ab;
    11'b00111010101: data <= 32'h3a62bc07;
    11'b00111010110: data <= 32'h3ec1bc05;
    11'b00111010111: data <= 32'h3e5d3b09;
    11'b00111011000: data <= 32'h3830408a;
    11'b00111011001: data <= 32'ha8e93dd4;
    11'b00111011010: data <= 32'h380eb66f;
    11'b00111011011: data <= 32'h3a70bd2a;
    11'b00111011100: data <= 32'hb24dbc7f;
    11'b00111011101: data <= 32'hbcdfbc94;
    11'b00111011110: data <= 32'hb6ffbe00;
    11'b00111011111: data <= 32'h3dccbcbd;
    11'b00111100000: data <= 32'h3f71b017;
    11'b00111100001: data <= 32'ha59c374e;
    11'b00111100010: data <= 32'hc0192fb9;
    11'b00111100011: data <= 32'hc055a747;
    11'b00111100100: data <= 32'hbc2d3934;
    11'b00111100101: data <= 32'hb8573bcf;
    11'b00111100110: data <= 32'hba68af94;
    11'b00111100111: data <= 32'hb81abd87;
    11'b00111101000: data <= 32'h3876b9b9;
    11'b00111101001: data <= 32'h3cb23e48;
    11'b00111101010: data <= 32'h3a3241ac;
    11'b00111101011: data <= 32'h353a3ee2;
    11'b00111101100: data <= 32'h37d0adeb;
    11'b00111101101: data <= 32'h374ab81d;
    11'b00111101110: data <= 32'hb59f2abc;
    11'b00111101111: data <= 32'hba16b0f7;
    11'b00111110000: data <= 32'h37b8bd10;
    11'b00111110001: data <= 32'h4093bedc;
    11'b00111110010: data <= 32'h4090bb00;
    11'b00111110011: data <= 32'h32a82bc3;
    11'b00111110100: data <= 32'hbe2f3074;
    11'b00111110101: data <= 32'hbd38a9ad;
    11'b00111110110: data <= 32'hb51930a9;
    11'b00111110111: data <= 32'hb86b2558;
    11'b00111111000: data <= 32'hbe85bc19;
    11'b00111111001: data <= 32'hbe7abf3d;
    11'b00111111010: data <= 32'hb195ba03;
    11'b00111111011: data <= 32'h3bda3ddc;
    11'b00111111100: data <= 32'h39c740d7;
    11'b00111111101: data <= 32'hacd73d52;
    11'b00111111110: data <= 32'hb519305f;
    11'b00111111111: data <= 32'hb528382c;
    11'b01000000000: data <= 32'hb9163d9e;
    11'b01000000001: data <= 32'hb84a3a4b;
    11'b01000000010: data <= 32'h3a5bbc13;
    11'b01000000011: data <= 32'h40abbf35;
    11'b01000000100: data <= 32'h4072b9ea;
    11'b01000000101: data <= 32'h3896389e;
    11'b01000000110: data <= 32'hb7973953;
    11'b01000000111: data <= 32'h2e4221e8;
    11'b01000001000: data <= 32'h395bb59a;
    11'b01000001001: data <= 32'hb63cb924;
    11'b01000001010: data <= 32'hc000bdc1;
    11'b01000001011: data <= 32'hbf8dbff6;
    11'b01000001100: data <= 32'ha8d3bc89;
    11'b01000001101: data <= 32'h3cea3853;
    11'b01000001110: data <= 32'h38913cbf;
    11'b01000001111: data <= 32'hba343796;
    11'b01000010000: data <= 32'hbcd730ff;
    11'b01000010001: data <= 32'hbb803cea;
    11'b01000010010: data <= 32'hbb1f4040;
    11'b01000010011: data <= 32'hba563c37;
    11'b01000010100: data <= 32'h3151bc23;
    11'b01000010101: data <= 32'h3dc1be41;
    11'b01000010110: data <= 32'h3e912160;
    11'b01000010111: data <= 32'h3a9c3e24;
    11'b01000011000: data <= 32'h38393d3f;
    11'b01000011001: data <= 32'h3ccc3164;
    11'b01000011010: data <= 32'h3d19b5cd;
    11'b01000011011: data <= 32'hb442b686;
    11'b01000011100: data <= 32'hbf59bb9d;
    11'b01000011101: data <= 32'hbd2cbeec;
    11'b01000011110: data <= 32'h3a66be6d;
    11'b01000011111: data <= 32'h3f11b936;
    11'b01000100000: data <= 32'h3831b030;
    11'b01000100001: data <= 32'hbc8eb505;
    11'b01000100010: data <= 32'hbda125c6;
    11'b01000100011: data <= 32'hbab53d24;
    11'b01000100100: data <= 32'hbb1b3f7b;
    11'b01000100101: data <= 32'hbd8b3812;
    11'b01000100110: data <= 32'hbc45bd7a;
    11'b01000100111: data <= 32'h2e74bd34;
    11'b01000101000: data <= 32'h3af4399a;
    11'b01000101001: data <= 32'h3aa1403e;
    11'b01000101010: data <= 32'h3b3b3e11;
    11'b01000101011: data <= 32'h3d86348d;
    11'b01000101100: data <= 32'h3c7b31c7;
    11'b01000101101: data <= 32'hb5c6398c;
    11'b01000101110: data <= 32'hbdb13379;
    11'b01000101111: data <= 32'hb695bc8b;
    11'b01000110000: data <= 32'h3e8ebf74;
    11'b01000110001: data <= 32'h404ebd91;
    11'b01000110010: data <= 32'h38dfb9f5;
    11'b01000110011: data <= 32'hbaa5b841;
    11'b01000110100: data <= 32'hb8edad58;
    11'b01000110101: data <= 32'h2c2f3aa5;
    11'b01000110110: data <= 32'hb8613be5;
    11'b01000110111: data <= 32'hbfb8b607;
    11'b01000111000: data <= 32'hc04fbf1c;
    11'b01000111001: data <= 32'hbae7bcf4;
    11'b01000111010: data <= 32'h365d39fd;
    11'b01000111011: data <= 32'h39303f13;
    11'b01000111100: data <= 32'h38693bc4;
    11'b01000111101: data <= 32'h396f31ec;
    11'b01000111110: data <= 32'h36423b76;
    11'b01000111111: data <= 32'hb9164009;
    11'b01001000000: data <= 32'hbc913daa;
    11'b01001000001: data <= 32'h2451b896;
    11'b01001000010: data <= 32'h3efbbf23;
    11'b01001000011: data <= 32'h3fddbd34;
    11'b01001000100: data <= 32'h396cb5d5;
    11'b01001000101: data <= 32'ha7e4add5;
    11'b01001000110: data <= 32'h3a08a907;
    11'b01001000111: data <= 32'h3d313505;
    11'b01001001000: data <= 32'ha95d33d8;
    11'b01001001001: data <= 32'hc032bac6;
    11'b01001001010: data <= 32'hc0eabf75;
    11'b01001001011: data <= 32'hbb25bd75;
    11'b01001001100: data <= 32'h38212d00;
    11'b01001001101: data <= 32'h37873892;
    11'b01001001110: data <= 32'hb099b015;
    11'b01001001111: data <= 32'hb40cb0f5;
    11'b01001010000: data <= 32'hb45c3da6;
    11'b01001010001: data <= 32'hbaa14188;
    11'b01001010010: data <= 32'hbcbe3f84;
    11'b01001010011: data <= 32'hb617b69c;
    11'b01001010100: data <= 32'h3b22bdf9;
    11'b01001010101: data <= 32'h3c9db892;
    11'b01001010110: data <= 32'h388638c7;
    11'b01001010111: data <= 32'h39d038b4;
    11'b01001011000: data <= 32'h3f852d59;
    11'b01001011001: data <= 32'h40413061;
    11'b01001011010: data <= 32'h34db346a;
    11'b01001011011: data <= 32'hbf69b692;
    11'b01001011100: data <= 32'hbf92bd96;
    11'b01001011101: data <= 32'had96bdeb;
    11'b01001011110: data <= 32'h3c42badf;
    11'b01001011111: data <= 32'h3680ba25;
    11'b01001100000: data <= 32'hb907bca8;
    11'b01001100001: data <= 32'hb8ffb872;
    11'b01001100010: data <= 32'hb3783d6a;
    11'b01001100011: data <= 32'hb9354118;
    11'b01001100100: data <= 32'hbdc73d9c;
    11'b01001100101: data <= 32'hbd6eb9d4;
    11'b01001100110: data <= 32'hb767bce0;
    11'b01001100111: data <= 32'h2f413285;
    11'b01001101000: data <= 32'h342a3d50;
    11'b01001101001: data <= 32'h3ba73ae2;
    11'b01001101010: data <= 32'h40362bb1;
    11'b01001101011: data <= 32'h40293609;
    11'b01001101100: data <= 32'h34483c81;
    11'b01001101101: data <= 32'hbdb03a42;
    11'b01001101110: data <= 32'hbba3b838;
    11'b01001101111: data <= 32'h3af0bd98;
    11'b01001110000: data <= 32'h3e13bdb4;
    11'b01001110001: data <= 32'h3631bdbb;
    11'b01001110010: data <= 32'hb8afbe24;
    11'b01001110011: data <= 32'hacb1ba22;
    11'b01001110100: data <= 32'h39553af7;
    11'b01001110101: data <= 32'ha96d3e87;
    11'b01001110110: data <= 32'hbe8936e7;
    11'b01001110111: data <= 32'hc07fbcd0;
    11'b01001111000: data <= 32'hbdeebc55;
    11'b01001111001: data <= 32'hb86f37af;
    11'b01001111010: data <= 32'hace63cce;
    11'b01001111011: data <= 32'h3872354f;
    11'b01001111100: data <= 32'h3d94b4a1;
    11'b01001111101: data <= 32'h3d363a2f;
    11'b01001111110: data <= 32'hac18407a;
    11'b01001111111: data <= 32'hbc5f400c;
    11'b01010000000: data <= 32'hb557344c;
    11'b01010000001: data <= 32'h3cbfbc70;
    11'b01010000010: data <= 32'h3d79bd0b;
    11'b01010000011: data <= 32'h3367bc41;
    11'b01010000100: data <= 32'hb039bc5a;
    11'b01010000101: data <= 32'h3c50b981;
    11'b01010000110: data <= 32'h3fd53529;
    11'b01010000111: data <= 32'h39cd39d9;
    11'b01010001000: data <= 32'hbe30b39b;
    11'b01010001001: data <= 32'hc0e7bd5f;
    11'b01010001010: data <= 32'hbe2cbc10;
    11'b01010001011: data <= 32'hb7a43072;
    11'b01010001100: data <= 32'hb413333b;
    11'b01010001101: data <= 32'hb140ba92;
    11'b01010001110: data <= 32'h355cbb46;
    11'b01010001111: data <= 32'h37543bb1;
    11'b01010010000: data <= 32'hb53e41ba;
    11'b01010010001: data <= 32'hbbd74111;
    11'b01010010010: data <= 32'hb6c8382c;
    11'b01010010011: data <= 32'h3877ba33;
    11'b01010010100: data <= 32'h3815b805;
    11'b01010010101: data <= 32'hb15b9dd2;
    11'b01010010110: data <= 32'h34f5b40c;
    11'b01010010111: data <= 32'h4021b7c0;
    11'b01010011000: data <= 32'h41b42637;
    11'b01010011001: data <= 32'h3cdb37b1;
    11'b01010011010: data <= 32'hbcd5a7ac;
    11'b01010011011: data <= 32'hbf63bacc;
    11'b01010011100: data <= 32'hb959bacd;
    11'b01010011101: data <= 32'h3233b779;
    11'b01010011110: data <= 32'hb3afbbae;
    11'b01010011111: data <= 32'hb9edbfc3;
    11'b01010100000: data <= 32'hb4a0be01;
    11'b01010100001: data <= 32'h34463a19;
    11'b01010100010: data <= 32'hb0c2412f;
    11'b01010100011: data <= 32'hbbcd4009;
    11'b01010100100: data <= 32'hbc412fe3;
    11'b01010100101: data <= 32'hb90bb884;
    11'b01010100110: data <= 32'hb8fc357f;
    11'b01010100111: data <= 32'hb9a53b9a;
    11'b01010101000: data <= 32'h35a533ea;
    11'b01010101001: data <= 32'h4073b7b5;
    11'b01010101010: data <= 32'h41982769;
    11'b01010101011: data <= 32'h3c913bfa;
    11'b01010101100: data <= 32'hba8a3bdf;
    11'b01010101101: data <= 32'hbac92f54;
    11'b01010101110: data <= 32'h37beb807;
    11'b01010101111: data <= 32'h3af4ba73;
    11'b01010110000: data <= 32'hb2b7be31;
    11'b01010110001: data <= 32'hbb36c0ab;
    11'b01010110010: data <= 32'habdebeeb;
    11'b01010110011: data <= 32'h3bcc3492;
    11'b01010110100: data <= 32'h385d3e7e;
    11'b01010110101: data <= 32'hbb0c3aff;
    11'b01010110110: data <= 32'hbec5b87a;
    11'b01010110111: data <= 32'hbe3fb7ec;
    11'b01010111000: data <= 32'hbd633a5a;
    11'b01010111001: data <= 32'hbc793c88;
    11'b01010111010: data <= 32'had37acdb;
    11'b01010111011: data <= 32'h3dd9bb31;
    11'b01010111100: data <= 32'h3f823069;
    11'b01010111101: data <= 32'h38fc3f4c;
    11'b01010111110: data <= 32'hb881403f;
    11'b01010111111: data <= 32'had113bf6;
    11'b01011000000: data <= 32'h3c66ad3d;
    11'b01011000001: data <= 32'h3b7db880;
    11'b01011000010: data <= 32'hb68dbc84;
    11'b01011000011: data <= 32'hb9d1bf21;
    11'b01011000100: data <= 32'h3a53bdfc;
    11'b01011000101: data <= 32'h404eb209;
    11'b01011000110: data <= 32'h3dab38c4;
    11'b01011000111: data <= 32'hb8e4acf7;
    11'b01011001000: data <= 32'hbf17bb71;
    11'b01011001001: data <= 32'hbe48b696;
    11'b01011001010: data <= 32'hbcd339bc;
    11'b01011001011: data <= 32'hbcbf3775;
    11'b01011001100: data <= 32'hb9ebbc6a;
    11'b01011001101: data <= 32'h34b7be88;
    11'b01011001110: data <= 32'h3a212ea5;
    11'b01011001111: data <= 32'h2f9f4093;
    11'b01011010000: data <= 32'hb7644129;
    11'b01011010001: data <= 32'h2cdd3ce8;
    11'b01011010010: data <= 32'h3a493258;
    11'b01011010011: data <= 32'h3314310f;
    11'b01011010100: data <= 32'hbb6325e2;
    11'b01011010101: data <= 32'hb848b9a4;
    11'b01011010110: data <= 32'h3e54bc35;
    11'b01011010111: data <= 32'h41fcb734;
    11'b01011011000: data <= 32'h3fb42fc7;
    11'b01011011001: data <= 32'hb44eb20c;
    11'b01011011010: data <= 32'hbcb1b8ce;
    11'b01011011011: data <= 32'hb8e9b07c;
    11'b01011011100: data <= 32'hb52d360f;
    11'b01011011101: data <= 32'hbb8db800;
    11'b01011011110: data <= 32'hbd0cc055;
    11'b01011011111: data <= 32'hb840c091;
    11'b01011100000: data <= 32'h340fb0fc;
    11'b01011100001: data <= 32'h2ee93ff2;
    11'b01011100010: data <= 32'hb5ef3ff7;
    11'b01011100011: data <= 32'hb49e3939;
    11'b01011100100: data <= 32'hb11b3290;
    11'b01011100101: data <= 32'hbad13b8e;
    11'b01011100110: data <= 32'hbe373ca4;
    11'b01011100111: data <= 32'hb8d82f59;
    11'b01011101000: data <= 32'h3eb7baac;
    11'b01011101001: data <= 32'h41c0b807;
    11'b01011101010: data <= 32'h3ee135d2;
    11'b01011101011: data <= 32'ha9cf387b;
    11'b01011101100: data <= 32'hb35b34aa;
    11'b01011101101: data <= 32'h39a1352a;
    11'b01011101110: data <= 32'h394f3266;
    11'b01011101111: data <= 32'hb96fbbf2;
    11'b01011110000: data <= 32'hbdcfc106;
    11'b01011110001: data <= 32'hb88ec0da;
    11'b01011110010: data <= 32'h396ab814;
    11'b01011110011: data <= 32'h39af3c3c;
    11'b01011110100: data <= 32'hb0ce3995;
    11'b01011110101: data <= 32'hb9beb544;
    11'b01011110110: data <= 32'hbbbd27ca;
    11'b01011110111: data <= 32'hbe293d99;
    11'b01011111000: data <= 32'hbfba3e65;
    11'b01011111001: data <= 32'hbbc12def;
    11'b01011111010: data <= 32'h3b87bc88;
    11'b01011111011: data <= 32'h3f47b826;
    11'b01011111100: data <= 32'h3b623bb6;
    11'b01011111101: data <= 32'ha8843e31;
    11'b01011111110: data <= 32'h38363c94;
    11'b01011111111: data <= 32'h3e423a16;
    11'b01100000000: data <= 32'h3c3036da;
    11'b01100000001: data <= 32'hb9dab8a0;
    11'b01100000010: data <= 32'hbd8ebf61;
    11'b01100000011: data <= 32'h28e9bfc8;
    11'b01100000100: data <= 32'h3eb5ba02;
    11'b01100000101: data <= 32'h3e3a2b11;
    11'b01100000110: data <= 32'h31b6b7d7;
    11'b01100000111: data <= 32'hba11bc1e;
    11'b01100001000: data <= 32'hbba8ac00;
    11'b01100001001: data <= 32'hbd3d3da8;
    11'b01100001010: data <= 32'hbf303cbe;
    11'b01100001011: data <= 32'hbdacb9d8;
    11'b01100001100: data <= 32'hb24ebf58;
    11'b01100001101: data <= 32'h37bfb925;
    11'b01100001110: data <= 32'h2d163d5b;
    11'b01100001111: data <= 32'hb06e3fda;
    11'b01100010000: data <= 32'h3a073d3e;
    11'b01100010001: data <= 32'h3e0c3b1a;
    11'b01100010010: data <= 32'h38803bce;
    11'b01100010011: data <= 32'hbccd385d;
    11'b01100010100: data <= 32'hbd3ab875;
    11'b01100010101: data <= 32'h399ebca5;
    11'b01100010110: data <= 32'h40e7ba48;
    11'b01100010111: data <= 32'h400bb788;
    11'b01100011000: data <= 32'h36c2baf6;
    11'b01100011001: data <= 32'hb499bbad;
    11'b01100011010: data <= 32'ha582308a;
    11'b01100011011: data <= 32'hb38e3cc9;
    11'b01100011100: data <= 32'hbce63617;
    11'b01100011101: data <= 32'hbecdbed5;
    11'b01100011110: data <= 32'hbc39c0ec;
    11'b01100011111: data <= 32'hb4d3bada;
    11'b01100100000: data <= 32'hb31d3c79;
    11'b01100100001: data <= 32'hb09f3d88;
    11'b01100100010: data <= 32'h38133891;
    11'b01100100011: data <= 32'h3a0c38bd;
    11'b01100100100: data <= 32'hb6753e18;
    11'b01100100101: data <= 32'hbf493ece;
    11'b01100100110: data <= 32'hbd84384a;
    11'b01100100111: data <= 32'h3aaab8fd;
    11'b01100101000: data <= 32'h40abb9a9;
    11'b01100101001: data <= 32'h3eb6b578;
    11'b01100101010: data <= 32'h3616b55f;
    11'b01100101011: data <= 32'h36ecb276;
    11'b01100101100: data <= 32'h3d3a38ce;
    11'b01100101101: data <= 32'h3c163c3d;
    11'b01100101110: data <= 32'hb8f5aead;
    11'b01100101111: data <= 32'hbee7c017;
    11'b01100110000: data <= 32'hbcc7c0ff;
    11'b01100110001: data <= 32'haf63bbeb;
    11'b01100110010: data <= 32'h32c7363b;
    11'b01100110011: data <= 32'h2c3d2d38;
    11'b01100110100: data <= 32'h30f3b964;
    11'b01100110101: data <= 32'h99552c34;
    11'b01100110110: data <= 32'hbc4d3f26;
    11'b01100110111: data <= 32'hc0414073;
    11'b01100111000: data <= 32'hbe493a2a;
    11'b01100111001: data <= 32'h3438b9bc;
    11'b01100111010: data <= 32'h3d17b98c;
    11'b01100111011: data <= 32'h390d3137;
    11'b01100111100: data <= 32'h28e33886;
    11'b01100111101: data <= 32'h3bd738fc;
    11'b01100111110: data <= 32'h407c3bff;
    11'b01100111111: data <= 32'h3eb73caf;
    11'b01101000000: data <= 32'hb6d7319e;
    11'b01101000001: data <= 32'hbe6cbd80;
    11'b01101000010: data <= 32'hb989bf29;
    11'b01101000011: data <= 32'h3a1abb1e;
    11'b01101000100: data <= 32'h3c0bb65e;
    11'b01101000101: data <= 32'h3616bcb3;
    11'b01101000110: data <= 32'h2a44bea7;
    11'b01101000111: data <= 32'hadd4b4f1;
    11'b01101001000: data <= 32'hbac43edd;
    11'b01101001001: data <= 32'hbf303faf;
    11'b01101001010: data <= 32'hbed12e73;
    11'b01101001011: data <= 32'hb946bd63;
    11'b01101001100: data <= 32'hb008ba88;
    11'b01101001101: data <= 32'hb81b3876;
    11'b01101001110: data <= 32'hb6133c2a;
    11'b01101001111: data <= 32'h3c5d3a5c;
    11'b01101010000: data <= 32'h40993bc4;
    11'b01101010001: data <= 32'h3d833dc2;
    11'b01101010010: data <= 32'hba573c60;
    11'b01101010011: data <= 32'hbe19a82b;
    11'b01101010100: data <= 32'ha9abb99a;
    11'b01101010101: data <= 32'h3e41b8aa;
    11'b01101010110: data <= 32'h3defba40;
    11'b01101010111: data <= 32'h3813bea9;
    11'b01101011000: data <= 32'h3499bf3e;
    11'b01101011001: data <= 32'h3942b3da;
    11'b01101011010: data <= 32'h345c3df5;
    11'b01101011011: data <= 32'hbb6c3ca3;
    11'b01101011100: data <= 32'hbe86baf5;
    11'b01101011101: data <= 32'hbd69bfe9;
    11'b01101011110: data <= 32'hbc17bb9e;
    11'b01101011111: data <= 32'hbc45382a;
    11'b01101100000: data <= 32'hb88e3902;
    11'b01101100001: data <= 32'h3a972552;
    11'b01101100010: data <= 32'h3e6f365c;
    11'b01101100011: data <= 32'h373f3e88;
    11'b01101100100: data <= 32'hbda54024;
    11'b01101100101: data <= 32'hbe333caf;
    11'b01101100110: data <= 32'h33302fbb;
    11'b01101100111: data <= 32'h3e58b468;
    11'b01101101000: data <= 32'h3c78b8da;
    11'b01101101001: data <= 32'h32ffbcdb;
    11'b01101101010: data <= 32'h3958bc86;
    11'b01101101011: data <= 32'h3f333247;
    11'b01101101100: data <= 32'h3e8d3d52;
    11'b01101101101: data <= 32'ha36e38a1;
    11'b01101101110: data <= 32'hbd88bd4b;
    11'b01101101111: data <= 32'hbdaec003;
    11'b01101110000: data <= 32'hbb7cbafb;
    11'b01101110001: data <= 32'hba042ec2;
    11'b01101110010: data <= 32'hb670b7de;
    11'b01101110011: data <= 32'h375fbd4e;
    11'b01101110100: data <= 32'h3a57b738;
    11'b01101110101: data <= 32'hb5023e5b;
    11'b01101110110: data <= 32'hbee740fe;
    11'b01101110111: data <= 32'hbe473e11;
    11'b01101111000: data <= 32'hac0e3220;
    11'b01101111001: data <= 32'h399cb1ca;
    11'b01101111010: data <= 32'ha5e3ae2c;
    11'b01101111011: data <= 32'hb72db4a3;
    11'b01101111100: data <= 32'h3b17b39b;
    11'b01101111101: data <= 32'h413d38ec;
    11'b01101111110: data <= 32'h40d63d3e;
    11'b01101111111: data <= 32'h362c38e8;
    11'b01110000000: data <= 32'hbc8eba97;
    11'b01110000001: data <= 32'hbb3cbcdf;
    11'b01110000010: data <= 32'hac31b74a;
    11'b01110000011: data <= 32'h2d4db57a;
    11'b01110000100: data <= 32'hac1abe79;
    11'b01110000101: data <= 32'h3435c0e6;
    11'b01110000110: data <= 32'h37f6bc4d;
    11'b01110000111: data <= 32'hb3e83d63;
    11'b01110001000: data <= 32'hbd574054;
    11'b01110001001: data <= 32'hbd9f3b0e;
    11'b01110001010: data <= 32'hb92eb6fd;
    11'b01110001011: data <= 32'hb878b51f;
    11'b01110001100: data <= 32'hbd3f35c1;
    11'b01110001101: data <= 32'hbc9c35a9;
    11'b01110001110: data <= 32'h3a442da4;
    11'b01110001111: data <= 32'h4144386a;
    11'b01110010000: data <= 32'h405b3d41;
    11'b01110010001: data <= 32'h2c2c3ccf;
    11'b01110010010: data <= 32'hbc3735fb;
    11'b01110010011: data <= 32'hb2e424da;
    11'b01110010100: data <= 32'h3aee3157;
    11'b01110010101: data <= 32'h3992b792;
    11'b01110010110: data <= 32'h2b12c01b;
    11'b01110010111: data <= 32'h3465c15f;
    11'b01110011000: data <= 32'h3b7dbc69;
    11'b01110011001: data <= 32'h39c33c5a;
    11'b01110011010: data <= 32'hb52f3d7d;
    11'b01110011011: data <= 32'hbbfdb1fa;
    11'b01110011100: data <= 32'hbc3abcc4;
    11'b01110011101: data <= 32'hbd8db775;
    11'b01110011110: data <= 32'hbfec3812;
    11'b01110011111: data <= 32'hbdf13322;
    11'b01110100000: data <= 32'h3728b83d;
    11'b01110100001: data <= 32'h3faab0b5;
    11'b01110100010: data <= 32'h3cbd3cae;
    11'b01110100011: data <= 32'hb93d3f7e;
    11'b01110100100: data <= 32'hbc673dff;
    11'b01110100101: data <= 32'h32823bdb;
    11'b01110100110: data <= 32'h3c95395e;
    11'b01110100111: data <= 32'h37d9b20a;
    11'b01110101000: data <= 32'hb56abe4d;
    11'b01110101001: data <= 32'h354dbfe3;
    11'b01110101010: data <= 32'h3f0db8b7;
    11'b01110101011: data <= 32'h3ffc3ba3;
    11'b01110101100: data <= 32'h3a013961;
    11'b01110101101: data <= 32'hb809bafa;
    11'b01110101110: data <= 32'hbbc4bd88;
    11'b01110101111: data <= 32'hbd17b4f4;
    11'b01110110000: data <= 32'hbeae3653;
    11'b01110110001: data <= 32'hbd25b8a3;
    11'b01110110010: data <= 32'h2e9fbf1e;
    11'b01110110011: data <= 32'h3c05bcac;
    11'b01110110100: data <= 32'h32d93abb;
    11'b01110110101: data <= 32'hbc894036;
    11'b01110110110: data <= 32'hbc4a3f41;
    11'b01110110111: data <= 32'h320b3c63;
    11'b01110111000: data <= 32'h38913a44;
    11'b01110111001: data <= 32'hb8593521;
    11'b01110111010: data <= 32'hbcb7b8a0;
    11'b01110111011: data <= 32'h339bbb36;
    11'b01110111100: data <= 32'h40b69f8f;
    11'b01110111101: data <= 32'h417b3b51;
    11'b01110111110: data <= 32'h3cf0376f;
    11'b01110111111: data <= 32'hb1f5b961;
    11'b01111000000: data <= 32'hb6d5b9b5;
    11'b01111000001: data <= 32'hb5833460;
    11'b01111000010: data <= 32'hb988345e;
    11'b01111000011: data <= 32'hba5dbdd2;
    11'b01111000100: data <= 32'haddbc1bb;
    11'b01111000101: data <= 32'h37febfa6;
    11'b01111000110: data <= 32'ha19c3781;
    11'b01111000111: data <= 32'hbb063ed8;
    11'b01111001000: data <= 32'hba133c85;
    11'b01111001001: data <= 32'hac4335ce;
    11'b01111001010: data <= 32'hb6c2381f;
    11'b01111001011: data <= 32'hbf2b3a15;
    11'b01111001100: data <= 32'hc01233db;
    11'b01111001101: data <= 32'haa29b4c1;
    11'b01111001110: data <= 32'h408a2d3d;
    11'b01111001111: data <= 32'h40ec3a5b;
    11'b01111010000: data <= 32'h3acc39dc;
    11'b01111010001: data <= 32'hb23d33de;
    11'b01111010010: data <= 32'h33d837aa;
    11'b01111010011: data <= 32'h39ed3c4b;
    11'b01111010100: data <= 32'h31e235f2;
    11'b01111010101: data <= 32'hb811bf08;
    11'b01111010110: data <= 32'hb174c223;
    11'b01111010111: data <= 32'h3910bfaf;
    11'b01111011000: data <= 32'h39583428;
    11'b01111011001: data <= 32'h2ce13b65;
    11'b01111011010: data <= 32'hb126ac7e;
    11'b01111011011: data <= 32'hb2afb910;
    11'b01111011100: data <= 32'hbc5c3230;
    11'b01111011101: data <= 32'hc0e23bc1;
    11'b01111011110: data <= 32'hc0cc365c;
    11'b01111011111: data <= 32'hb628b8f7;
    11'b01111100000: data <= 32'h3e2ab857;
    11'b01111100001: data <= 32'h3d6c3759;
    11'b01111100010: data <= 32'had7e3c6e;
    11'b01111100011: data <= 32'hb6ac3cbc;
    11'b01111100100: data <= 32'h39973dbc;
    11'b01111100101: data <= 32'h3d1e3ea0;
    11'b01111100110: data <= 32'h346739b1;
    11'b01111100111: data <= 32'hba70bcfe;
    11'b01111101000: data <= 32'hb4b3c086;
    11'b01111101001: data <= 32'h3c9abce5;
    11'b01111101010: data <= 32'h3ef034a3;
    11'b01111101011: data <= 32'h3c973298;
    11'b01111101100: data <= 32'h3752bbf3;
    11'b01111101101: data <= 32'ha196bc7d;
    11'b01111101110: data <= 32'hbb5c334e;
    11'b01111101111: data <= 32'hc01e3c0e;
    11'b01111110000: data <= 32'hc01cade7;
    11'b01111110001: data <= 32'hb8b3be91;
    11'b01111110010: data <= 32'h38f9be3c;
    11'b01111110011: data <= 32'h314ba7ac;
    11'b01111110100: data <= 32'hbae63cb6;
    11'b01111110101: data <= 32'hb8433dab;
    11'b01111110110: data <= 32'h3a8b3e01;
    11'b01111110111: data <= 32'h3c0e3eb5;
    11'b01111111000: data <= 32'hb81c3c74;
    11'b01111111001: data <= 32'hbe88b3cb;
    11'b01111111010: data <= 32'hb88fbbf1;
    11'b01111111011: data <= 32'h3e25b599;
    11'b01111111100: data <= 32'h40bf369c;
    11'b01111111101: data <= 32'h3e6eaf08;
    11'b01111111110: data <= 32'h39ebbc63;
    11'b01111111111: data <= 32'h378bb9b5;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    