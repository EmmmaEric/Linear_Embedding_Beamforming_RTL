
module memory_rom_47(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3c6d3c82;
    11'b00000000001: data <= 32'h398538e3;
    11'b00000000010: data <= 32'hb8ebb94a;
    11'b00000000011: data <= 32'hb8bcbf1a;
    11'b00000000100: data <= 32'h3c53bd5d;
    11'b00000000101: data <= 32'h40af3054;
    11'b00000000110: data <= 32'h3f0d38f9;
    11'b00000000111: data <= 32'h34f8b71d;
    11'b00000001000: data <= 32'hb842bcf7;
    11'b00000001001: data <= 32'hbacab6a6;
    11'b00000001010: data <= 32'hbd74398c;
    11'b00000001011: data <= 32'hbe9d2d48;
    11'b00000001100: data <= 32'hbafcbec3;
    11'b00000001101: data <= 32'h3579c04b;
    11'b00000001110: data <= 32'h3726b740;
    11'b00000001111: data <= 32'hb86c3dfe;
    11'b00000010000: data <= 32'hbb6c3fa8;
    11'b00000010001: data <= 32'h26463d3a;
    11'b00000010010: data <= 32'h39973c09;
    11'b00000010011: data <= 32'hb4863b93;
    11'b00000010100: data <= 32'hbe7234b1;
    11'b00000010101: data <= 32'hbc02b8a9;
    11'b00000010110: data <= 32'h3d5db849;
    11'b00000010111: data <= 32'h41a9345c;
    11'b00000011000: data <= 32'h40203701;
    11'b00000011001: data <= 32'h37d8b554;
    11'b00000011010: data <= 32'hab9ab8d5;
    11'b00000011011: data <= 32'h306c353f;
    11'b00000011100: data <= 32'hb18d3b2f;
    11'b00000011101: data <= 32'hbaf1b751;
    11'b00000011110: data <= 32'hba96c121;
    11'b00000011111: data <= 32'haca5c1a0;
    11'b00000100000: data <= 32'h31bdba8d;
    11'b00000100001: data <= 32'hb5553c39;
    11'b00000100010: data <= 32'hb8043c56;
    11'b00000100011: data <= 32'h290334af;
    11'b00000100100: data <= 32'h9daf3652;
    11'b00000100101: data <= 32'hbd883c74;
    11'b00000100110: data <= 32'hc1003c11;
    11'b00000100111: data <= 32'hbdb12ce5;
    11'b00000101000: data <= 32'h3c5db5de;
    11'b00000101001: data <= 32'h40af2fbb;
    11'b00000101010: data <= 32'h3d883844;
    11'b00000101011: data <= 32'h3061361e;
    11'b00000101100: data <= 32'h35a23818;
    11'b00000101101: data <= 32'h3ca53cfa;
    11'b00000101110: data <= 32'h3a943cf5;
    11'b00000101111: data <= 32'hb6aab804;
    11'b00000110000: data <= 32'hbab5c110;
    11'b00000110001: data <= 32'ha1dcc122;
    11'b00000110010: data <= 32'h39f6ba04;
    11'b00000110011: data <= 32'h38e0377c;
    11'b00000110100: data <= 32'h342caf9e;
    11'b00000110101: data <= 32'h31fcbb49;
    11'b00000110110: data <= 32'hb607b24e;
    11'b00000110111: data <= 32'hbf373ca2;
    11'b00000111000: data <= 32'hc15f3ca8;
    11'b00000111001: data <= 32'hbe6bb204;
    11'b00000111010: data <= 32'h3732bc0c;
    11'b00000111011: data <= 32'h3c9eb636;
    11'b00000111100: data <= 32'h314e3908;
    11'b00000111101: data <= 32'hb71b3c31;
    11'b00000111110: data <= 32'h38763d27;
    11'b00000111111: data <= 32'h3e983f00;
    11'b00001000000: data <= 32'h3bc63e40;
    11'b00001000001: data <= 32'hb9ab2a93;
    11'b00001000010: data <= 32'hbc66be3c;
    11'b00001000011: data <= 32'h3469be30;
    11'b00001000100: data <= 32'h3e6eb540;
    11'b00001000101: data <= 32'h3e5c28ab;
    11'b00001000110: data <= 32'h3b40bbd6;
    11'b00001000111: data <= 32'h37d0be02;
    11'b00001001000: data <= 32'haa6fb3f9;
    11'b00001001001: data <= 32'hbcc43d06;
    11'b00001001010: data <= 32'hc0093aaa;
    11'b00001001011: data <= 32'hbdc5bc52;
    11'b00001001100: data <= 32'hb2bbc00f;
    11'b00001001101: data <= 32'h9c54bc03;
    11'b00001001110: data <= 32'hba3e3813;
    11'b00001001111: data <= 32'hba113c44;
    11'b00001010000: data <= 32'h38e63c6d;
    11'b00001010001: data <= 32'h3dd43de9;
    11'b00001010010: data <= 32'h34193eb5;
    11'b00001010011: data <= 32'hbe603b12;
    11'b00001010100: data <= 32'hbe45b3e3;
    11'b00001010101: data <= 32'h36c3b6d1;
    11'b00001010110: data <= 32'h400d2e22;
    11'b00001010111: data <= 32'h3f60ae8d;
    11'b00001011000: data <= 32'h3bd1bc50;
    11'b00001011001: data <= 32'h3a4dbc91;
    11'b00001011010: data <= 32'h3aa535c5;
    11'b00001011011: data <= 32'h2ec53e19;
    11'b00001011100: data <= 32'hbb6a370e;
    11'b00001011101: data <= 32'hbc5ebf67;
    11'b00001011110: data <= 32'hb86fc14d;
    11'b00001011111: data <= 32'hb794bd37;
    11'b00001100000: data <= 32'hbadd31f7;
    11'b00001100001: data <= 32'hb7eb3510;
    11'b00001100010: data <= 32'h397c98d9;
    11'b00001100011: data <= 32'h3b6b38a1;
    11'b00001100100: data <= 32'hb9ad3e2a;
    11'b00001100101: data <= 32'hc0e03e10;
    11'b00001100110: data <= 32'hbfdb38d5;
    11'b00001100111: data <= 32'h33932bb5;
    11'b00001101000: data <= 32'h3e5c3079;
    11'b00001101001: data <= 32'h3c51aa85;
    11'b00001101010: data <= 32'h35e3b873;
    11'b00001101011: data <= 32'h3b49b212;
    11'b00001101100: data <= 32'h3f013ceb;
    11'b00001101101: data <= 32'h3d213f84;
    11'b00001101110: data <= 32'hb092362a;
    11'b00001101111: data <= 32'hbb02bf5c;
    11'b00001110000: data <= 32'hb81ec0aa;
    11'b00001110001: data <= 32'haf3fbc12;
    11'b00001110010: data <= 32'haf02b07b;
    11'b00001110011: data <= 32'h32b9ba45;
    11'b00001110100: data <= 32'h3b02bd82;
    11'b00001110101: data <= 32'h38c0b5aa;
    11'b00001110110: data <= 32'hbc803d4c;
    11'b00001110111: data <= 32'hc1233ea2;
    11'b00001111000: data <= 32'hbfe23868;
    11'b00001111001: data <= 32'hb1b8b5be;
    11'b00001111010: data <= 32'h37f3b4a3;
    11'b00001111011: data <= 32'hb4caa3e0;
    11'b00001111100: data <= 32'hb870277d;
    11'b00001111101: data <= 32'h3aa8386e;
    11'b00001111110: data <= 32'h406c3ec9;
    11'b00001111111: data <= 32'h3e964026;
    11'b00010000000: data <= 32'hb1a83a0c;
    11'b00010000001: data <= 32'hbc1cbb9a;
    11'b00010000010: data <= 32'hb4aabca7;
    11'b00010000011: data <= 32'h3911b42c;
    11'b00010000100: data <= 32'h3a7bb46b;
    11'b00010000101: data <= 32'h3aa5be65;
    11'b00010000110: data <= 32'h3c67c05e;
    11'b00010000111: data <= 32'h3a48b98e;
    11'b00010001000: data <= 32'hb8a83d1c;
    11'b00010001001: data <= 32'hbf123d89;
    11'b00010001010: data <= 32'hbdfbb253;
    11'b00010001011: data <= 32'hb859bd23;
    11'b00010001100: data <= 32'hb8d6bb14;
    11'b00010001101: data <= 32'hbddcaeb0;
    11'b00010001110: data <= 32'hbcbe303e;
    11'b00010001111: data <= 32'h39a536d7;
    11'b00010010000: data <= 32'h40203d44;
    11'b00010010001: data <= 32'h3c623fa2;
    11'b00010010010: data <= 32'hbb813d38;
    11'b00010010011: data <= 32'hbde234c5;
    11'b00010010100: data <= 32'hb0c831ad;
    11'b00010010101: data <= 32'h3c5b380a;
    11'b00010010110: data <= 32'h3c67b25e;
    11'b00010010111: data <= 32'h3a8fbee7;
    11'b00010011000: data <= 32'h3ca6c004;
    11'b00010011001: data <= 32'h3da0b3c9;
    11'b00010011010: data <= 32'h392f3e07;
    11'b00010011011: data <= 32'hb7613c15;
    11'b00010011100: data <= 32'hba48bbb6;
    11'b00010011101: data <= 32'hb920bfb3;
    11'b00010011110: data <= 32'hbc5abc85;
    11'b00010011111: data <= 32'hbefcb39f;
    11'b00010100000: data <= 32'hbc7ab642;
    11'b00010100001: data <= 32'h39beb8eb;
    11'b00010100010: data <= 32'h3e4e32e5;
    11'b00010100011: data <= 32'h316e3da4;
    11'b00010100100: data <= 32'hbf213eab;
    11'b00010100101: data <= 32'hbf563c99;
    11'b00010100110: data <= 32'hb2423b19;
    11'b00010100111: data <= 32'h3ab93a50;
    11'b00010101000: data <= 32'h3665ab2f;
    11'b00010101001: data <= 32'h2752bd04;
    11'b00010101010: data <= 32'h3b79bc84;
    11'b00010101011: data <= 32'h401838d6;
    11'b00010101100: data <= 32'h3f413f60;
    11'b00010101101: data <= 32'h387e3af8;
    11'b00010101110: data <= 32'hb496bc68;
    11'b00010101111: data <= 32'hb791beaa;
    11'b00010110000: data <= 32'hba3bb980;
    11'b00010110001: data <= 32'hbc6ab3a1;
    11'b00010110010: data <= 32'hb76fbcdb;
    11'b00010110011: data <= 32'h3b32bfe1;
    11'b00010110100: data <= 32'h3cc1bbbb;
    11'b00010110101: data <= 32'hb5bb3afc;
    11'b00010110110: data <= 32'hbfe13e92;
    11'b00010110111: data <= 32'hbedb3c92;
    11'b00010111000: data <= 32'hb51a38dc;
    11'b00010111001: data <= 32'h22293724;
    11'b00010111010: data <= 32'hbba3a053;
    11'b00010111011: data <= 32'hbc95b92f;
    11'b00010111100: data <= 32'h3813b4f2;
    11'b00010111101: data <= 32'h409c3c80;
    11'b00010111110: data <= 32'h406f3fc9;
    11'b00010111111: data <= 32'h39993bea;
    11'b00011000000: data <= 32'hb4e7b754;
    11'b00011000001: data <= 32'hb31ab833;
    11'b00011000010: data <= 32'ha8ba3515;
    11'b00011000011: data <= 32'hb09ba2ff;
    11'b00011000100: data <= 32'h3287bf38;
    11'b00011000101: data <= 32'h3c41c1a0;
    11'b00011000110: data <= 32'h3cb0be0a;
    11'b00011000111: data <= 32'ha908392c;
    11'b00011001000: data <= 32'hbcd13d42;
    11'b00011001001: data <= 32'hbc0336a6;
    11'b00011001010: data <= 32'hb51fb524;
    11'b00011001011: data <= 32'hbaccb1d4;
    11'b00011001100: data <= 32'hc04eac1c;
    11'b00011001101: data <= 32'hc004b620;
    11'b00011001110: data <= 32'h30fbb38e;
    11'b00011001111: data <= 32'h40253a55;
    11'b00011010000: data <= 32'h3eca3e46;
    11'b00011010001: data <= 32'ha6fe3cbc;
    11'b00011010010: data <= 32'hba123858;
    11'b00011010011: data <= 32'hac053ac5;
    11'b00011010100: data <= 32'h38503d5c;
    11'b00011010101: data <= 32'h351d355c;
    11'b00011010110: data <= 32'h3402bf44;
    11'b00011010111: data <= 32'h3b95c15a;
    11'b00011011000: data <= 32'h3dd8bc86;
    11'b00011011001: data <= 32'h3b893ad1;
    11'b00011011010: data <= 32'h301b3b83;
    11'b00011011011: data <= 32'ha4eeb6f8;
    11'b00011011100: data <= 32'haedbbc6c;
    11'b00011011101: data <= 32'hbcc1b7e3;
    11'b00011011110: data <= 32'hc0f7ab8a;
    11'b00011011111: data <= 32'hc01db8db;
    11'b00011100000: data <= 32'h2eabbc23;
    11'b00011100001: data <= 32'h3e45b538;
    11'b00011100010: data <= 32'h39b73a53;
    11'b00011100011: data <= 32'hbbe53cd5;
    11'b00011100100: data <= 32'hbcc33ce6;
    11'b00011100101: data <= 32'h9e033e74;
    11'b00011100110: data <= 32'h386b3f22;
    11'b00011100111: data <= 32'hb0b738b5;
    11'b00011101000: data <= 32'hb859bd3f;
    11'b00011101001: data <= 32'h372abf0d;
    11'b00011101010: data <= 32'h3efeb25f;
    11'b00011101011: data <= 32'h3fab3d04;
    11'b00011101100: data <= 32'h3cdd39ba;
    11'b00011101101: data <= 32'h3977ba64;
    11'b00011101110: data <= 32'h331ebc46;
    11'b00011101111: data <= 32'hbaa1ac1c;
    11'b00011110000: data <= 32'hbf51322c;
    11'b00011110001: data <= 32'hbd6abc4d;
    11'b00011110010: data <= 32'h356dc05f;
    11'b00011110011: data <= 32'h3c85be4e;
    11'b00011110100: data <= 32'h9d06222f;
    11'b00011110101: data <= 32'hbd893bc5;
    11'b00011110110: data <= 32'hbc693c94;
    11'b00011110111: data <= 32'h2e183d63;
    11'b00011111000: data <= 32'h2c473dbf;
    11'b00011111001: data <= 32'hbd2938d7;
    11'b00011111010: data <= 32'hbf24b95f;
    11'b00011111011: data <= 32'hb3e2ba43;
    11'b00011111100: data <= 32'h3eff3826;
    11'b00011111101: data <= 32'h40723da3;
    11'b00011111110: data <= 32'h3d8e3923;
    11'b00011111111: data <= 32'h39aeb7b0;
    11'b00100000000: data <= 32'h37a5b093;
    11'b00100000001: data <= 32'hab753c03;
    11'b00100000010: data <= 32'hb9ec39a0;
    11'b00100000011: data <= 32'hb80abd7f;
    11'b00100000100: data <= 32'h3894c1d1;
    11'b00100000101: data <= 32'h3ba7c059;
    11'b00100000110: data <= 32'h213fb507;
    11'b00100000111: data <= 32'hbab238bf;
    11'b00100001000: data <= 32'hb5763628;
    11'b00100001001: data <= 32'h3623351e;
    11'b00100001010: data <= 32'hb7af393a;
    11'b00100001011: data <= 32'hc0b4378a;
    11'b00100001100: data <= 32'hc171b486;
    11'b00100001101: data <= 32'hba03b6e2;
    11'b00100001110: data <= 32'h3dac3689;
    11'b00100001111: data <= 32'h3ea53c00;
    11'b00100010000: data <= 32'h38c03870;
    11'b00100010001: data <= 32'h30613230;
    11'b00100010010: data <= 32'h387d3c53;
    11'b00100010011: data <= 32'h38e6403b;
    11'b00100010100: data <= 32'ha5fa3d00;
    11'b00100010101: data <= 32'hb362bcf5;
    11'b00100010110: data <= 32'h373cc16f;
    11'b00100010111: data <= 32'h3bdabf08;
    11'b00100011000: data <= 32'h3945a7c3;
    11'b00100011001: data <= 32'h35643470;
    11'b00100011010: data <= 32'h39f3b853;
    11'b00100011011: data <= 32'h3aafb986;
    11'b00100011100: data <= 32'hb9092f60;
    11'b00100011101: data <= 32'hc13c373d;
    11'b00100011110: data <= 32'hc187b455;
    11'b00100011111: data <= 32'hba2fbb2f;
    11'b00100100000: data <= 32'h3b91b84b;
    11'b00100100001: data <= 32'h38eb2faa;
    11'b00100100010: data <= 32'hb88534f2;
    11'b00100100011: data <= 32'hb81f392c;
    11'b00100100100: data <= 32'h38903f19;
    11'b00100100101: data <= 32'h3aa4412d;
    11'b00100100110: data <= 32'hb1663e1d;
    11'b00100100111: data <= 32'hbab2b9e1;
    11'b00100101000: data <= 32'hb079befc;
    11'b00100101001: data <= 32'h3bdbb93a;
    11'b00100101010: data <= 32'h3d7f389f;
    11'b00100101011: data <= 32'h3d5e2f8f;
    11'b00100101100: data <= 32'h3e0abc51;
    11'b00100101101: data <= 32'h3cfdbbb5;
    11'b00100101110: data <= 32'hb3593576;
    11'b00100101111: data <= 32'hbfa43a35;
    11'b00100110000: data <= 32'hbfaeb736;
    11'b00100110001: data <= 32'hb5aebf11;
    11'b00100110010: data <= 32'h38a0bec6;
    11'b00100110011: data <= 32'hb418ba03;
    11'b00100110100: data <= 32'hbd09ac57;
    11'b00100110101: data <= 32'hb92737be;
    11'b00100110110: data <= 32'h39bd3dd3;
    11'b00100110111: data <= 32'h38ff4046;
    11'b00100111000: data <= 32'hbc0f3d95;
    11'b00100111001: data <= 32'hbfe5b12c;
    11'b00100111010: data <= 32'hbb91b915;
    11'b00100111011: data <= 32'h3a5a3593;
    11'b00100111100: data <= 32'h3e383bb2;
    11'b00100111101: data <= 32'h3ddc26a9;
    11'b00100111110: data <= 32'h3de8bc19;
    11'b00100111111: data <= 32'h3d99b57e;
    11'b00101000000: data <= 32'h37c93d27;
    11'b00101000001: data <= 32'hb9a93da0;
    11'b00101000010: data <= 32'hba6db82c;
    11'b00101000011: data <= 32'h2f73c0a7;
    11'b00101000100: data <= 32'h369ec07c;
    11'b00101000101: data <= 32'hb7cabc40;
    11'b00101000110: data <= 32'hbc19b65d;
    11'b00101000111: data <= 32'ha55cb3d8;
    11'b00101001000: data <= 32'h3c80354a;
    11'b00101001001: data <= 32'h35483c70;
    11'b00101001010: data <= 32'hbf893c17;
    11'b00101001011: data <= 32'hc1b8323a;
    11'b00101001100: data <= 32'hbdebab24;
    11'b00101001101: data <= 32'h37393873;
    11'b00101001110: data <= 32'h3bf039b7;
    11'b00101001111: data <= 32'h38abb171;
    11'b00101010000: data <= 32'h3987b8f5;
    11'b00101010001: data <= 32'h3d08394e;
    11'b00101010010: data <= 32'h3c6f40b3;
    11'b00101010011: data <= 32'h32ea400a;
    11'b00101010100: data <= 32'hb29ab51b;
    11'b00101010101: data <= 32'h31e4c033;
    11'b00101010110: data <= 32'h359cbf01;
    11'b00101010111: data <= 32'haf46b8d9;
    11'b00101011000: data <= 32'hadc6b81f;
    11'b00101011001: data <= 32'h3c09bc77;
    11'b00101011010: data <= 32'h3eb3baf0;
    11'b00101011011: data <= 32'h34cc3400;
    11'b00101011100: data <= 32'hc02a3a53;
    11'b00101011101: data <= 32'hc1ae3448;
    11'b00101011110: data <= 32'hbd7db3f9;
    11'b00101011111: data <= 32'h3074b014;
    11'b00101100000: data <= 32'h9eacae62;
    11'b00101100001: data <= 32'hb9f8b84a;
    11'b00101100010: data <= 32'hb469b547;
    11'b00101100011: data <= 32'h3c223d0b;
    11'b00101100100: data <= 32'h3d6f418d;
    11'b00101100101: data <= 32'h356b4070;
    11'b00101100110: data <= 32'hb83d2c92;
    11'b00101100111: data <= 32'hb520bca8;
    11'b00101101000: data <= 32'h330db7dd;
    11'b00101101001: data <= 32'h366b34d7;
    11'b00101101010: data <= 32'h3a57b6eb;
    11'b00101101011: data <= 32'h3ef9bea8;
    11'b00101101100: data <= 32'h401ebd98;
    11'b00101101101: data <= 32'h39193193;
    11'b00101101110: data <= 32'hbd913bfd;
    11'b00101101111: data <= 32'hbf6e32dd;
    11'b00101110000: data <= 32'hb96abb1e;
    11'b00101110001: data <= 32'h2208bc8a;
    11'b00101110010: data <= 32'hbaf5bb98;
    11'b00101110011: data <= 32'hbec1bb7d;
    11'b00101110100: data <= 32'hb9c9b7be;
    11'b00101110101: data <= 32'h3c233b88;
    11'b00101110110: data <= 32'h3d10406b;
    11'b00101110111: data <= 32'hb4333f5e;
    11'b00101111000: data <= 32'hbdf636b0;
    11'b00101111001: data <= 32'hbc6dac70;
    11'b00101111010: data <= 32'ha83c3a03;
    11'b00101111011: data <= 32'h384d3c13;
    11'b00101111100: data <= 32'h3b26b592;
    11'b00101111101: data <= 32'h3e7bbed1;
    11'b00101111110: data <= 32'h4006bc22;
    11'b00101111111: data <= 32'h3c9b3b59;
    11'b00110000000: data <= 32'hb2b33e68;
    11'b00110000001: data <= 32'hb81433a9;
    11'b00110000010: data <= 32'h3058bd6f;
    11'b00110000011: data <= 32'h2a5cbe90;
    11'b00110000100: data <= 32'hbcb3bcca;
    11'b00110000101: data <= 32'hbedfbc79;
    11'b00110000110: data <= 32'hb548bc30;
    11'b00110000111: data <= 32'h3d98b144;
    11'b00110001000: data <= 32'h3c573bb8;
    11'b00110001001: data <= 32'hbc013c83;
    11'b00110001010: data <= 32'hc0a03867;
    11'b00110001011: data <= 32'hbe683888;
    11'b00110001100: data <= 32'hb4893cec;
    11'b00110001101: data <= 32'h2e2c3c20;
    11'b00110001110: data <= 32'h26f7b7a6;
    11'b00110001111: data <= 32'h391ebdae;
    11'b00110010000: data <= 32'h3e2ab20d;
    11'b00110010001: data <= 32'h3e283f96;
    11'b00110010010: data <= 32'h3a094064;
    11'b00110010011: data <= 32'h35d83670;
    11'b00110010100: data <= 32'h37eebcd3;
    11'b00110010101: data <= 32'h2d4cbca0;
    11'b00110010110: data <= 32'hbb63b895;
    11'b00110010111: data <= 32'hbbc9bb7c;
    11'b00110011000: data <= 32'h38c0bec0;
    11'b00110011001: data <= 32'h3fc6bd8f;
    11'b00110011010: data <= 32'h3c3fb19f;
    11'b00110011011: data <= 32'hbce93897;
    11'b00110011100: data <= 32'hc09537e6;
    11'b00110011101: data <= 32'hbd6d37d1;
    11'b00110011110: data <= 32'hb55a3a19;
    11'b00110011111: data <= 32'hb97d359c;
    11'b00110100000: data <= 32'hbd4ababe;
    11'b00110100001: data <= 32'hb8d5bcb4;
    11'b00110100010: data <= 32'h3bcb365b;
    11'b00110100011: data <= 32'h3e8140a0;
    11'b00110100100: data <= 32'h3bda4095;
    11'b00110100101: data <= 32'h347e38a0;
    11'b00110100110: data <= 32'h3118b75e;
    11'b00110100111: data <= 32'ha9022fac;
    11'b00110101000: data <= 32'hb7c038d5;
    11'b00110101001: data <= 32'hb07db7fd;
    11'b00110101010: data <= 32'h3d3fc017;
    11'b00110101011: data <= 32'h4084c006;
    11'b00110101100: data <= 32'h3cf0b819;
    11'b00110101101: data <= 32'hb9963898;
    11'b00110101110: data <= 32'hbd2e369b;
    11'b00110101111: data <= 32'hb68bab23;
    11'b00110110000: data <= 32'haf18b112;
    11'b00110110001: data <= 32'hbd61b78d;
    11'b00110110010: data <= 32'hc0b2bcd3;
    11'b00110110011: data <= 32'hbd53bcdf;
    11'b00110110100: data <= 32'h39d13292;
    11'b00110110101: data <= 32'h3dea3ef2;
    11'b00110110110: data <= 32'h37cb3ebe;
    11'b00110110111: data <= 32'hb87538b3;
    11'b00110111000: data <= 32'hb8a836ce;
    11'b00110111001: data <= 32'hb47e3dc2;
    11'b00110111010: data <= 32'hb4963e76;
    11'b00110111011: data <= 32'h2b10b02b;
    11'b00110111100: data <= 32'h3cbfc000;
    11'b00110111101: data <= 32'h4008bf09;
    11'b00110111110: data <= 32'h3dc12ce4;
    11'b00110111111: data <= 32'h34733c6c;
    11'b00111000000: data <= 32'h2ff83705;
    11'b00111000001: data <= 32'h39b0b855;
    11'b00111000010: data <= 32'h33ceb9ca;
    11'b00111000011: data <= 32'hbe25b9cd;
    11'b00111000100: data <= 32'hc0fabcf0;
    11'b00111000101: data <= 32'hbc81be08;
    11'b00111000110: data <= 32'h3be4b9a3;
    11'b00111000111: data <= 32'h3d3236db;
    11'b00111001000: data <= 32'hb3783949;
    11'b00111001001: data <= 32'hbd9f3612;
    11'b00111001010: data <= 32'hbc563b60;
    11'b00111001011: data <= 32'hb6b54011;
    11'b00111001100: data <= 32'hb8013f67;
    11'b00111001101: data <= 32'hb90daf71;
    11'b00111001110: data <= 32'h30e9bed4;
    11'b00111001111: data <= 32'h3cf9bbab;
    11'b00111010000: data <= 32'h3de33c2f;
    11'b00111010001: data <= 32'h3c553ed3;
    11'b00111010010: data <= 32'h3c793838;
    11'b00111010011: data <= 32'h3d50b88c;
    11'b00111010100: data <= 32'h376db65b;
    11'b00111010101: data <= 32'hbd0aabce;
    11'b00111010110: data <= 32'hbf3dba2c;
    11'b00111010111: data <= 32'hb3d0bf2f;
    11'b00111011000: data <= 32'h3e1dbf07;
    11'b00111011001: data <= 32'h3cecbaa7;
    11'b00111011010: data <= 32'hb8c1b1e3;
    11'b00111011011: data <= 32'hbe132dbf;
    11'b00111011100: data <= 32'hba873a63;
    11'b00111011101: data <= 32'hb31a3e99;
    11'b00111011110: data <= 32'hbb963cff;
    11'b00111011111: data <= 32'hbf37b766;
    11'b00111100000: data <= 32'hbcd4bdc3;
    11'b00111100001: data <= 32'h35c6b476;
    11'b00111100010: data <= 32'h3d233e4e;
    11'b00111100011: data <= 32'h3cf63f2b;
    11'b00111100100: data <= 32'h3c8b37e1;
    11'b00111100101: data <= 32'h3c74b02c;
    11'b00111100110: data <= 32'h363539a0;
    11'b00111100111: data <= 32'hba7e3ce8;
    11'b00111101000: data <= 32'hbb5b9f8d;
    11'b00111101001: data <= 32'h3888bf63;
    11'b00111101010: data <= 32'h3f68c093;
    11'b00111101011: data <= 32'h3cefbd25;
    11'b00111101100: data <= 32'hb56fb5a2;
    11'b00111101101: data <= 32'hb989acc1;
    11'b00111101110: data <= 32'h337733ea;
    11'b00111101111: data <= 32'h354939a6;
    11'b00111110000: data <= 32'hbd1e35be;
    11'b00111110001: data <= 32'hc16fbac3;
    11'b00111110010: data <= 32'hc021bd69;
    11'b00111110011: data <= 32'hae71b360;
    11'b00111110100: data <= 32'h3c083ca8;
    11'b00111110101: data <= 32'h39db3c67;
    11'b00111110110: data <= 32'h34e631e4;
    11'b00111110111: data <= 32'h356636b6;
    11'b00111111000: data <= 32'h2fd93f99;
    11'b00111111001: data <= 32'hb82d40c3;
    11'b00111111010: data <= 32'hb82938f3;
    11'b00111111011: data <= 32'h38ccbe81;
    11'b00111111100: data <= 32'h3e2dc003;
    11'b00111111101: data <= 32'h3c90b9e0;
    11'b00111111110: data <= 32'h34d9319e;
    11'b00111111111: data <= 32'h38c7a853;
    11'b01000000000: data <= 32'h3e05b4cf;
    11'b01000000001: data <= 32'h3bd2a6b5;
    11'b01000000010: data <= 32'hbd03a9e8;
    11'b01000000011: data <= 32'hc1a3bab1;
    11'b01000000100: data <= 32'hbfb3bd84;
    11'b01000000101: data <= 32'h2f08ba8a;
    11'b01000000110: data <= 32'h3a93a01b;
    11'b01000000111: data <= 32'ha7dcad11;
    11'b01000001000: data <= 32'hb962b583;
    11'b01000001001: data <= 32'hb4e2394f;
    11'b01000001010: data <= 32'h9d6440e2;
    11'b01000001011: data <= 32'hb815416b;
    11'b01000001100: data <= 32'hbb3839d7;
    11'b01000001101: data <= 32'hb4a6bd2f;
    11'b01000001110: data <= 32'h38fdbcb2;
    11'b01000001111: data <= 32'h3ab53557;
    11'b01000010000: data <= 32'h3a9c3b31;
    11'b01000010001: data <= 32'h3e1d2c23;
    11'b01000010010: data <= 32'h407db819;
    11'b01000010011: data <= 32'h3d6424e5;
    11'b01000010100: data <= 32'hbb3a377d;
    11'b01000010101: data <= 32'hc038b3c2;
    11'b01000010110: data <= 32'hbbd0bd51;
    11'b01000010111: data <= 32'h3a02be46;
    11'b01000011000: data <= 32'h3a33bcca;
    11'b01000011001: data <= 32'hb854bc4b;
    11'b01000011010: data <= 32'hbc2abab2;
    11'b01000011011: data <= 32'hb22d36d1;
    11'b01000011100: data <= 32'h34c5400f;
    11'b01000011101: data <= 32'hb9124026;
    11'b01000011110: data <= 32'hbf0d350d;
    11'b01000011111: data <= 32'hbe49bc35;
    11'b01000100000: data <= 32'hb6deb5fb;
    11'b01000100001: data <= 32'h36633c60;
    11'b01000100010: data <= 32'h3aa13c95;
    11'b01000100011: data <= 32'h3e15aa1d;
    11'b01000100100: data <= 32'h4013b5ff;
    11'b01000100101: data <= 32'h3cfa3a78;
    11'b01000100110: data <= 32'hb7823ea9;
    11'b01000100111: data <= 32'hbc7e399e;
    11'b01000101000: data <= 32'h28f2bc5c;
    11'b01000101001: data <= 32'h3cf3bfa0;
    11'b01000101010: data <= 32'h39d5be80;
    11'b01000101011: data <= 32'hb877bd2b;
    11'b01000101100: data <= 32'hb828bc18;
    11'b01000101101: data <= 32'h3a0cb024;
    11'b01000101110: data <= 32'h3c1f3c09;
    11'b01000101111: data <= 32'hb9333c08;
    11'b01000110000: data <= 32'hc0e7b34d;
    11'b01000110001: data <= 32'hc0cdbb8b;
    11'b01000110010: data <= 32'hbbddad5b;
    11'b01000110011: data <= 32'h29673bd3;
    11'b01000110100: data <= 32'h349b388a;
    11'b01000110101: data <= 32'h3908b836;
    11'b01000110110: data <= 32'h3c78b0d8;
    11'b01000110111: data <= 32'h3aa23f08;
    11'b01000111000: data <= 32'hb1ba4194;
    11'b01000111001: data <= 32'hb8183dd4;
    11'b01000111010: data <= 32'h35c4b9da;
    11'b01000111011: data <= 32'h3c3ebe3b;
    11'b01000111100: data <= 32'h37c1bc18;
    11'b01000111101: data <= 32'hb3c6b947;
    11'b01000111110: data <= 32'h380fbadd;
    11'b01000111111: data <= 32'h3ffbb953;
    11'b01001000000: data <= 32'h3f5b2e08;
    11'b01001000001: data <= 32'hb6f33533;
    11'b01001000010: data <= 32'hc0e6b5e7;
    11'b01001000011: data <= 32'hc071bac0;
    11'b01001000100: data <= 32'hb9b2b59d;
    11'b01001000101: data <= 32'hab0e2d1a;
    11'b01001000110: data <= 32'hb769b898;
    11'b01001000111: data <= 32'hb80ebcf5;
    11'b01001001000: data <= 32'h32c8b085;
    11'b01001001001: data <= 32'h38484055;
    11'b01001001010: data <= 32'hacc3422e;
    11'b01001001011: data <= 32'hb8b73e39;
    11'b01001001100: data <= 32'hb3e0b71d;
    11'b01001001101: data <= 32'h3211b9cd;
    11'b01001001110: data <= 32'ha39331ba;
    11'b01001001111: data <= 32'h21ba34e2;
    11'b01001010000: data <= 32'h3d1eb8ae;
    11'b01001010001: data <= 32'h4171bb84;
    11'b01001010010: data <= 32'h407db09c;
    11'b01001010011: data <= 32'hacda3861;
    11'b01001010100: data <= 32'hbee730fc;
    11'b01001010101: data <= 32'hbca1b8c8;
    11'b01001010110: data <= 32'h309cba76;
    11'b01001010111: data <= 32'h2c78bb6a;
    11'b01001011000: data <= 32'hbc0cbe44;
    11'b01001011001: data <= 32'hbc8cbf45;
    11'b01001011010: data <= 32'h2713b70f;
    11'b01001011011: data <= 32'h39f43ee0;
    11'b01001011100: data <= 32'ha3c640b9;
    11'b01001011101: data <= 32'hbc913baf;
    11'b01001011110: data <= 32'hbd4ab5be;
    11'b01001011111: data <= 32'hbaf12e41;
    11'b01001100000: data <= 32'hb8ae3cb8;
    11'b01001100001: data <= 32'hae9b3acd;
    11'b01001100010: data <= 32'h3cd9b89f;
    11'b01001100011: data <= 32'h40e2bbb3;
    11'b01001100100: data <= 32'h40013555;
    11'b01001100101: data <= 32'h332e3e16;
    11'b01001100110: data <= 32'hb9c83c69;
    11'b01001100111: data <= 32'h2d20b225;
    11'b01001101000: data <= 32'h3b6bbbd3;
    11'b01001101001: data <= 32'h3153bd18;
    11'b01001101010: data <= 32'hbca7bef6;
    11'b01001101011: data <= 32'hbb64bfac;
    11'b01001101100: data <= 32'h39e1bb2e;
    11'b01001101101: data <= 32'h3de13975;
    11'b01001101110: data <= 32'h31063c5d;
    11'b01001101111: data <= 32'hbe7d3003;
    11'b01001110000: data <= 32'hc019b690;
    11'b01001110001: data <= 32'hbd9c37f9;
    11'b01001110010: data <= 32'hbb4e3d78;
    11'b01001110011: data <= 32'hb8b83840;
    11'b01001110100: data <= 32'h34d5bc21;
    11'b01001110101: data <= 32'h3d5ebb7c;
    11'b01001110110: data <= 32'h3d3f3c2c;
    11'b01001110111: data <= 32'h357b410b;
    11'b01001111000: data <= 32'ha5fb3f71;
    11'b01001111001: data <= 32'h39983237;
    11'b01001111010: data <= 32'h3c1db910;
    11'b01001111011: data <= 32'ha7cfb928;
    11'b01001111100: data <= 32'hbc2cbba7;
    11'b01001111101: data <= 32'hb110be05;
    11'b01001111110: data <= 32'h3f55bd0c;
    11'b01001111111: data <= 32'h4097b4d5;
    11'b01010000000: data <= 32'h37372f82;
    11'b01010000001: data <= 32'hbe4bb4fe;
    11'b01010000010: data <= 32'hbf52b631;
    11'b01010000011: data <= 32'hbc0b36aa;
    11'b01010000100: data <= 32'hba6e39fb;
    11'b01010000101: data <= 32'hbcbcb735;
    11'b01010000110: data <= 32'hbb1ebf17;
    11'b01010000111: data <= 32'h3107bc2f;
    11'b01010001000: data <= 32'h39a73d70;
    11'b01010001001: data <= 32'h3574418b;
    11'b01010001010: data <= 32'h2c703f7d;
    11'b01010001011: data <= 32'h362a352f;
    11'b01010001100: data <= 32'h35742c66;
    11'b01010001101: data <= 32'hb87538da;
    11'b01010001110: data <= 32'hbb8a3459;
    11'b01010001111: data <= 32'h37b5bb51;
    11'b01010010000: data <= 32'h40ffbd9c;
    11'b01010010001: data <= 32'h414db988;
    11'b01010010010: data <= 32'h39a728a5;
    11'b01010010011: data <= 32'hbb8d1393;
    11'b01010010100: data <= 32'hb9c3affc;
    11'b01010010101: data <= 32'h2d9b3059;
    11'b01010010110: data <= 32'hb5e3ade1;
    11'b01010010111: data <= 32'hbe53bd7f;
    11'b01010011000: data <= 32'hbe9cc0aa;
    11'b01010011001: data <= 32'hb569bd32;
    11'b01010011010: data <= 32'h39623bbf;
    11'b01010011011: data <= 32'h364f3ffe;
    11'b01010011100: data <= 32'hb4b93c3e;
    11'b01010011101: data <= 32'hb7e02f7e;
    11'b01010011110: data <= 32'hb91539e1;
    11'b01010011111: data <= 32'hbc903ee6;
    11'b01010100000: data <= 32'hbc433c87;
    11'b01010100001: data <= 32'h36edb915;
    11'b01010100010: data <= 32'h405bbd90;
    11'b01010100011: data <= 32'h4072b671;
    11'b01010100100: data <= 32'h39f23a44;
    11'b01010100101: data <= 32'hadfe3ac9;
    11'b01010100110: data <= 32'h39003508;
    11'b01010100111: data <= 32'h3cc02665;
    11'b01010101000: data <= 32'h2680b6b0;
    11'b01010101001: data <= 32'hbeadbe0a;
    11'b01010101010: data <= 32'hbe7dc095;
    11'b01010101011: data <= 32'h2f8cbe21;
    11'b01010101100: data <= 32'h3d172c98;
    11'b01010101101: data <= 32'h38db3906;
    11'b01010101110: data <= 32'hb967ada9;
    11'b01010101111: data <= 32'hbca4b3f6;
    11'b01010110000: data <= 32'hbc8b3c2e;
    11'b01010110001: data <= 32'hbd7b402e;
    11'b01010110010: data <= 32'hbd833c58;
    11'b01010110011: data <= 32'hb5b7bb78;
    11'b01010110100: data <= 32'h3be8bd9a;
    11'b01010110101: data <= 32'h3cec31a8;
    11'b01010110110: data <= 32'h384f3ec3;
    11'b01010110111: data <= 32'h37ef3e49;
    11'b01010111000: data <= 32'h3da9392b;
    11'b01010111001: data <= 32'h3e573407;
    11'b01010111010: data <= 32'h249e2f75;
    11'b01010111011: data <= 32'hbe48b932;
    11'b01010111100: data <= 32'hbc07be64;
    11'b01010111101: data <= 32'h3c5dbe4f;
    11'b01010111110: data <= 32'h401eba4f;
    11'b01010111111: data <= 32'h3b12b817;
    11'b01011000000: data <= 32'hb985bac1;
    11'b01011000001: data <= 32'hbc06b739;
    11'b01011000010: data <= 32'hb9743bbc;
    11'b01011000011: data <= 32'hbc103e89;
    11'b01011000100: data <= 32'hbeaf342b;
    11'b01011000101: data <= 32'hbdadbe7e;
    11'b01011000110: data <= 32'hb5b1be16;
    11'b01011000111: data <= 32'h34a1380f;
    11'b01011001000: data <= 32'h34643fe7;
    11'b01011001001: data <= 32'h388c3e23;
    11'b01011001010: data <= 32'h3d1c3895;
    11'b01011001011: data <= 32'h3c57397a;
    11'b01011001100: data <= 32'hb70b3cf6;
    11'b01011001101: data <= 32'hbdff39d4;
    11'b01011001110: data <= 32'hb64eb94e;
    11'b01011001111: data <= 32'h3f0fbdb3;
    11'b01011010000: data <= 32'h40c1bc89;
    11'b01011010001: data <= 32'h3bdaba37;
    11'b01011010010: data <= 32'hb49bba0c;
    11'b01011010011: data <= 32'ha27ab493;
    11'b01011010100: data <= 32'h387239cb;
    11'b01011010101: data <= 32'hb3a33add;
    11'b01011010110: data <= 32'hbf07b929;
    11'b01011010111: data <= 32'hc03bc053;
    11'b01011011000: data <= 32'hbc2bbea6;
    11'b01011011001: data <= 32'h9ec734ca;
    11'b01011011010: data <= 32'h32383d37;
    11'b01011011011: data <= 32'h33ab38c7;
    11'b01011011100: data <= 32'h37e9290d;
    11'b01011011101: data <= 32'h30fe3c23;
    11'b01011011110: data <= 32'hbc0a408e;
    11'b01011011111: data <= 32'hbe373f23;
    11'b01011100000: data <= 32'hb4e2ad8b;
    11'b01011100001: data <= 32'h3e21bcf4;
    11'b01011100010: data <= 32'h3f63baf3;
    11'b01011100011: data <= 32'h39bdb0dd;
    11'b01011100100: data <= 32'h340d216d;
    11'b01011100101: data <= 32'h3cfa306f;
    11'b01011100110: data <= 32'h3f6a38ab;
    11'b01011100111: data <= 32'h37af3704;
    11'b01011101000: data <= 32'hbe85bad9;
    11'b01011101001: data <= 32'hc02fc013;
    11'b01011101010: data <= 32'hb9d8be85;
    11'b01011101011: data <= 32'h3793b4e4;
    11'b01011101100: data <= 32'h36132652;
    11'b01011101101: data <= 32'hb089b9fe;
    11'b01011101110: data <= 32'hb32bb962;
    11'b01011101111: data <= 32'hb6793c63;
    11'b01011110000: data <= 32'hbcbd4144;
    11'b01011110001: data <= 32'hbe943f9d;
    11'b01011110010: data <= 32'hbaa3b329;
    11'b01011110011: data <= 32'h36f1bcc8;
    11'b01011110100: data <= 32'h394ab4e0;
    11'b01011110101: data <= 32'h30ed3a21;
    11'b01011110110: data <= 32'h388d3a34;
    11'b01011110111: data <= 32'h4007370d;
    11'b01011111000: data <= 32'h40df3917;
    11'b01011111001: data <= 32'h396c39eb;
    11'b01011111010: data <= 32'hbdcbad9a;
    11'b01011111011: data <= 32'hbdffbcab;
    11'b01011111100: data <= 32'h3301bd45;
    11'b01011111101: data <= 32'h3d1cbb01;
    11'b01011111110: data <= 32'h3925bc56;
    11'b01011111111: data <= 32'hb489bed8;
    11'b01100000000: data <= 32'hb444bc80;
    11'b01100000001: data <= 32'ha96d3b2f;
    11'b01100000010: data <= 32'hb96a4066;
    11'b01100000011: data <= 32'hbe623c87;
    11'b01100000100: data <= 32'hbe61bb39;
    11'b01100000101: data <= 32'hbaf8bd3e;
    11'b01100000110: data <= 32'hb8072f44;
    11'b01100000111: data <= 32'hb6703cd8;
    11'b01100001000: data <= 32'h37bd3a9f;
    11'b01100001001: data <= 32'h3f9533ce;
    11'b01100001010: data <= 32'h400c3a0e;
    11'b01100001011: data <= 32'h343c3e4a;
    11'b01100001100: data <= 32'hbd793cf9;
    11'b01100001101: data <= 32'hbaa48d0c;
    11'b01100001110: data <= 32'h3c12bab2;
    11'b01100001111: data <= 32'h3ebcbc1b;
    11'b01100010000: data <= 32'h3931bd78;
    11'b01100010001: data <= 32'hb0ffbefc;
    11'b01100010010: data <= 32'h3735bc30;
    11'b01100010011: data <= 32'h3c903913;
    11'b01100010100: data <= 32'h354e3d91;
    11'b01100010101: data <= 32'hbd52304d;
    11'b01100010110: data <= 32'hc021be17;
    11'b01100010111: data <= 32'hbe48bd8f;
    11'b01100011000: data <= 32'hbbae3076;
    11'b01100011001: data <= 32'hb8f63a5e;
    11'b01100011010: data <= 32'h2f24aa2f;
    11'b01100011011: data <= 32'h3c66b814;
    11'b01100011100: data <= 32'h3c2539f8;
    11'b01100011101: data <= 32'hb60140b9;
    11'b01100011110: data <= 32'hbd8c409d;
    11'b01100011111: data <= 32'hb8603a29;
    11'b01100100000: data <= 32'h3c15b758;
    11'b01100100001: data <= 32'h3ce2b980;
    11'b01100100010: data <= 32'h31ddb9f2;
    11'b01100100011: data <= 32'h278dbbac;
    11'b01100100100: data <= 32'h3dcab892;
    11'b01100100101: data <= 32'h40e337a0;
    11'b01100100110: data <= 32'h3d163a89;
    11'b01100100111: data <= 32'hbbb2b4a8;
    11'b01100101000: data <= 32'hbfbcbdea;
    11'b01100101001: data <= 32'hbd14bcba;
    11'b01100101010: data <= 32'hb801b003;
    11'b01100101011: data <= 32'hb6a3b30a;
    11'b01100101100: data <= 32'hb473bd96;
    11'b01100101101: data <= 32'h342abddc;
    11'b01100101110: data <= 32'h348b3833;
    11'b01100101111: data <= 32'hb9254126;
    11'b01100110000: data <= 32'hbd5840e4;
    11'b01100110001: data <= 32'hba0a3994;
    11'b01100110010: data <= 32'h31efb64f;
    11'b01100110011: data <= 32'h2902af16;
    11'b01100110100: data <= 32'hb9133442;
    11'b01100110101: data <= 32'h277fa789;
    11'b01100110110: data <= 32'h4018b167;
    11'b01100110111: data <= 32'h421b36cb;
    11'b01100111000: data <= 32'h3e503aa7;
    11'b01100111001: data <= 32'hb9ad32f7;
    11'b01100111010: data <= 32'hbd40b8fe;
    11'b01100111011: data <= 32'hb410b8eb;
    11'b01100111100: data <= 32'h3701b5b9;
    11'b01100111101: data <= 32'haa90bc8e;
    11'b01100111110: data <= 32'hb7e1c0ca;
    11'b01100111111: data <= 32'ha877c024;
    11'b01101000000: data <= 32'h3646328d;
    11'b01101000001: data <= 32'hb16e4030;
    11'b01101000010: data <= 32'hbc2e3e83;
    11'b01101000011: data <= 32'hbcafad27;
    11'b01101000100: data <= 32'hbb4db8c8;
    11'b01101000101: data <= 32'hbcad35b3;
    11'b01101000110: data <= 32'hbd8c3b70;
    11'b01101000111: data <= 32'hb353344c;
    11'b01101001000: data <= 32'h3f70b4f5;
    11'b01101001001: data <= 32'h413b353c;
    11'b01101001010: data <= 32'h3c6d3d45;
    11'b01101001011: data <= 32'hb9913d50;
    11'b01101001100: data <= 32'hb8de38b6;
    11'b01101001101: data <= 32'h39df2e40;
    11'b01101001110: data <= 32'h3c4fb495;
    11'b01101001111: data <= 32'h27cabd51;
    11'b01101010000: data <= 32'hb869c0db;
    11'b01101010001: data <= 32'h3593bfed;
    11'b01101010010: data <= 32'h3d61a629;
    11'b01101010011: data <= 32'h3b093d06;
    11'b01101010100: data <= 32'hb82f377b;
    11'b01101010101: data <= 32'hbd83bb5b;
    11'b01101010110: data <= 32'hbdfdba27;
    11'b01101010111: data <= 32'hbe96384a;
    11'b01101011000: data <= 32'hbe973aa3;
    11'b01101011001: data <= 32'hb8dbb5ec;
    11'b01101011010: data <= 32'h3c21bc5e;
    11'b01101011011: data <= 32'h3df72a92;
    11'b01101011100: data <= 32'h34423f3f;
    11'b01101011101: data <= 32'hba8a4084;
    11'b01101011110: data <= 32'hb26d3d9c;
    11'b01101011111: data <= 32'h3c213898;
    11'b01101100000: data <= 32'h3adc2ee2;
    11'b01101100001: data <= 32'hb71eb955;
    11'b01101100010: data <= 32'hb903be21;
    11'b01101100011: data <= 32'h3c21bd54;
    11'b01101100100: data <= 32'h40feace1;
    11'b01101100101: data <= 32'h3f8538a8;
    11'b01101100110: data <= 32'h9c71b37a;
    11'b01101100111: data <= 32'hbc8ebc81;
    11'b01101101000: data <= 32'hbc96b89a;
    11'b01101101001: data <= 32'hbc723826;
    11'b01101101010: data <= 32'hbd3b3058;
    11'b01101101011: data <= 32'hbb35be37;
    11'b01101101100: data <= 32'h2f64c03c;
    11'b01101101101: data <= 32'h37bdb5d3;
    11'b01101101110: data <= 32'hb41f3f7b;
    11'b01101101111: data <= 32'hba7640a9;
    11'b01101110000: data <= 32'hb1ce3d25;
    11'b01101110001: data <= 32'h382c386e;
    11'b01101110010: data <= 32'hb0a738e4;
    11'b01101110011: data <= 32'hbd59367f;
    11'b01101110100: data <= 32'hbad6b5ef;
    11'b01101110101: data <= 32'h3dbeb962;
    11'b01101110110: data <= 32'h420fabd2;
    11'b01101110111: data <= 32'h405a3651;
    11'b01101111000: data <= 32'h32fbaa43;
    11'b01101111001: data <= 32'hb873b775;
    11'b01101111010: data <= 32'hacb92bea;
    11'b01101111011: data <= 32'h281a384b;
    11'b01101111100: data <= 32'hb992b86c;
    11'b01101111101: data <= 32'hbc1bc0ee;
    11'b01101111110: data <= 32'hb5aac17e;
    11'b01101111111: data <= 32'h3459b9b1;
    11'b01110000000: data <= 32'h14683d8b;
    11'b01110000001: data <= 32'hb7663dd5;
    11'b01110000010: data <= 32'hb5653553;
    11'b01110000011: data <= 32'hb51c2fe0;
    11'b01110000100: data <= 32'hbd093bd7;
    11'b01110000101: data <= 32'hc0493ce0;
    11'b01110000110: data <= 32'hbcc833aa;
    11'b01110000111: data <= 32'h3ccfb8a1;
    11'b01110001000: data <= 32'h4112b1fc;
    11'b01110001001: data <= 32'h3e3f38f8;
    11'b01110001010: data <= 32'h288f3a44;
    11'b01110001011: data <= 32'h2a8d391f;
    11'b01110001100: data <= 32'h3c2d3ad4;
    11'b01110001101: data <= 32'h3bc939f3;
    11'b01110001110: data <= 32'hb5cbb943;
    11'b01110001111: data <= 32'hbc57c0e3;
    11'b01110010000: data <= 32'hb306c11b;
    11'b01110010001: data <= 32'h3b70ba47;
    11'b01110010010: data <= 32'h3b69390e;
    11'b01110010011: data <= 32'h30e131d4;
    11'b01110010100: data <= 32'hb5ceba5d;
    11'b01110010101: data <= 32'hba3db4fe;
    11'b01110010110: data <= 32'hbebe3c86;
    11'b01110010111: data <= 32'hc0b03d67;
    11'b01110011000: data <= 32'hbde0adf4;
    11'b01110011001: data <= 32'h3705bcdc;
    11'b01110011010: data <= 32'h3d3bb874;
    11'b01110011011: data <= 32'h372d3b37;
    11'b01110011100: data <= 32'hb5a93e35;
    11'b01110011101: data <= 32'h36813d9d;
    11'b01110011110: data <= 32'h3e3b3d43;
    11'b01110011111: data <= 32'h3c463c5b;
    11'b01110100000: data <= 32'hb956a808;
    11'b01110100001: data <= 32'hbcf9bdd4;
    11'b01110100010: data <= 32'h3365be9f;
    11'b01110100011: data <= 32'h3f8fb899;
    11'b01110100100: data <= 32'h3f7e26c0;
    11'b01110100101: data <= 32'h3998b9c2;
    11'b01110100110: data <= 32'haf44bd4d;
    11'b01110100111: data <= 32'hb6ecb50c;
    11'b01110101000: data <= 32'hbc493cb6;
    11'b01110101001: data <= 32'hbf2a3b33;
    11'b01110101010: data <= 32'hbe13bc3d;
    11'b01110101011: data <= 32'hb66cc05c;
    11'b01110101100: data <= 32'h2f37bc22;
    11'b01110101101: data <= 32'hb67e3b26;
    11'b01110101110: data <= 32'hb88c3e61;
    11'b01110101111: data <= 32'h377c3ce3;
    11'b01110110000: data <= 32'h3d2c3c80;
    11'b01110110001: data <= 32'h34e23d88;
    11'b01110110010: data <= 32'hbdf33bb9;
    11'b01110110011: data <= 32'hbe38afda;
    11'b01110110100: data <= 32'h382bb94f;
    11'b01110110101: data <= 32'h40b8b4f5;
    11'b01110110110: data <= 32'h403cb1aa;
    11'b01110110111: data <= 32'h3a67ba40;
    11'b01110111000: data <= 32'h34dbbb6e;
    11'b01110111001: data <= 32'h3898336a;
    11'b01110111010: data <= 32'h33583d2b;
    11'b01110111011: data <= 32'hbad835cc;
    11'b01110111100: data <= 32'hbd82bf86;
    11'b01110111101: data <= 32'hbae5c189;
    11'b01110111110: data <= 32'hb57dbd3c;
    11'b01110111111: data <= 32'hb6f93831;
    11'b01111000000: data <= 32'hb5703a2a;
    11'b01111000001: data <= 32'h36923014;
    11'b01111000010: data <= 32'h3911363b;
    11'b01111000011: data <= 32'hb9893dea;
    11'b01111000100: data <= 32'hc0873eff;
    11'b01111000101: data <= 32'hbf7d39cf;
    11'b01111000110: data <= 32'h359db418;
    11'b01111000111: data <= 32'h3f94b491;
    11'b01111001000: data <= 32'h3d85a932;
    11'b01111001001: data <= 32'h3578b0f3;
    11'b01111001010: data <= 32'h39312858;
    11'b01111001011: data <= 32'h3e9b3bfd;
    11'b01111001100: data <= 32'h3d9c3e13;
    11'b01111001101: data <= 32'hb1ff33d7;
    11'b01111001110: data <= 32'hbcffbf79;
    11'b01111001111: data <= 32'hba67c0f2;
    11'b01111010000: data <= 32'h2de3bc93;
    11'b01111010001: data <= 32'h35092152;
    11'b01111010010: data <= 32'h33dfb763;
    11'b01111010011: data <= 32'h3709bce6;
    11'b01111010100: data <= 32'h32a8b647;
    11'b01111010101: data <= 32'hbc6f3da6;
    11'b01111010110: data <= 32'hc0c73fbb;
    11'b01111010111: data <= 32'hbfd03908;
    11'b01111011000: data <= 32'hb285b979;
    11'b01111011001: data <= 32'h39aab8e2;
    11'b01111011010: data <= 32'h2a983129;
    11'b01111011011: data <= 32'hb6633849;
    11'b01111011100: data <= 32'h3a1d3a24;
    11'b01111011101: data <= 32'h40653da5;
    11'b01111011110: data <= 32'h3ef93ee6;
    11'b01111011111: data <= 32'hb4013999;
    11'b01111100000: data <= 32'hbd59bb59;
    11'b01111100001: data <= 32'hb705bd81;
    11'b01111100010: data <= 32'h3b7eb8b4;
    11'b01111100011: data <= 32'h3cd7b575;
    11'b01111100100: data <= 32'h3a20bd87;
    11'b01111100101: data <= 32'h38d4c004;
    11'b01111100110: data <= 32'h36d5b95f;
    11'b01111100111: data <= 32'hb8383d6f;
    11'b01111101000: data <= 32'hbea13e49;
    11'b01111101001: data <= 32'hbeb3b227;
    11'b01111101010: data <= 32'hba4abe4a;
    11'b01111101011: data <= 32'hb7ecbc4b;
    11'b01111101100: data <= 32'hbc433213;
    11'b01111101101: data <= 32'hbb61394b;
    11'b01111101110: data <= 32'h398538e9;
    11'b01111101111: data <= 32'h40093c4b;
    11'b01111110000: data <= 32'h3c9b3ee2;
    11'b01111110001: data <= 32'hbbb93dc9;
    11'b01111110010: data <= 32'hbe8e36a8;
    11'b01111110011: data <= 32'hb0deaf70;
    11'b01111110100: data <= 32'h3dc823bc;
    11'b01111110101: data <= 32'h3de5b605;
    11'b01111110110: data <= 32'h3a06be16;
    11'b01111110111: data <= 32'h3a23bf3e;
    11'b01111111000: data <= 32'h3ccfb435;
    11'b01111111001: data <= 32'h3a243dd3;
    11'b01111111010: data <= 32'hb7513c44;
    11'b01111111011: data <= 32'hbcb3bc0e;
    11'b01111111100: data <= 32'hbc31c057;
    11'b01111111101: data <= 32'hbc15bd12;
    11'b01111111110: data <= 32'hbd492643;
    11'b01111111111: data <= 32'hbafa292c;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    