
module memory_rom_35(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbe18b6e8;
    11'b00000000001: data <= 32'hbafab21b;
    11'b00000000010: data <= 32'h3b1d34a9;
    11'b00000000011: data <= 32'h3d7d3d1a;
    11'b00000000100: data <= 32'hb5443ec8;
    11'b00000000101: data <= 32'hc0403c0b;
    11'b00000000110: data <= 32'hbf423511;
    11'b00000000111: data <= 32'ha4f03866;
    11'b00000001000: data <= 32'h3c513a8a;
    11'b00000001001: data <= 32'h3b7ead19;
    11'b00000001010: data <= 32'h3ad7bd23;
    11'b00000001011: data <= 32'h3da6bad5;
    11'b00000001100: data <= 32'h3e543c55;
    11'b00000001101: data <= 32'h39da4011;
    11'b00000001110: data <= 32'hb1ae3890;
    11'b00000001111: data <= 32'hb3e8be6e;
    11'b00000010000: data <= 32'hb03cc03a;
    11'b00000010001: data <= 32'hb967bc6d;
    11'b00000010010: data <= 32'hbc67b84d;
    11'b00000010011: data <= 32'hb205bbcb;
    11'b00000010100: data <= 32'h3d1fbc23;
    11'b00000010101: data <= 32'h3c89297f;
    11'b00000010110: data <= 32'hbb9d3c8b;
    11'b00000010111: data <= 32'hc1393c8f;
    11'b00000011000: data <= 32'hbfee38f9;
    11'b00000011001: data <= 32'hb3943842;
    11'b00000011010: data <= 32'h357c37db;
    11'b00000011011: data <= 32'hb4b0b390;
    11'b00000011100: data <= 32'hb462baf3;
    11'b00000011101: data <= 32'h3c091da2;
    11'b00000011110: data <= 32'h3fea3f74;
    11'b00000011111: data <= 32'h3dad40cf;
    11'b00000100000: data <= 32'h333f3a13;
    11'b00000100001: data <= 32'hb343bc6c;
    11'b00000100010: data <= 32'hadd4bcb4;
    11'b00000100011: data <= 32'hb1cfb323;
    11'b00000100100: data <= 32'hb1cfb5d8;
    11'b00000100101: data <= 32'h3978beaf;
    11'b00000100110: data <= 32'h3ec4c034;
    11'b00000100111: data <= 32'h3cb3b9d2;
    11'b00000101000: data <= 32'hba7d3afd;
    11'b00000101001: data <= 32'hc0363c1f;
    11'b00000101010: data <= 32'hbdc4324b;
    11'b00000101011: data <= 32'hb4b9b44c;
    11'b00000101100: data <= 32'hb89db465;
    11'b00000101101: data <= 32'hbe8ab830;
    11'b00000101110: data <= 32'hbd31b961;
    11'b00000101111: data <= 32'h39313432;
    11'b00000110000: data <= 32'h3fe83f49;
    11'b00000110001: data <= 32'h3cf34071;
    11'b00000110010: data <= 32'hb4de3bed;
    11'b00000110011: data <= 32'hba0caf7d;
    11'b00000110100: data <= 32'hb0fd33f1;
    11'b00000110101: data <= 32'h34953b17;
    11'b00000110110: data <= 32'h36e1a9e6;
    11'b00000110111: data <= 32'h3c16bfb1;
    11'b00000111000: data <= 32'h3f1fc0a1;
    11'b00000111001: data <= 32'h3de3b8a4;
    11'b00000111010: data <= 32'h2cde3c7a;
    11'b00000111011: data <= 32'hba903b0f;
    11'b00000111100: data <= 32'hb709b7db;
    11'b00000111101: data <= 32'hb03bbc87;
    11'b00000111110: data <= 32'hbc94babe;
    11'b00000111111: data <= 32'hc09bb9c4;
    11'b00001000000: data <= 32'hbe50bb16;
    11'b00001000001: data <= 32'h3910b5f7;
    11'b00001000010: data <= 32'h3ee13abf;
    11'b00001000011: data <= 32'h37ae3df0;
    11'b00001000100: data <= 32'hbd0d3c3f;
    11'b00001000101: data <= 32'hbd8f3a00;
    11'b00001000110: data <= 32'hb4a23d3f;
    11'b00001000111: data <= 32'h34fd3e28;
    11'b00001001000: data <= 32'h313a30ee;
    11'b00001001001: data <= 32'h36febecf;
    11'b00001001010: data <= 32'h3d79bec3;
    11'b00001001011: data <= 32'h3f23346f;
    11'b00001001100: data <= 32'h3ca43eb1;
    11'b00001001101: data <= 32'h37d13ab9;
    11'b00001001110: data <= 32'h36e8bace;
    11'b00001001111: data <= 32'h2fe9bd2e;
    11'b00001010000: data <= 32'hbc69b93b;
    11'b00001010001: data <= 32'hbffcb8ac;
    11'b00001010010: data <= 32'hbc09bd67;
    11'b00001010011: data <= 32'h3be7be2b;
    11'b00001010100: data <= 32'h3de4b838;
    11'b00001010101: data <= 32'hb26a38be;
    11'b00001010110: data <= 32'hbf513b47;
    11'b00001010111: data <= 32'hbe253bfb;
    11'b00001011000: data <= 32'hb4e53db5;
    11'b00001011001: data <= 32'hb0693d79;
    11'b00001011010: data <= 32'hbb4e2bb9;
    11'b00001011011: data <= 32'hba93bd28;
    11'b00001011100: data <= 32'h38fdba7a;
    11'b00001011101: data <= 32'h3f7b3c75;
    11'b00001011110: data <= 32'h3f144012;
    11'b00001011111: data <= 32'h3c283af8;
    11'b00001100000: data <= 32'h3937b8ca;
    11'b00001100001: data <= 32'h3439b805;
    11'b00001100010: data <= 32'hb8ea358d;
    11'b00001100011: data <= 32'hbc5aaccc;
    11'b00001100100: data <= 32'haec8bee2;
    11'b00001100101: data <= 32'h3d9cc106;
    11'b00001100110: data <= 32'h3d96bdd4;
    11'b00001100111: data <= 32'hb4562d7e;
    11'b00001101000: data <= 32'hbdd73943;
    11'b00001101001: data <= 32'hbb283893;
    11'b00001101010: data <= 32'ha9a03958;
    11'b00001101011: data <= 32'hb9d338d3;
    11'b00001101100: data <= 32'hc04cb386;
    11'b00001101101: data <= 32'hc007bc0e;
    11'b00001101110: data <= 32'ha551b613;
    11'b00001101111: data <= 32'h3eba3cce;
    11'b00001110000: data <= 32'h3e4d3f1a;
    11'b00001110001: data <= 32'h38a63a78;
    11'b00001110010: data <= 32'h31392c5e;
    11'b00001110011: data <= 32'h32633a79;
    11'b00001110100: data <= 32'hae453e86;
    11'b00001110101: data <= 32'hb577387c;
    11'b00001110110: data <= 32'h35a9befa;
    11'b00001110111: data <= 32'h3dc4c166;
    11'b00001111000: data <= 32'h3dbdbda3;
    11'b00001111001: data <= 32'h34f433de;
    11'b00001111010: data <= 32'hb4a237cd;
    11'b00001111011: data <= 32'h3486b097;
    11'b00001111100: data <= 32'h3750b4b2;
    11'b00001111101: data <= 32'hbc25acc2;
    11'b00001111110: data <= 32'hc18eb68a;
    11'b00001111111: data <= 32'hc0d7bc09;
    11'b00010000000: data <= 32'hb178b9d6;
    11'b00010000001: data <= 32'h3d7b3584;
    11'b00010000010: data <= 32'h3a653af8;
    11'b00010000011: data <= 32'hb70c383e;
    11'b00010000100: data <= 32'hb87e3936;
    11'b00010000101: data <= 32'h2c5c3f4d;
    11'b00010000110: data <= 32'h2e9440e0;
    11'b00010000111: data <= 32'hb5983b8f;
    11'b00010001000: data <= 32'haea5bdbd;
    11'b00010001001: data <= 32'h3b0dc01e;
    11'b00010001010: data <= 32'h3d9ab82f;
    11'b00010001011: data <= 32'h3c613ae9;
    11'b00010001100: data <= 32'h3bb73745;
    11'b00010001101: data <= 32'h3d55b91f;
    11'b00010001110: data <= 32'h3b93b97d;
    11'b00010001111: data <= 32'hbaeca495;
    11'b00010010000: data <= 32'hc0eab0d8;
    11'b00010010001: data <= 32'hbf6ebc95;
    11'b00010010010: data <= 32'h32e4be60;
    11'b00010010011: data <= 32'h3c87bbb5;
    11'b00010010100: data <= 32'h2290b2fd;
    11'b00010010101: data <= 32'hbcd42e5a;
    11'b00010010110: data <= 32'hbabf39db;
    11'b00010010111: data <= 32'h30893fb6;
    11'b00010011000: data <= 32'ha9eb409f;
    11'b00010011001: data <= 32'hbc7f3ae3;
    11'b00010011010: data <= 32'hbd29bc14;
    11'b00010011011: data <= 32'hac6ebc63;
    11'b00010011100: data <= 32'h3cb037cb;
    11'b00010011101: data <= 32'h3e013d73;
    11'b00010011110: data <= 32'h3e0436cd;
    11'b00010011111: data <= 32'h3e8fb93f;
    11'b00010100000: data <= 32'h3c97b1f1;
    11'b00010100001: data <= 32'hb5b43b33;
    11'b00010100010: data <= 32'hbdf2387b;
    11'b00010100011: data <= 32'hba7bbcb9;
    11'b00010100100: data <= 32'h3a16c0aa;
    11'b00010100101: data <= 32'h3c16bf86;
    11'b00010100110: data <= 32'hb4acbad3;
    11'b00010100111: data <= 32'hbc79b44b;
    11'b00010101000: data <= 32'hb4bf3423;
    11'b00010101001: data <= 32'h38bd3c7e;
    11'b00010101010: data <= 32'hb4b43dbe;
    11'b00010101011: data <= 32'hc037372d;
    11'b00010101100: data <= 32'hc0f0b9da;
    11'b00010101101: data <= 32'hbb06b76d;
    11'b00010101110: data <= 32'h3a7c3abd;
    11'b00010101111: data <= 32'h3ce73cd9;
    11'b00010110000: data <= 32'h3c0e3242;
    11'b00010110001: data <= 32'h3c54b538;
    11'b00010110010: data <= 32'h3bed3ae8;
    11'b00010110011: data <= 32'h31294056;
    11'b00010110100: data <= 32'hb8893d8d;
    11'b00010110101: data <= 32'hae25bbd9;
    11'b00010110110: data <= 32'h3b69c0cf;
    11'b00010110111: data <= 32'h3b5fbf40;
    11'b00010111000: data <= 32'ha8a2b95d;
    11'b00010111001: data <= 32'hb2f9b629;
    11'b00010111010: data <= 32'h3adfb752;
    11'b00010111011: data <= 32'h3d392457;
    11'b00010111100: data <= 32'hb56c382c;
    11'b00010111101: data <= 32'hc12f3042;
    11'b00010111110: data <= 32'hc1bcb8f6;
    11'b00010111111: data <= 32'hbc37b810;
    11'b00011000000: data <= 32'h380c342e;
    11'b00011000001: data <= 32'h37053571;
    11'b00011000010: data <= 32'hb018b4df;
    11'b00011000011: data <= 32'h30a0a8bf;
    11'b00011000100: data <= 32'h39af3ed8;
    11'b00011000101: data <= 32'h36fd41f4;
    11'b00011000110: data <= 32'hb4ac3f64;
    11'b00011000111: data <= 32'hb45db8ff;
    11'b00011001000: data <= 32'h36b0bef1;
    11'b00011001001: data <= 32'h3959ba9f;
    11'b00011001010: data <= 32'h36f43023;
    11'b00011001011: data <= 32'h3ac8b463;
    11'b00011001100: data <= 32'h3fb3bc03;
    11'b00011001101: data <= 32'h3fadb910;
    11'b00011001110: data <= 32'hac6434b6;
    11'b00011001111: data <= 32'hc0713507;
    11'b00011010000: data <= 32'hc073b86d;
    11'b00011010001: data <= 32'hb830bc30;
    11'b00011010010: data <= 32'h3652bab8;
    11'b00011010011: data <= 32'hb61bba2c;
    11'b00011010100: data <= 32'hbc83bb37;
    11'b00011010101: data <= 32'hb6b4aedf;
    11'b00011010110: data <= 32'h39763ef7;
    11'b00011010111: data <= 32'h37744198;
    11'b00011011000: data <= 32'hb9ee3ea8;
    11'b00011011001: data <= 32'hbcf0b4f7;
    11'b00011011010: data <= 32'hb86eb9f4;
    11'b00011011011: data <= 32'h33b4364c;
    11'b00011011100: data <= 32'h39233b3c;
    11'b00011011101: data <= 32'h3d2fb1c4;
    11'b00011011110: data <= 32'h4069bcac;
    11'b00011011111: data <= 32'h4024b736;
    11'b00011100000: data <= 32'h36073bc7;
    11'b00011100001: data <= 32'hbce43c24;
    11'b00011100010: data <= 32'hbbe9b5ea;
    11'b00011100011: data <= 32'h349abe32;
    11'b00011100100: data <= 32'h36c7be96;
    11'b00011100101: data <= 32'hba7abda0;
    11'b00011100110: data <= 32'hbd63bd1e;
    11'b00011100111: data <= 32'hb015b87f;
    11'b00011101000: data <= 32'h3c803b3f;
    11'b00011101001: data <= 32'h37113f08;
    11'b00011101010: data <= 32'hbdd63c05;
    11'b00011101011: data <= 32'hc091b160;
    11'b00011101100: data <= 32'hbd8ba1dc;
    11'b00011101101: data <= 32'hb2003c30;
    11'b00011101110: data <= 32'h355e3c18;
    11'b00011101111: data <= 32'h3a21b60c;
    11'b00011110000: data <= 32'h3e0dbc3b;
    11'b00011110001: data <= 32'h3ecc3506;
    11'b00011110010: data <= 32'h3a02402f;
    11'b00011110011: data <= 32'hb3173f9c;
    11'b00011110100: data <= 32'h2299aac6;
    11'b00011110101: data <= 32'h39e7be27;
    11'b00011110110: data <= 32'h361cbe1d;
    11'b00011110111: data <= 32'hba13bc7f;
    11'b00011111000: data <= 32'hb9f2bce5;
    11'b00011111001: data <= 32'h3ae7bc9a;
    11'b00011111010: data <= 32'h3f89b44b;
    11'b00011111011: data <= 32'h386f388e;
    11'b00011111100: data <= 32'hbf44364b;
    11'b00011111101: data <= 32'hc13eb0a0;
    11'b00011111110: data <= 32'hbdfd3045;
    11'b00011111111: data <= 32'hb5f83a2d;
    11'b00100000000: data <= 32'hb5a23567;
    11'b00100000001: data <= 32'hb6f4bb61;
    11'b00100000010: data <= 32'h3521bba4;
    11'b00100000011: data <= 32'h3c7b3bf9;
    11'b00100000100: data <= 32'h3b4e41aa;
    11'b00100000101: data <= 32'h331940aa;
    11'b00100000110: data <= 32'h30d033b4;
    11'b00100000111: data <= 32'h370dbb74;
    11'b00100001000: data <= 32'h2e24b7cf;
    11'b00100001001: data <= 32'hb7ebae0a;
    11'b00100001010: data <= 32'h3005ba99;
    11'b00100001011: data <= 32'h3f68be45;
    11'b00100001100: data <= 32'h4101bc44;
    11'b00100001101: data <= 32'h3a8d25fc;
    11'b00100001110: data <= 32'hbddf355b;
    11'b00100001111: data <= 32'hbfb4ac3d;
    11'b00100010000: data <= 32'hba21b217;
    11'b00100010001: data <= 32'hb300aeab;
    11'b00100010010: data <= 32'hbc27b97d;
    11'b00100010011: data <= 32'hbe43be37;
    11'b00100010100: data <= 32'hb880bc4b;
    11'b00100010101: data <= 32'h3a9b3c0b;
    11'b00100010110: data <= 32'h3b664134;
    11'b00100010111: data <= 32'ha2903ff0;
    11'b00100011000: data <= 32'hb87e352f;
    11'b00100011001: data <= 32'hb6d0ac4b;
    11'b00100011010: data <= 32'hb62c3ad2;
    11'b00100011011: data <= 32'hb6253bfa;
    11'b00100011100: data <= 32'h3829b714;
    11'b00100011101: data <= 32'h402cbebd;
    11'b00100011110: data <= 32'h4110bc5d;
    11'b00100011111: data <= 32'h3c4e36db;
    11'b00100100000: data <= 32'hb8a43b69;
    11'b00100100001: data <= 32'hb8a231b6;
    11'b00100100010: data <= 32'h35a7b870;
    11'b00100100011: data <= 32'h2f1dba91;
    11'b00100100100: data <= 32'hbd93bd1f;
    11'b00100100101: data <= 32'hbfeebf6b;
    11'b00100100110: data <= 32'hb881bd91;
    11'b00100100111: data <= 32'h3c6e343b;
    11'b00100101000: data <= 32'h3ba63dd9;
    11'b00100101001: data <= 32'hb8853c20;
    11'b00100101010: data <= 32'hbdf1312b;
    11'b00100101011: data <= 32'hbcde3899;
    11'b00100101100: data <= 32'hba433ec7;
    11'b00100101101: data <= 32'hb8e33db5;
    11'b00100101110: data <= 32'h2adbb72b;
    11'b00100101111: data <= 32'h3d3bbe74;
    11'b00100110000: data <= 32'h3f92b814;
    11'b00100110001: data <= 32'h3c9d3d92;
    11'b00100110010: data <= 32'h35193efd;
    11'b00100110011: data <= 32'h38d73804;
    11'b00100110100: data <= 32'h3c86b88c;
    11'b00100110101: data <= 32'h34b7b9e5;
    11'b00100110110: data <= 32'hbd74bb6b;
    11'b00100110111: data <= 32'hbe4bbe47;
    11'b00100111000: data <= 32'h33c6bed3;
    11'b00100111001: data <= 32'h3f3eba6d;
    11'b00100111010: data <= 32'h3c692e5d;
    11'b00100111011: data <= 32'hbb2d2d08;
    11'b00100111100: data <= 32'hbf4faca2;
    11'b00100111101: data <= 32'hbd1939bc;
    11'b00100111110: data <= 32'hba463e7e;
    11'b00100111111: data <= 32'hbc3d3ba4;
    11'b00101000000: data <= 32'hbc2ebb56;
    11'b00101000001: data <= 32'haa2abe3f;
    11'b00101000010: data <= 32'h3bbd2ec6;
    11'b00101000011: data <= 32'h3c214038;
    11'b00101000100: data <= 32'h39e34046;
    11'b00101000101: data <= 32'h3b9f3948;
    11'b00101000110: data <= 32'h3c53b103;
    11'b00101000111: data <= 32'h2f1b32d2;
    11'b00101001000: data <= 32'hbca03407;
    11'b00101001001: data <= 32'hba70baa7;
    11'b00101001010: data <= 32'h3cb9bf4a;
    11'b00101001011: data <= 32'h40ccbe38;
    11'b00101001100: data <= 32'h3d1db94b;
    11'b00101001101: data <= 32'hb98eb430;
    11'b00101001110: data <= 32'hbcd4b032;
    11'b00101001111: data <= 32'hb693372b;
    11'b00101010000: data <= 32'hb4fb3b03;
    11'b00101010001: data <= 32'hbdc82099;
    11'b00101010010: data <= 32'hc03bbe1d;
    11'b00101010011: data <= 32'hbc98be8b;
    11'b00101010100: data <= 32'h35bc330b;
    11'b00101010101: data <= 32'h3aef3fc0;
    11'b00101010110: data <= 32'h385d3eb5;
    11'b00101010111: data <= 32'h3657374a;
    11'b00101011000: data <= 32'h353336b7;
    11'b00101011001: data <= 32'hb59b3df1;
    11'b00101011010: data <= 32'hbc283e3d;
    11'b00101011011: data <= 32'hb5afaf10;
    11'b00101011100: data <= 32'h3dd8bee7;
    11'b00101011101: data <= 32'h40afbe6d;
    11'b00101011110: data <= 32'h3d26b6f2;
    11'b00101011111: data <= 32'hacaf31d3;
    11'b00101100000: data <= 32'h2c872d2e;
    11'b00101100001: data <= 32'h3b5f2ec2;
    11'b00101100010: data <= 32'h35f930b9;
    11'b00101100011: data <= 32'hbe38b8ed;
    11'b00101100100: data <= 32'hc115bf14;
    11'b00101100101: data <= 32'hbd61bf02;
    11'b00101100110: data <= 32'h373bb4a4;
    11'b00101100111: data <= 32'h3abb3aed;
    11'b00101101000: data <= 32'h2815382a;
    11'b00101101001: data <= 32'hb802ac51;
    11'b00101101010: data <= 32'hb7a93a5b;
    11'b00101101011: data <= 32'hb9b540a6;
    11'b00101101100: data <= 32'hbc744068;
    11'b00101101101: data <= 32'hb8f62f5b;
    11'b00101101110: data <= 32'h3a00be42;
    11'b00101101111: data <= 32'h3e10bc48;
    11'b00101110000: data <= 32'h3c0b377f;
    11'b00101110001: data <= 32'h38613bee;
    11'b00101110010: data <= 32'h3cf93637;
    11'b00101110011: data <= 32'h3fb9a242;
    11'b00101110100: data <= 32'h3aa22c58;
    11'b00101110101: data <= 32'hbd99b546;
    11'b00101110110: data <= 32'hc05abd4b;
    11'b00101110111: data <= 32'hb90fbeec;
    11'b00101111000: data <= 32'h3c73bc4f;
    11'b00101111001: data <= 32'h3bd5b7a7;
    11'b00101111010: data <= 32'hb5ceb96d;
    11'b00101111011: data <= 32'hbbbdb8e4;
    11'b00101111100: data <= 32'hb8ce3a36;
    11'b00101111101: data <= 32'hb8b04096;
    11'b00101111110: data <= 32'hbd0a3f6d;
    11'b00101111111: data <= 32'hbdc9b472;
    11'b00110000000: data <= 32'hb8a5be00;
    11'b00110000001: data <= 32'h3569b6c6;
    11'b00110000010: data <= 32'h38613d17;
    11'b00110000011: data <= 32'h3a2b3dc4;
    11'b00110000100: data <= 32'h3e843739;
    11'b00110000101: data <= 32'h40143078;
    11'b00110000110: data <= 32'h3a1a3a1b;
    11'b00110000111: data <= 32'hbcaa3a89;
    11'b00110001000: data <= 32'hbd9ab564;
    11'b00110001001: data <= 32'h35c0bdf2;
    11'b00110001010: data <= 32'h3f05be6e;
    11'b00110001011: data <= 32'h3c5dbd18;
    11'b00110001100: data <= 32'hb604bcd9;
    11'b00110001101: data <= 32'hb8a1bab0;
    11'b00110001110: data <= 32'h33213759;
    11'b00110001111: data <= 32'h2fb53e3c;
    11'b00110010000: data <= 32'hbd1f3b1f;
    11'b00110010001: data <= 32'hc08dbb71;
    11'b00110010010: data <= 32'hbed8be24;
    11'b00110010011: data <= 32'hb7eeb05c;
    11'b00110010100: data <= 32'h314c3d3b;
    11'b00110010101: data <= 32'h38053c1e;
    11'b00110010110: data <= 32'h3c6328a4;
    11'b00110010111: data <= 32'h3d3335c7;
    11'b00110011000: data <= 32'h347b3f25;
    11'b00110011001: data <= 32'hbc1d404d;
    11'b00110011010: data <= 32'hba8a3914;
    11'b00110011011: data <= 32'h3a93bc7f;
    11'b00110011100: data <= 32'h3f06be31;
    11'b00110011101: data <= 32'h3b59bc53;
    11'b00110011110: data <= 32'hada8ba9e;
    11'b00110011111: data <= 32'h3732b911;
    11'b00110100000: data <= 32'h3e4f2eb5;
    11'b00110100001: data <= 32'h3c4a39da;
    11'b00110100010: data <= 32'hbc592ed9;
    11'b00110100011: data <= 32'hc11ebcf6;
    11'b00110100100: data <= 32'hbfcebe05;
    11'b00110100101: data <= 32'hb80bb573;
    11'b00110100110: data <= 32'h2da137b2;
    11'b00110100111: data <= 32'ha6b5b095;
    11'b00110101000: data <= 32'h3043ba17;
    11'b00110101001: data <= 32'h35da367a;
    11'b00110101010: data <= 32'hb11640ea;
    11'b00110101011: data <= 32'hbbf241b0;
    11'b00110101100: data <= 32'hba793c07;
    11'b00110101101: data <= 32'h3597bae8;
    11'b00110101110: data <= 32'h3b66bbda;
    11'b00110101111: data <= 32'h35edb06c;
    11'b00110110000: data <= 32'h31e82d17;
    11'b00110110001: data <= 32'h3dbeb406;
    11'b00110110010: data <= 32'h414aadab;
    11'b00110110011: data <= 32'h3edf36a4;
    11'b00110110100: data <= 32'hba3d3133;
    11'b00110110101: data <= 32'hc049ba76;
    11'b00110110110: data <= 32'hbce0bcea;
    11'b00110110111: data <= 32'h32e3ba34;
    11'b00110111000: data <= 32'h3499b94f;
    11'b00110111001: data <= 32'hb78abda1;
    11'b00110111010: data <= 32'hb844be23;
    11'b00110111011: data <= 32'h261231f4;
    11'b00110111100: data <= 32'hac4640b4;
    11'b00110111101: data <= 32'hbb4b40ff;
    11'b00110111110: data <= 32'hbd2738c6;
    11'b00110111111: data <= 32'hba2bbab1;
    11'b00111000000: data <= 32'hb522b4c5;
    11'b00111000001: data <= 32'hb5ab3aab;
    11'b00111000010: data <= 32'h313839e3;
    11'b00111000011: data <= 32'h3ee8b03e;
    11'b00111000100: data <= 32'h418db02e;
    11'b00111000101: data <= 32'h3eba3a3d;
    11'b00111000110: data <= 32'hb8683c5d;
    11'b00111000111: data <= 32'hbd5633b6;
    11'b00111001000: data <= 32'hadafb99e;
    11'b00111001001: data <= 32'h3c2ebc16;
    11'b00111001010: data <= 32'h3788bd62;
    11'b00111001011: data <= 32'hb925bff4;
    11'b00111001100: data <= 32'hb73ebf5d;
    11'b00111001101: data <= 32'h38feb15e;
    11'b00111001110: data <= 32'h39803e55;
    11'b00111001111: data <= 32'hb9273daf;
    11'b00111010000: data <= 32'hbf3ab315;
    11'b00111010001: data <= 32'hbf15bb9d;
    11'b00111010010: data <= 32'hbce52f6b;
    11'b00111010011: data <= 32'hbafc3c9b;
    11'b00111010100: data <= 32'hb2103866;
    11'b00111010101: data <= 32'h3c9eb89a;
    11'b00111010110: data <= 32'h3fd2b20b;
    11'b00111010111: data <= 32'h3c403de8;
    11'b00111011000: data <= 32'hb7e4408e;
    11'b00111011001: data <= 32'hb9353d32;
    11'b00111011010: data <= 32'h3912b0e1;
    11'b00111011011: data <= 32'h3d1abaa0;
    11'b00111011100: data <= 32'h34b6bc69;
    11'b00111011101: data <= 32'hb8efbe38;
    11'b00111011110: data <= 32'h33dfbe2b;
    11'b00111011111: data <= 32'h3f47b740;
    11'b00111100000: data <= 32'h3ef03967;
    11'b00111100001: data <= 32'hb310366a;
    11'b00111100010: data <= 32'hbfa3ba1b;
    11'b00111100011: data <= 32'hbfcabb8b;
    11'b00111100100: data <= 32'hbce130c6;
    11'b00111100101: data <= 32'hbb3e3938;
    11'b00111100110: data <= 32'hb962b73b;
    11'b00111100111: data <= 32'h3001bde1;
    11'b00111101000: data <= 32'h3a7ab678;
    11'b00111101001: data <= 32'h364c3fb5;
    11'b00111101010: data <= 32'hb80941cb;
    11'b00111101011: data <= 32'hb6eb3ec4;
    11'b00111101100: data <= 32'h37be2fb0;
    11'b00111101101: data <= 32'h3908b459;
    11'b00111101110: data <= 32'hb580ae80;
    11'b00111101111: data <= 32'hb8f7b772;
    11'b00111110000: data <= 32'h3bd9bb89;
    11'b00111110001: data <= 32'h419bb8a2;
    11'b00111110010: data <= 32'h40dd31b0;
    11'b00111110011: data <= 32'h30f63087;
    11'b00111110100: data <= 32'hbdd8b841;
    11'b00111110101: data <= 32'hbca4b8be;
    11'b00111110110: data <= 32'hb5959800;
    11'b00111110111: data <= 32'hb816b2ff;
    11'b00111111000: data <= 32'hbc2abe7f;
    11'b00111111001: data <= 32'hb991c0a6;
    11'b00111111010: data <= 32'h3137b9f9;
    11'b00111111011: data <= 32'h34403eff;
    11'b00111111100: data <= 32'hb60140fe;
    11'b00111111101: data <= 32'hb90f3caa;
    11'b00111111110: data <= 32'hb588a293;
    11'b00111111111: data <= 32'hb81f3569;
    11'b01000000000: data <= 32'hbcb13c02;
    11'b01000000001: data <= 32'hba8637b3;
    11'b01000000010: data <= 32'h3ca3b8b4;
    11'b01000000011: data <= 32'h41c3b91d;
    11'b01000000100: data <= 32'h40a4346e;
    11'b01000000101: data <= 32'h344a3a21;
    11'b01000000110: data <= 32'hb9b13665;
    11'b01000000111: data <= 32'h2d962a99;
    11'b01000001000: data <= 32'h3a09a851;
    11'b01000001001: data <= 32'had67ba02;
    11'b01000001010: data <= 32'hbccfc04f;
    11'b01000001011: data <= 32'hbae3c134;
    11'b01000001100: data <= 32'h3736bc24;
    11'b01000001101: data <= 32'h3b0e3c0f;
    11'b01000001110: data <= 32'h20ee3d42;
    11'b01000001111: data <= 32'hbb3e2e29;
    11'b01000010000: data <= 32'hbca6b5ef;
    11'b01000010001: data <= 32'hbd7c39bf;
    11'b01000010010: data <= 32'hbed53e2f;
    11'b01000010011: data <= 32'hbca438e7;
    11'b01000010100: data <= 32'h38c3baf3;
    11'b01000010101: data <= 32'h3fdfba6b;
    11'b01000010110: data <= 32'h3de939b1;
    11'b01000010111: data <= 32'h2df93ef7;
    11'b01000011000: data <= 32'hacdd3da3;
    11'b01000011001: data <= 32'h3c123947;
    11'b01000011010: data <= 32'h3d3932c2;
    11'b01000011011: data <= 32'hacb3b7c4;
    11'b01000011100: data <= 32'hbd0abe94;
    11'b01000011101: data <= 32'hb6e5c03b;
    11'b01000011110: data <= 32'h3da5bc71;
    11'b01000011111: data <= 32'h3f7f3132;
    11'b01000100000: data <= 32'h38322e7d;
    11'b01000100001: data <= 32'hbb36ba28;
    11'b01000100010: data <= 32'hbd22b896;
    11'b01000100011: data <= 32'hbd383a7e;
    11'b01000100100: data <= 32'hbe653d42;
    11'b01000100101: data <= 32'hbde0b048;
    11'b01000100110: data <= 32'hb61abec8;
    11'b01000100111: data <= 32'h3929bc85;
    11'b01000101000: data <= 32'h37cd3c09;
    11'b01000101001: data <= 32'hb0d6408c;
    11'b01000101010: data <= 32'h31ab3f04;
    11'b01000101011: data <= 32'h3c873abc;
    11'b01000101100: data <= 32'h3b79391c;
    11'b01000101101: data <= 32'hb9023793;
    11'b01000101110: data <= 32'hbd8bb655;
    11'b01000101111: data <= 32'h2f7bbcd1;
    11'b01000110000: data <= 32'h408fbbeb;
    11'b01000110001: data <= 32'h4112b58a;
    11'b01000110010: data <= 32'h3ae4b6ad;
    11'b01000110011: data <= 32'hb83abaad;
    11'b01000110100: data <= 32'hb82bb557;
    11'b01000110101: data <= 32'hb4b43a42;
    11'b01000110110: data <= 32'hbb573943;
    11'b01000110111: data <= 32'hbe5abcaa;
    11'b01000111000: data <= 32'hbcc6c10d;
    11'b01000111001: data <= 32'hb40dbdec;
    11'b01000111010: data <= 32'h29603ad3;
    11'b01000111011: data <= 32'hb13c3f81;
    11'b01000111100: data <= 32'h2db73c70;
    11'b01000111101: data <= 32'h384b374b;
    11'b01000111110: data <= 32'ha9d33c0d;
    11'b01000111111: data <= 32'hbdbe3e3a;
    11'b01001000000: data <= 32'hbe873a59;
    11'b01001000001: data <= 32'h3444b81f;
    11'b01001000010: data <= 32'h40aebafe;
    11'b01001000011: data <= 32'h40a8b577;
    11'b01001000100: data <= 32'h3a1ca970;
    11'b01001000101: data <= 32'h21b8ae1b;
    11'b01001000110: data <= 32'h399e3495;
    11'b01001000111: data <= 32'h3c293aaf;
    11'b01001001000: data <= 32'hb0b63262;
    11'b01001001001: data <= 32'hbe2cbea7;
    11'b01001001010: data <= 32'hbdb9c176;
    11'b01001001011: data <= 32'hb33abe6f;
    11'b01001001100: data <= 32'h36f334b5;
    11'b01001001101: data <= 32'h31d439b9;
    11'b01001001110: data <= 32'hace1b1bc;
    11'b01001001111: data <= 32'hb142b3d8;
    11'b01001010000: data <= 32'hbacc3cac;
    11'b01001010001: data <= 32'hbfb5404e;
    11'b01001010010: data <= 32'hbf793cc5;
    11'b01001010011: data <= 32'hb135b851;
    11'b01001010100: data <= 32'h3dc6bbc7;
    11'b01001010101: data <= 32'h3d23a630;
    11'b01001010110: data <= 32'h341b3a41;
    11'b01001010111: data <= 32'h36963ab9;
    11'b01001011000: data <= 32'h3eaf3afe;
    11'b01001011001: data <= 32'h3f763c1b;
    11'b01001011010: data <= 32'h30d535ff;
    11'b01001011011: data <= 32'hbe06bca7;
    11'b01001011100: data <= 32'hbc78c023;
    11'b01001011101: data <= 32'h386ebd7e;
    11'b01001011110: data <= 32'h3d50b530;
    11'b01001011111: data <= 32'h3987b835;
    11'b01001100000: data <= 32'hace4bd4a;
    11'b01001100001: data <= 32'hb548ba1b;
    11'b01001100010: data <= 32'hba4e3c88;
    11'b01001100011: data <= 32'hbeb1400f;
    11'b01001100100: data <= 32'hbf9b3933;
    11'b01001100101: data <= 32'hbb54bcf5;
    11'b01001100110: data <= 32'h2e63bd2f;
    11'b01001100111: data <= 32'h2378339c;
    11'b01001101000: data <= 32'hb53d3d42;
    11'b01001101001: data <= 32'h380b3cbc;
    11'b01001101010: data <= 32'h3f8a3b96;
    11'b01001101011: data <= 32'h3ee23ce7;
    11'b01001101100: data <= 32'hb3c13c86;
    11'b01001101101: data <= 32'hbe7b2e74;
    11'b01001101110: data <= 32'hb913bb13;
    11'b01001101111: data <= 32'h3d89bb2e;
    11'b01001110000: data <= 32'h3febb92d;
    11'b01001110001: data <= 32'h3ba3bc8b;
    11'b01001110010: data <= 32'h2fbcbe8e;
    11'b01001110011: data <= 32'h3429b9c3;
    11'b01001110100: data <= 32'h336f3c4e;
    11'b01001110101: data <= 32'hb9e13dd4;
    11'b01001110110: data <= 32'hbea7b4f5;
    11'b01001110111: data <= 32'hbe17c018;
    11'b01001111000: data <= 32'hbb0ebe6b;
    11'b01001111001: data <= 32'hb9a5328e;
    11'b01001111010: data <= 32'hb89f3c38;
    11'b01001111011: data <= 32'h35dd3846;
    11'b01001111100: data <= 32'h3d8c354c;
    11'b01001111101: data <= 32'h3ac63d06;
    11'b01001111110: data <= 32'hbc0e4000;
    11'b01001111111: data <= 32'hbf633d75;
    11'b01010000000: data <= 32'hb68c2e49;
    11'b01010000001: data <= 32'h3e33b804;
    11'b01010000010: data <= 32'h3f16b87d;
    11'b01010000011: data <= 32'h3943baef;
    11'b01010000100: data <= 32'h3580bc29;
    11'b01010000101: data <= 32'h3d16b125;
    11'b01010000110: data <= 32'h3e8a3c80;
    11'b01010000111: data <= 32'h35733bba;
    11'b01010001000: data <= 32'hbd37bb07;
    11'b01010001001: data <= 32'hbe97c084;
    11'b01010001010: data <= 32'hbbb5be48;
    11'b01010001011: data <= 32'hb7daacb3;
    11'b01010001100: data <= 32'hb5352e0c;
    11'b01010001101: data <= 32'h3279ba87;
    11'b01010001110: data <= 32'h3984b96c;
    11'b01010001111: data <= 32'h18dd3c49;
    11'b01010010000: data <= 32'hbe1140e9;
    11'b01010010001: data <= 32'hbfd83f7f;
    11'b01010010010: data <= 32'hb8cb349b;
    11'b01010010011: data <= 32'h3ab1b772;
    11'b01010010100: data <= 32'h3962b399;
    11'b01010010101: data <= 32'hb0d0ace2;
    11'b01010010110: data <= 32'h3648ae35;
    11'b01010010111: data <= 32'h4029370c;
    11'b01010011000: data <= 32'h41243cef;
    11'b01010011001: data <= 32'h3b1a3b93;
    11'b01010011010: data <= 32'hbc57b85c;
    11'b01010011011: data <= 32'hbd3cbe37;
    11'b01010011100: data <= 32'hb3b8bc34;
    11'b01010011101: data <= 32'h35fbb572;
    11'b01010011110: data <= 32'h320ebbcd;
    11'b01010011111: data <= 32'h30ebc025;
    11'b01010100000: data <= 32'h3601bde7;
    11'b01010100001: data <= 32'had693a7d;
    11'b01010100010: data <= 32'hbcf44092;
    11'b01010100011: data <= 32'hbef43da1;
    11'b01010100100: data <= 32'hbc0db582;
    11'b01010100101: data <= 32'hb54aba38;
    11'b01010100110: data <= 32'hb9b32a54;
    11'b01010100111: data <= 32'hbc2a387d;
    11'b01010101000: data <= 32'h331135f7;
    11'b01010101001: data <= 32'h40723813;
    11'b01010101010: data <= 32'h41093cdc;
    11'b01010101011: data <= 32'h38d33d8b;
    11'b01010101100: data <= 32'hbca43852;
    11'b01010101101: data <= 32'hba80b41f;
    11'b01010101110: data <= 32'h393fb3ff;
    11'b01010101111: data <= 32'h3c83b5cf;
    11'b01010110000: data <= 32'h376fbdfb;
    11'b01010110001: data <= 32'h319ec0ff;
    11'b01010110010: data <= 32'h3970be58;
    11'b01010110011: data <= 32'h3a13396e;
    11'b01010110100: data <= 32'hb25e3ecd;
    11'b01010110101: data <= 32'hbcae3696;
    11'b01010110110: data <= 32'hbd2dbce9;
    11'b01010110111: data <= 32'hbcd1bc6e;
    11'b01010111000: data <= 32'hbe3b30d3;
    11'b01010111001: data <= 32'hbdf73868;
    11'b01010111010: data <= 32'ha885aebf;
    11'b01010111011: data <= 32'h3ed6b221;
    11'b01010111100: data <= 32'h3e8c3b68;
    11'b01010111101: data <= 32'hb2ec3fab;
    11'b01010111110: data <= 32'hbda53eba;
    11'b01010111111: data <= 32'hb7d13aec;
    11'b01011000000: data <= 32'h3c233644;
    11'b01011000001: data <= 32'h3c56af56;
    11'b01011000010: data <= 32'h2ec7bccc;
    11'b01011000011: data <= 32'h2e71bfb0;
    11'b01011000100: data <= 32'h3d6bbc0e;
    11'b01011000101: data <= 32'h400f39fa;
    11'b01011000110: data <= 32'h3c193c8e;
    11'b01011000111: data <= 32'hb832b55e;
    11'b01011001000: data <= 32'hbcd8be62;
    11'b01011001001: data <= 32'hbcfdbc24;
    11'b01011001010: data <= 32'hbd973076;
    11'b01011001011: data <= 32'hbd15ad72;
    11'b01011001100: data <= 32'hb250bd44;
    11'b01011001101: data <= 32'h3bb2bd67;
    11'b01011001110: data <= 32'h392b36d1;
    11'b01011001111: data <= 32'hbaf14040;
    11'b01011010000: data <= 32'hbe0d4047;
    11'b01011010001: data <= 32'hb7273c8f;
    11'b01011010010: data <= 32'h39073818;
    11'b01011010011: data <= 32'h3025338c;
    11'b01011010100: data <= 32'hbac6b5f9;
    11'b01011010101: data <= 32'hb1c4baed;
    11'b01011010110: data <= 32'h3f8bb46e;
    11'b01011010111: data <= 32'h41cd3aeb;
    11'b01011011000: data <= 32'h3ebe3b66;
    11'b01011011001: data <= 32'hb15fb4a1;
    11'b01011011010: data <= 32'hba75bc2a;
    11'b01011011011: data <= 32'hb7edb626;
    11'b01011011100: data <= 32'hb7453290;
    11'b01011011101: data <= 32'hb923badf;
    11'b01011011110: data <= 32'hb313c100;
    11'b01011011111: data <= 32'h37d4c093;
    11'b01011100000: data <= 32'h34b1a67c;
    11'b01011100001: data <= 32'hb9fc3f63;
    11'b01011100010: data <= 32'hbcb83e91;
    11'b01011100011: data <= 32'hb8493774;
    11'b01011100100: data <= 32'hb3722f98;
    11'b01011100101: data <= 32'hbcb437e8;
    11'b01011100110: data <= 32'hbf98363d;
    11'b01011100111: data <= 32'hb8b8b0f0;
    11'b01011101000: data <= 32'h3f86a92e;
    11'b01011101001: data <= 32'h41a13a21;
    11'b01011101010: data <= 32'h3d963c3c;
    11'b01011101011: data <= 32'hb48237c5;
    11'b01011101100: data <= 32'hb5463157;
    11'b01011101101: data <= 32'h380538bd;
    11'b01011101110: data <= 32'h381d375c;
    11'b01011101111: data <= 32'hb241bcc7;
    11'b01011110000: data <= 32'hb3ebc1c9;
    11'b01011110001: data <= 32'h3822c0dd;
    11'b01011110010: data <= 32'h3aa1b159;
    11'b01011110011: data <= 32'h321f3d0b;
    11'b01011110100: data <= 32'hb6ee3882;
    11'b01011110101: data <= 32'hb815b8d6;
    11'b01011110110: data <= 32'hbb21b614;
    11'b01011110111: data <= 32'hbff838ed;
    11'b01011111000: data <= 32'hc0da3900;
    11'b01011111001: data <= 32'hbb47b548;
    11'b01011111010: data <= 32'h3d5ab900;
    11'b01011111011: data <= 32'h3f7634e7;
    11'b01011111100: data <= 32'h36be3d10;
    11'b01011111101: data <= 32'hb9843d8b;
    11'b01011111110: data <= 32'h9d7e3d0a;
    11'b01011111111: data <= 32'h3c623d69;
    11'b01100000000: data <= 32'h3a1b3aa1;
    11'b01100000001: data <= 32'hb6b8bab9;
    11'b01100000010: data <= 32'hb78cc086;
    11'b01100000011: data <= 32'h3aecbef6;
    11'b01100000100: data <= 32'h3f5a28b1;
    11'b01100000101: data <= 32'h3d8839ad;
    11'b01100000110: data <= 32'h35dfb5f5;
    11'b01100000111: data <= 32'hb405bd04;
    11'b01100001000: data <= 32'hbabeb755;
    11'b01100001001: data <= 32'hbf2839d0;
    11'b01100001010: data <= 32'hc04234e8;
    11'b01100001011: data <= 32'hbbbfbd12;
    11'b01100001100: data <= 32'h38d5befa;
    11'b01100001101: data <= 32'h39abb5f0;
    11'b01100001110: data <= 32'hb8003d00;
    11'b01100001111: data <= 32'hbba83edf;
    11'b01100010000: data <= 32'h302a3e06;
    11'b01100010001: data <= 32'h3bf03dc8;
    11'b01100010010: data <= 32'h2dc73c7a;
    11'b01100010011: data <= 32'hbd48a519;
    11'b01100010100: data <= 32'hbb8abc3e;
    11'b01100010101: data <= 32'h3c8aba00;
    11'b01100010110: data <= 32'h411c3550;
    11'b01100010111: data <= 32'h400d36e0;
    11'b01100011000: data <= 32'h39fdb8e5;
    11'b01100011001: data <= 32'h30aebbea;
    11'b01100011010: data <= 32'had2d2fec;
    11'b01100011011: data <= 32'hb9ca3bdc;
    11'b01100011100: data <= 32'hbd15b1d2;
    11'b01100011101: data <= 32'hba7fc08c;
    11'b01100011110: data <= 32'h2dcdc159;
    11'b01100011111: data <= 32'h2dadbb2c;
    11'b01100100000: data <= 32'hb96c3b5f;
    11'b01100100001: data <= 32'hb9ba3cc2;
    11'b01100100010: data <= 32'h331939dc;
    11'b01100100011: data <= 32'h36e63adf;
    11'b01100100100: data <= 32'hbc123cd5;
    11'b01100100101: data <= 32'hc0be3a1f;
    11'b01100100110: data <= 32'hbde1ae7d;
    11'b01100100111: data <= 32'h3c1bb2b7;
    11'b01100101000: data <= 32'h40d4359f;
    11'b01100101001: data <= 32'h3ea4366c;
    11'b01100101010: data <= 32'h37c1b09b;
    11'b01100101011: data <= 32'h37aa1aa8;
    11'b01100101100: data <= 32'h3b6f3c68;
    11'b01100101101: data <= 32'h378f3d90;
    11'b01100101110: data <= 32'hb827b5d8;
    11'b01100101111: data <= 32'hb98bc12d;
    11'b01100110000: data <= 32'ha4eac188;
    11'b01100110001: data <= 32'h350bbb82;
    11'b01100110010: data <= 32'h268e371a;
    11'b01100110011: data <= 32'h26c42e59;
    11'b01100110100: data <= 32'h36d4b85c;
    11'b01100110101: data <= 32'ha85d2bf1;
    11'b01100110110: data <= 32'hbef33ca8;
    11'b01100110111: data <= 32'hc1be3c71;
    11'b01100111000: data <= 32'hbef92718;
    11'b01100111001: data <= 32'h3865b84b;
    11'b01100111010: data <= 32'h3dc8ad80;
    11'b01100111011: data <= 32'h37fb36a9;
    11'b01100111100: data <= 32'hb291383b;
    11'b01100111101: data <= 32'h39043bdc;
    11'b01100111110: data <= 32'h3e6f3f70;
    11'b01100111111: data <= 32'h3c133f14;
    11'b01101000000: data <= 32'hb773a79b;
    11'b01101000001: data <= 32'hbaf4bfb9;
    11'b01101000010: data <= 32'h3065bfa5;
    11'b01101000011: data <= 32'h3c47b7a5;
    11'b01101000100: data <= 32'h3c552c50;
    11'b01101000101: data <= 32'h3abdbb3f;
    11'b01101000110: data <= 32'h39ffbdf0;
    11'b01101000111: data <= 32'h29b7b501;
    11'b01101001000: data <= 32'hbdff3cca;
    11'b01101001001: data <= 32'hc0e23bc9;
    11'b01101001010: data <= 32'hbe53b918;
    11'b01101001011: data <= 32'ha59fbdff;
    11'b01101001100: data <= 32'h3361ba50;
    11'b01101001101: data <= 32'hb9a234a3;
    11'b01101001110: data <= 32'hba443a43;
    11'b01101001111: data <= 32'h39403cbd;
    11'b01101010000: data <= 32'h3eaf3f6d;
    11'b01101010001: data <= 32'h390d3f8b;
    11'b01101010010: data <= 32'hbcbe3932;
    11'b01101010011: data <= 32'hbd74b96e;
    11'b01101010100: data <= 32'h3436b935;
    11'b01101010101: data <= 32'h3ea93062;
    11'b01101010110: data <= 32'h3eb1ad2d;
    11'b01101010111: data <= 32'h3caabd2e;
    11'b01101011000: data <= 32'h3c1dbe10;
    11'b01101011001: data <= 32'h39932c07;
    11'b01101011010: data <= 32'hb63b3ddd;
    11'b01101011011: data <= 32'hbd553933;
    11'b01101011100: data <= 32'hbc6cbdf1;
    11'b01101011101: data <= 32'hb626c0ba;
    11'b01101011110: data <= 32'hb831bd2a;
    11'b01101011111: data <= 32'hbcc12576;
    11'b01101100000: data <= 32'hba393534;
    11'b01101100001: data <= 32'h39ef35e9;
    11'b01101100010: data <= 32'h3d253c2e;
    11'b01101100011: data <= 32'hb4a23eaf;
    11'b01101100100: data <= 32'hc0513d17;
    11'b01101100101: data <= 32'hbf953669;
    11'b01101100110: data <= 32'h31153292;
    11'b01101100111: data <= 32'h3e3736c7;
    11'b01101101000: data <= 32'h3d11acfa;
    11'b01101101001: data <= 32'h39b3bc08;
    11'b01101101010: data <= 32'h3c59b9e4;
    11'b01101101011: data <= 32'h3e303b94;
    11'b01101101100: data <= 32'h3b513f99;
    11'b01101101101: data <= 32'hb4303815;
    11'b01101101110: data <= 32'hb986bf2a;
    11'b01101101111: data <= 32'hb6edc0d6;
    11'b01101110000: data <= 32'hb7a5bcba;
    11'b01101110001: data <= 32'hb9ceb321;
    11'b01101110010: data <= 32'hb0dfb8f2;
    11'b01101110011: data <= 32'h3bddbc05;
    11'b01101110100: data <= 32'h3b3fac50;
    11'b01101110101: data <= 32'hbbb83d3c;
    11'b01101110110: data <= 32'hc13f3e1c;
    11'b01101110111: data <= 32'hc01e39a3;
    11'b01101111000: data <= 32'hb04230aa;
    11'b01101111001: data <= 32'h39b13048;
    11'b01101111010: data <= 32'h246fae4e;
    11'b01101111011: data <= 32'hb481b73f;
    11'b01101111100: data <= 32'h3b443146;
    11'b01101111101: data <= 32'h40393eb1;
    11'b01101111110: data <= 32'h3e84406c;
    11'b01101111111: data <= 32'h2d6939b2;
    11'b01110000000: data <= 32'hb973bcef;
    11'b01110000001: data <= 32'hb4ccbdf0;
    11'b01110000010: data <= 32'h304fb6ff;
    11'b01110000011: data <= 32'h3310b46f;
    11'b01110000100: data <= 32'h390cbdfc;
    11'b01110000101: data <= 32'h3d1ec036;
    11'b01110000110: data <= 32'h3b39ba0c;
    11'b01110000111: data <= 32'hba693c79;
    11'b01110001000: data <= 32'hc0423d91;
    11'b01110001001: data <= 32'hbe923257;
    11'b01110001010: data <= 32'hb65fb95f;
    11'b01110001011: data <= 32'hb5f6b834;
    11'b01110001100: data <= 32'hbd5fb361;
    11'b01110001101: data <= 32'hbcc3b164;
    11'b01110001110: data <= 32'h396e36a6;
    11'b01110001111: data <= 32'h404d3e7c;
    11'b01110010000: data <= 32'h3da34039;
    11'b01110010001: data <= 32'hb74d3c72;
    11'b01110010010: data <= 32'hbc72af17;
    11'b01110010011: data <= 32'hb260ac9f;
    11'b01110010100: data <= 32'h39b93827;
    11'b01110010101: data <= 32'h3aa6b066;
    11'b01110010110: data <= 32'h3b61bf5c;
    11'b01110010111: data <= 32'h3d8fc0a0;
    11'b01110011000: data <= 32'h3d41b8c1;
    11'b01110011001: data <= 32'h31f63d2d;
    11'b01110011010: data <= 32'hbb063c67;
    11'b01110011011: data <= 32'hba96b8c9;
    11'b01110011100: data <= 32'hb73abe1d;
    11'b01110011101: data <= 32'hbc40bc08;
    11'b01110011110: data <= 32'hc005b610;
    11'b01110011111: data <= 32'hbdbdb6de;
    11'b01110100000: data <= 32'h3918b49c;
    11'b01110100001: data <= 32'h3f303978;
    11'b01110100010: data <= 32'h388f3e42;
    11'b01110100011: data <= 32'hbd923daa;
    11'b01110100100: data <= 32'hbe853b1d;
    11'b01110100101: data <= 32'hb3493bd0;
    11'b01110100110: data <= 32'h3a073c5f;
    11'b01110100111: data <= 32'h382e2818;
    11'b01110101000: data <= 32'h35d0be4c;
    11'b01110101001: data <= 32'h3c8fbe90;
    11'b01110101010: data <= 32'h3f633316;
    11'b01110101011: data <= 32'h3d993eda;
    11'b01110101100: data <= 32'h36433b60;
    11'b01110101101: data <= 32'had98bc09;
    11'b01110101110: data <= 32'hb4b1bea7;
    11'b01110101111: data <= 32'hbc19ba8a;
    11'b01110110000: data <= 32'hbeb9b5a1;
    11'b01110110001: data <= 32'hbb4fbc4b;
    11'b01110110010: data <= 32'h3ad4be44;
    11'b01110110011: data <= 32'h3d9eb902;
    11'b01110110100: data <= 32'hb1713ada;
    11'b01110110101: data <= 32'hbfb23db4;
    11'b01110110110: data <= 32'hbef33cbe;
    11'b01110110111: data <= 32'hb4a63c4b;
    11'b01110111000: data <= 32'h31dc3b9a;
    11'b01110111001: data <= 32'hb90c2b20;
    11'b01110111010: data <= 32'hba90bc1a;
    11'b01110111011: data <= 32'h38d4b9b1;
    11'b01110111100: data <= 32'h40473bfd;
    11'b01110111101: data <= 32'h402e3ff7;
    11'b01110111110: data <= 32'h3b573b83;
    11'b01110111111: data <= 32'h2f67b988;
    11'b01111000000: data <= 32'had66ba99;
    11'b01111000001: data <= 32'hb6df2ea1;
    11'b01111000010: data <= 32'hb9efaa5f;
    11'b01111000011: data <= 32'hae56bea5;
    11'b01111000100: data <= 32'h3c8bc144;
    11'b01111000101: data <= 32'h3d0bbe0e;
    11'b01111000110: data <= 32'hb2de36cc;
    11'b01111000111: data <= 32'hbe173cb4;
    11'b01111001000: data <= 32'hbca73998;
    11'b01111001001: data <= 32'hb2cf34cc;
    11'b01111001010: data <= 32'hb8d73497;
    11'b01111001011: data <= 32'hbfcbacb8;
    11'b01111001100: data <= 32'hbfc7b924;
    11'b01111001101: data <= 32'h2dc8b494;
    11'b01111001110: data <= 32'h400c3c2b;
    11'b01111001111: data <= 32'h3f8d3f0e;
    11'b01111010000: data <= 32'h37453c15;
    11'b01111010001: data <= 32'hb47f3071;
    11'b01111010010: data <= 32'h25233853;
    11'b01111010011: data <= 32'h32de3d26;
    11'b01111010100: data <= 32'h20513689;
    11'b01111010101: data <= 32'h349abf42;
    11'b01111010110: data <= 32'h3c9ac1b3;
    11'b01111010111: data <= 32'h3d8cbddb;
    11'b01111011000: data <= 32'h37db382f;
    11'b01111011001: data <= 32'hb5303af1;
    11'b01111011010: data <= 32'haf50b053;
    11'b01111011011: data <= 32'h2d02b94b;
    11'b01111011100: data <= 32'hbc4db494;
    11'b01111011101: data <= 32'hc140b11b;
    11'b01111011110: data <= 32'hc0abb946;
    11'b01111011111: data <= 32'hacf0b9ca;
    11'b01111100000: data <= 32'h3e833153;
    11'b01111100001: data <= 32'h3c1c3bf0;
    11'b01111100010: data <= 32'hb86a3bba;
    11'b01111100011: data <= 32'hbb073b2b;
    11'b01111100100: data <= 32'h27063e63;
    11'b01111100101: data <= 32'h37474015;
    11'b01111100110: data <= 32'haafd3a08;
    11'b01111100111: data <= 32'hb251bde9;
    11'b01111101000: data <= 32'h3994c057;
    11'b01111101001: data <= 32'h3e3fb8e7;
    11'b01111101010: data <= 32'h3dc93c01;
    11'b01111101011: data <= 32'h3b9b395c;
    11'b01111101100: data <= 32'h3ab0b9ac;
    11'b01111101101: data <= 32'h376cbc14;
    11'b01111101110: data <= 32'hbb7bb1cb;
    11'b01111101111: data <= 32'hc0982974;
    11'b01111110000: data <= 32'hbf45bbae;
    11'b01111110001: data <= 32'h3176bef2;
    11'b01111110010: data <= 32'h3ce5bc93;
    11'b01111110011: data <= 32'h310629ec;
    11'b01111110100: data <= 32'hbd22399d;
    11'b01111110101: data <= 32'hbc523c3c;
    11'b01111110110: data <= 32'h2ecf3ed5;
    11'b01111110111: data <= 32'h32853fca;
    11'b01111111000: data <= 32'hbb893a47;
    11'b01111111001: data <= 32'hbd7ebb57;
    11'b01111111010: data <= 32'hadb5bc8d;
    11'b01111111011: data <= 32'h3e2c3573;
    11'b01111111100: data <= 32'h3fe53d87;
    11'b01111111101: data <= 32'h3e0038a0;
    11'b01111111110: data <= 32'h3c8ab974;
    11'b01111111111: data <= 32'h39d2b715;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    