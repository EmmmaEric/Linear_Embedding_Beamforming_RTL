
module memory_rom_46(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3ab13d5d;
    11'b00000000001: data <= 32'h385039f4;
    11'b00000000010: data <= 32'hb751ba41;
    11'b00000000011: data <= 32'hb215bf73;
    11'b00000000100: data <= 32'h3d66bc48;
    11'b00000000101: data <= 32'h40833925;
    11'b00000000110: data <= 32'h3e563be9;
    11'b00000000111: data <= 32'h365fb5e7;
    11'b00000001000: data <= 32'hb401bd4f;
    11'b00000001001: data <= 32'hb9e9b8b4;
    11'b00000001010: data <= 32'hbdee3618;
    11'b00000001011: data <= 32'hbe86b480;
    11'b00000001100: data <= 32'hb7b7bf5e;
    11'b00000001101: data <= 32'h3a6ac00a;
    11'b00000001110: data <= 32'h3843b579;
    11'b00000001111: data <= 32'hbaf03d60;
    11'b00000010000: data <= 32'hbd483eab;
    11'b00000010001: data <= 32'hb4213d1f;
    11'b00000010010: data <= 32'h37673c8b;
    11'b00000010011: data <= 32'hb7bf3ae5;
    11'b00000010100: data <= 32'hbe8dac35;
    11'b00000010101: data <= 32'hbacaba4b;
    11'b00000010110: data <= 32'h3db7b35b;
    11'b00000010111: data <= 32'h41683b0f;
    11'b00000011000: data <= 32'h3faa3aff;
    11'b00000011001: data <= 32'h3865b30b;
    11'b00000011010: data <= 32'h2cb0b8d0;
    11'b00000011011: data <= 32'h2c0e35a1;
    11'b00000011100: data <= 32'hb5d93ab4;
    11'b00000011101: data <= 32'hb9fbb91c;
    11'b00000011110: data <= 32'hb3d4c15e;
    11'b00000011111: data <= 32'h3854c184;
    11'b00000100000: data <= 32'h35a1ba0d;
    11'b00000100001: data <= 32'hb8733bae;
    11'b00000100010: data <= 32'hb9cd3b95;
    11'b00000100011: data <= 32'ha64334b3;
    11'b00000100100: data <= 32'hadef3629;
    11'b00000100101: data <= 32'hbe613a4a;
    11'b00000100110: data <= 32'hc153372b;
    11'b00000100111: data <= 32'hbd9bb387;
    11'b00000101000: data <= 32'h3c98afa9;
    11'b00000101001: data <= 32'h40853906;
    11'b00000101010: data <= 32'h3ced3a91;
    11'b00000101011: data <= 32'h2a5a3671;
    11'b00000101100: data <= 32'h337a389e;
    11'b00000101101: data <= 32'h3ae83de0;
    11'b00000101110: data <= 32'h38413d8b;
    11'b00000101111: data <= 32'hb4c6b8ad;
    11'b00000110000: data <= 32'hb445c14f;
    11'b00000110001: data <= 32'h3862c102;
    11'b00000110010: data <= 32'h3b1fb88d;
    11'b00000110011: data <= 32'h37e138b7;
    11'b00000110100: data <= 32'h347dabd6;
    11'b00000110101: data <= 32'h3616baca;
    11'b00000110110: data <= 32'hb53bb45c;
    11'b00000110111: data <= 32'hc00839ea;
    11'b00000111000: data <= 32'hc1c03868;
    11'b00000111001: data <= 32'hbe17b845;
    11'b00000111010: data <= 32'h394bbb1e;
    11'b00000111011: data <= 32'h3cd7b00b;
    11'b00000111100: data <= 32'h25e13935;
    11'b00000111101: data <= 32'hb94a3b6b;
    11'b00000111110: data <= 32'h34433d85;
    11'b00000111111: data <= 32'h3ceb4022;
    11'b00001000000: data <= 32'h38db3ef0;
    11'b00001000001: data <= 32'hb9a2aedf;
    11'b00001000010: data <= 32'hb9ddbf0c;
    11'b00001000011: data <= 32'h38ddbdca;
    11'b00001000100: data <= 32'h3e9127fc;
    11'b00001000101: data <= 32'h3e2d3616;
    11'b00001000110: data <= 32'h3c63ba17;
    11'b00001000111: data <= 32'h3a6cbd70;
    11'b00001001000: data <= 32'h1a64b406;
    11'b00001001001: data <= 32'hbdc13bbf;
    11'b00001001010: data <= 32'hc04d35f3;
    11'b00001001011: data <= 32'hbcafbd7c;
    11'b00001001100: data <= 32'h3397c00d;
    11'b00001001101: data <= 32'h32cdbbd2;
    11'b00001001110: data <= 32'hbafd3543;
    11'b00001001111: data <= 32'hbbc43b04;
    11'b00001010000: data <= 32'h35c03cdb;
    11'b00001010001: data <= 32'h3c673f0a;
    11'b00001010010: data <= 32'haf843ec4;
    11'b00001010011: data <= 32'hbeff381c;
    11'b00001010100: data <= 32'hbde5b8a8;
    11'b00001010101: data <= 32'h3811b529;
    11'b00001010110: data <= 32'h3fd53847;
    11'b00001010111: data <= 32'h3f4934ca;
    11'b00001011000: data <= 32'h3cc0babb;
    11'b00001011001: data <= 32'h3c11bb89;
    11'b00001011010: data <= 32'h39da3848;
    11'b00001011011: data <= 32'hb35b3e0b;
    11'b00001011100: data <= 32'hbc003337;
    11'b00001011101: data <= 32'hb94cc018;
    11'b00001011110: data <= 32'h2898c16a;
    11'b00001011111: data <= 32'hb1c1bd7e;
    11'b00001100000: data <= 32'hbb079ab8;
    11'b00001100001: data <= 32'hb866326f;
    11'b00001100010: data <= 32'h395f30b5;
    11'b00001100011: data <= 32'h3a393a25;
    11'b00001100100: data <= 32'hbc203d66;
    11'b00001100101: data <= 32'hc16c3b96;
    11'b00001100110: data <= 32'hc017312f;
    11'b00001100111: data <= 32'h33162f17;
    11'b00001101000: data <= 32'h3e1637b8;
    11'b00001101001: data <= 32'h3c4031e1;
    11'b00001101010: data <= 32'h37adb769;
    11'b00001101011: data <= 32'h3b73238e;
    11'b00001101100: data <= 32'h3dc53e56;
    11'b00001101101: data <= 32'h3abc4039;
    11'b00001101110: data <= 32'hb32f3575;
    11'b00001101111: data <= 32'hb746bff5;
    11'b00001110000: data <= 32'h1d97c0c6;
    11'b00001110001: data <= 32'h2f13bc10;
    11'b00001110010: data <= 32'hace4b122;
    11'b00001110011: data <= 32'h3607b9c4;
    11'b00001110100: data <= 32'h3c9fbc9d;
    11'b00001110101: data <= 32'h393cb2db;
    11'b00001110110: data <= 32'hbd8f3c32;
    11'b00001110111: data <= 32'hc1bc3c3c;
    11'b00001111000: data <= 32'hc0152ee9;
    11'b00001111001: data <= 32'hae03b63a;
    11'b00001111010: data <= 32'h3861b195;
    11'b00001111011: data <= 32'hb4a5ad23;
    11'b00001111100: data <= 32'hb860addd;
    11'b00001111101: data <= 32'h398e39ca;
    11'b00001111110: data <= 32'h3f284047;
    11'b00001111111: data <= 32'h3c9d40c4;
    11'b00010000000: data <= 32'hb56c3991;
    11'b00010000001: data <= 32'hba5ebc9c;
    11'b00010000010: data <= 32'ha7babcca;
    11'b00010000011: data <= 32'h3967af66;
    11'b00010000100: data <= 32'h3aceae12;
    11'b00010000101: data <= 32'h3ca3bd87;
    11'b00010000110: data <= 32'h3e33bf92;
    11'b00010000111: data <= 32'h3b52b808;
    11'b00010001000: data <= 32'hbaca3c7d;
    11'b00010001001: data <= 32'hc00e3bb8;
    11'b00010001010: data <= 32'hbda8b829;
    11'b00010001011: data <= 32'hb401bd7d;
    11'b00010001100: data <= 32'hb662bbf4;
    11'b00010001101: data <= 32'hbda2b6b7;
    11'b00010001110: data <= 32'hbcbdb017;
    11'b00010001111: data <= 32'h38cb3894;
    11'b00010010000: data <= 32'h3ee93ef1;
    11'b00010010001: data <= 32'h39364033;
    11'b00010010010: data <= 32'hbcce3c44;
    11'b00010010011: data <= 32'hbdffa78c;
    11'b00010010100: data <= 32'hb1d33089;
    11'b00010010101: data <= 32'h3ba339d7;
    11'b00010010110: data <= 32'h3c79297c;
    11'b00010010111: data <= 32'h3cb4be09;
    11'b00010011000: data <= 32'h3e49bed4;
    11'b00010011001: data <= 32'h3db22c96;
    11'b00010011010: data <= 32'h34d83e73;
    11'b00010011011: data <= 32'hb9623b26;
    11'b00010011100: data <= 32'hb873bc75;
    11'b00010011101: data <= 32'hb2a0c009;
    11'b00010011110: data <= 32'hba8bbd5a;
    11'b00010011111: data <= 32'hbe9db8e5;
    11'b00010100000: data <= 32'hbc05b901;
    11'b00010100001: data <= 32'h3ab2b718;
    11'b00010100010: data <= 32'h3df63870;
    11'b00010100011: data <= 32'hb09f3da7;
    11'b00010100100: data <= 32'hc0353cf4;
    11'b00010100101: data <= 32'hc01339c8;
    11'b00010100110: data <= 32'hb6193a97;
    11'b00010100111: data <= 32'h39313b9e;
    11'b00010101000: data <= 32'h366d27a7;
    11'b00010101001: data <= 32'h34d2bce0;
    11'b00010101010: data <= 32'h3ca3bb2e;
    11'b00010101011: data <= 32'h3f773c27;
    11'b00010101100: data <= 32'h3d784063;
    11'b00010101101: data <= 32'h35b83bc1;
    11'b00010101110: data <= 32'ha92abc90;
    11'b00010101111: data <= 32'hae62beea;
    11'b00010110000: data <= 32'hb8e5bab6;
    11'b00010110001: data <= 32'hbc1ab793;
    11'b00010110010: data <= 32'hb1fdbd26;
    11'b00010110011: data <= 32'h3d3bbee8;
    11'b00010110100: data <= 32'h3d79b976;
    11'b00010110101: data <= 32'hb8583a36;
    11'b00010110110: data <= 32'hc0903cb3;
    11'b00010110111: data <= 32'hbfad39f1;
    11'b00010111000: data <= 32'hb7103830;
    11'b00010111001: data <= 32'had823701;
    11'b00010111010: data <= 32'hbb73b2f3;
    11'b00010111011: data <= 32'hbbcfbb0e;
    11'b00010111100: data <= 32'h388ab209;
    11'b00010111101: data <= 32'h40033e69;
    11'b00010111110: data <= 32'h3ef540c3;
    11'b00010111111: data <= 32'h37753c75;
    11'b00011000000: data <= 32'hb265b81f;
    11'b00011000001: data <= 32'hae8bb87a;
    11'b00011000010: data <= 32'haebe34d9;
    11'b00011000011: data <= 32'hb063a9f8;
    11'b00011000100: data <= 32'h38bfbee1;
    11'b00011000101: data <= 32'h3e9ac107;
    11'b00011000110: data <= 32'h3de2bcdd;
    11'b00011000111: data <= 32'hb1d238ff;
    11'b00011001000: data <= 32'hbdd93c15;
    11'b00011001001: data <= 32'hbc4531f4;
    11'b00011001010: data <= 32'hb3c0b622;
    11'b00011001011: data <= 32'hba55b5cc;
    11'b00011001100: data <= 32'hc02db83f;
    11'b00011001101: data <= 32'hbf80ba7b;
    11'b00011001110: data <= 32'h329fb23b;
    11'b00011001111: data <= 32'h3f693ce7;
    11'b00011010000: data <= 32'h3d413f9a;
    11'b00011010001: data <= 32'hb4943c98;
    11'b00011010010: data <= 32'hbade35d6;
    11'b00011010011: data <= 32'hb3d03a82;
    11'b00011010100: data <= 32'h33873db3;
    11'b00011010101: data <= 32'h33a8364c;
    11'b00011010110: data <= 32'h3920bee2;
    11'b00011010111: data <= 32'h3e08c0cf;
    11'b00011011000: data <= 32'h3eafba43;
    11'b00011011001: data <= 32'h39db3c27;
    11'b00011011010: data <= 32'had143b8b;
    11'b00011011011: data <= 32'h2ce6b6e7;
    11'b00011011100: data <= 32'h3051bc68;
    11'b00011011101: data <= 32'hbc39b9e9;
    11'b00011011110: data <= 32'hc0d2b8c7;
    11'b00011011111: data <= 32'hbf7ebc29;
    11'b00011100000: data <= 32'h3548bbe3;
    11'b00011100001: data <= 32'h3e682638;
    11'b00011100010: data <= 32'h382e3b6c;
    11'b00011100011: data <= 32'hbce93bb7;
    11'b00011100100: data <= 32'hbdb53b80;
    11'b00011100101: data <= 32'hb5ad3e4c;
    11'b00011100110: data <= 32'h30d63f71;
    11'b00011100111: data <= 32'hb45c3850;
    11'b00011101000: data <= 32'hb3d0bd9b;
    11'b00011101001: data <= 32'h3a94be7d;
    11'b00011101010: data <= 32'h3f00320c;
    11'b00011101011: data <= 32'h3e643e91;
    11'b00011101100: data <= 32'h3c1f3baf;
    11'b00011101101: data <= 32'h3ab9b911;
    11'b00011101110: data <= 32'h372bbbf4;
    11'b00011101111: data <= 32'hba61b3bd;
    11'b00011110000: data <= 32'hbf50b2bc;
    11'b00011110001: data <= 32'hbc57bd63;
    11'b00011110010: data <= 32'h3a78c01e;
    11'b00011110011: data <= 32'h3dc7bd2a;
    11'b00011110100: data <= 32'ha165225a;
    11'b00011110101: data <= 32'hbe40392e;
    11'b00011110110: data <= 32'hbd4b3b05;
    11'b00011110111: data <= 32'hb25a3d58;
    11'b00011111000: data <= 32'hb3f33daa;
    11'b00011111001: data <= 32'hbd9234ec;
    11'b00011111010: data <= 32'hbe62bc2e;
    11'b00011111011: data <= 32'hac4aba87;
    11'b00011111100: data <= 32'h3e633b1d;
    11'b00011111101: data <= 32'h3f733f6f;
    11'b00011111110: data <= 32'h3cdc3b69;
    11'b00011111111: data <= 32'h3a60b50c;
    11'b00100000000: data <= 32'h37f2a85d;
    11'b00100000001: data <= 32'hb46c3bbd;
    11'b00100000010: data <= 32'hbb01382f;
    11'b00100000011: data <= 32'hb225bdd1;
    11'b00100000100: data <= 32'h3cc5c16e;
    11'b00100000101: data <= 32'h3d9fbfa6;
    11'b00100000110: data <= 32'h2cdbb4d7;
    11'b00100000111: data <= 32'hbb92365c;
    11'b00100001000: data <= 32'hb6a534d1;
    11'b00100001001: data <= 32'h34e13656;
    11'b00100001010: data <= 32'hb8e83843;
    11'b00100001011: data <= 32'hc0cdaaca;
    11'b00100001100: data <= 32'hc130baf2;
    11'b00100001101: data <= 32'hb916b8a7;
    11'b00100001110: data <= 32'h3d3039ac;
    11'b00100001111: data <= 32'h3d9c3d59;
    11'b00100010000: data <= 32'h3753395a;
    11'b00100010001: data <= 32'h2dde3301;
    11'b00100010010: data <= 32'h35013cb8;
    11'b00100010011: data <= 32'h30624065;
    11'b00100010100: data <= 32'hb4b73cd9;
    11'b00100010101: data <= 32'h29d7bd0e;
    11'b00100010110: data <= 32'h3c22c11b;
    11'b00100010111: data <= 32'h3d5cbe00;
    11'b00100011000: data <= 32'h392f2f61;
    11'b00100011001: data <= 32'h344d357e;
    11'b00100011010: data <= 32'h3ac1b5df;
    11'b00100011011: data <= 32'h3bb7b7df;
    11'b00100011100: data <= 32'hb925a61c;
    11'b00100011101: data <= 32'hc14fb01a;
    11'b00100011110: data <= 32'hc146baee;
    11'b00100011111: data <= 32'hb872bc2d;
    11'b00100100000: data <= 32'h3c2ab513;
    11'b00100100001: data <= 32'h38933403;
    11'b00100100010: data <= 32'hb8f631b9;
    11'b00100100011: data <= 32'hb923382a;
    11'b00100100100: data <= 32'h31803f6f;
    11'b00100100101: data <= 32'h33e64169;
    11'b00100100110: data <= 32'hb7f83dce;
    11'b00100100111: data <= 32'hb941bb38;
    11'b00100101000: data <= 32'h33d7bef0;
    11'b00100101001: data <= 32'h3c68b6bf;
    11'b00100101010: data <= 32'h3cdc3ae9;
    11'b00100101011: data <= 32'h3d23367b;
    11'b00100101100: data <= 32'h3ed6b9d0;
    11'b00100101101: data <= 32'h3db4b958;
    11'b00100101110: data <= 32'hb4d4348d;
    11'b00100101111: data <= 32'hc0123575;
    11'b00100110000: data <= 32'hbf18bae0;
    11'b00100110001: data <= 32'h2926bf35;
    11'b00100110010: data <= 32'h3b76be1b;
    11'b00100110011: data <= 32'hadb2ba4e;
    11'b00100110100: data <= 32'hbcdcb56e;
    11'b00100110101: data <= 32'hb9db3557;
    11'b00100110110: data <= 32'h36283e51;
    11'b00100110111: data <= 32'h30934071;
    11'b00100111000: data <= 32'hbd2f3c8e;
    11'b00100111001: data <= 32'hbf90b8b6;
    11'b00100111010: data <= 32'hba43ba98;
    11'b00100111011: data <= 32'h399b381e;
    11'b00100111100: data <= 32'h3d3c3d1b;
    11'b00100111101: data <= 32'h3db23577;
    11'b00100111110: data <= 32'h3ea8b971;
    11'b00100111111: data <= 32'h3dc2a748;
    11'b00101000000: data <= 32'h32293d75;
    11'b00101000001: data <= 32'hbbfb3cde;
    11'b00101000010: data <= 32'hb95ab97f;
    11'b00101000011: data <= 32'h38f8c07e;
    11'b00101000100: data <= 32'h3b1fc032;
    11'b00101000101: data <= 32'hb3e1bc91;
    11'b00101000110: data <= 32'hbb4eb8e2;
    11'b00101000111: data <= 32'h287eb3c6;
    11'b00101001000: data <= 32'h3c1b388d;
    11'b00101001001: data <= 32'h2cfd3c9f;
    11'b00101001010: data <= 32'hc02138b3;
    11'b00101001011: data <= 32'hc1aab6ed;
    11'b00101001100: data <= 32'hbdb7b5ff;
    11'b00101001101: data <= 32'h35253924;
    11'b00101001110: data <= 32'h3a813b4d;
    11'b00101001111: data <= 32'h38daa937;
    11'b00101010000: data <= 32'h3a7ab743;
    11'b00101010001: data <= 32'h3c553b64;
    11'b00101010010: data <= 32'h388f4112;
    11'b00101010011: data <= 32'hb3554008;
    11'b00101010100: data <= 32'hb031b5c4;
    11'b00101010101: data <= 32'h3919c006;
    11'b00101010110: data <= 32'h39c7be87;
    11'b00101010111: data <= 32'h2512b8eb;
    11'b00101011000: data <= 32'h266cb82f;
    11'b00101011001: data <= 32'h3cebbaf7;
    11'b00101011010: data <= 32'h3f4bb7b2;
    11'b00101011011: data <= 32'h338034f6;
    11'b00101011100: data <= 32'hc06a3517;
    11'b00101011101: data <= 32'hc1a8b5b7;
    11'b00101011110: data <= 32'hbd21b854;
    11'b00101011111: data <= 32'h3145adfc;
    11'b00101100000: data <= 32'h2341ae5e;
    11'b00101100001: data <= 32'hb8e5b97e;
    11'b00101100010: data <= 32'hb244b615;
    11'b00101100011: data <= 32'h39e23dd6;
    11'b00101100100: data <= 32'h39c64203;
    11'b00101100101: data <= 32'hb0e74079;
    11'b00101100110: data <= 32'hb843aa42;
    11'b00101100111: data <= 32'hab80bcd3;
    11'b00101101000: data <= 32'h3527b6e1;
    11'b00101101001: data <= 32'h35373620;
    11'b00101101010: data <= 32'h3af4b406;
    11'b00101101011: data <= 32'h4021bcfc;
    11'b00101101100: data <= 32'h40a0bb53;
    11'b00101101101: data <= 32'h38a434f7;
    11'b00101101110: data <= 32'hbe4f395f;
    11'b00101101111: data <= 32'hbf6fb247;
    11'b00101110000: data <= 32'hb771bc10;
    11'b00101110001: data <= 32'h3420bc6b;
    11'b00101110010: data <= 32'hb927bc77;
    11'b00101110011: data <= 32'hbdc8bd1f;
    11'b00101110100: data <= 32'hb8c9b905;
    11'b00101110101: data <= 32'h3a733c96;
    11'b00101110110: data <= 32'h3a0840dd;
    11'b00101110111: data <= 32'hb9453ef4;
    11'b00101111000: data <= 32'hbe2f2d3f;
    11'b00101111001: data <= 32'hbc41b4eb;
    11'b00101111010: data <= 32'hb23a39d3;
    11'b00101111011: data <= 32'h34dd3c71;
    11'b00101111100: data <= 32'h3b99b0be;
    11'b00101111101: data <= 32'h3fd0bd3f;
    11'b00101111110: data <= 32'h4060b88d;
    11'b00101111111: data <= 32'h3b5f3c98;
    11'b00110000000: data <= 32'hb86e3e11;
    11'b00110000001: data <= 32'hb8632fad;
    11'b00110000010: data <= 32'h36debd31;
    11'b00110000011: data <= 32'h3676be5d;
    11'b00110000100: data <= 32'hbb1cbdb2;
    11'b00110000101: data <= 32'hbdbbbddc;
    11'b00110000110: data <= 32'haddabc5f;
    11'b00110000111: data <= 32'h3d9c30aa;
    11'b00110001000: data <= 32'h3ac73cb7;
    11'b00110001001: data <= 32'hbce73b0e;
    11'b00110001010: data <= 32'hc0c12853;
    11'b00110001011: data <= 32'hbebc3298;
    11'b00110001100: data <= 32'hb8583c90;
    11'b00110001101: data <= 32'hb0283c1b;
    11'b00110001110: data <= 32'h3034b76a;
    11'b00110001111: data <= 32'h3b7abcfc;
    11'b00110010000: data <= 32'h3e2f30ed;
    11'b00110010001: data <= 32'h3c5a4060;
    11'b00110010010: data <= 32'h3420409c;
    11'b00110010011: data <= 32'h34513780;
    11'b00110010100: data <= 32'h39f9bc48;
    11'b00110010101: data <= 32'h354abc70;
    11'b00110010110: data <= 32'hba39ba14;
    11'b00110010111: data <= 32'hb9f5bc81;
    11'b00110011000: data <= 32'h3b99be12;
    11'b00110011001: data <= 32'h4066bb75;
    11'b00110011010: data <= 32'h3c492bbe;
    11'b00110011011: data <= 32'hbd4e34ae;
    11'b00110011100: data <= 32'hc0b0a43d;
    11'b00110011101: data <= 32'hbdb731d8;
    11'b00110011110: data <= 32'hb7df3960;
    11'b00110011111: data <= 32'hb9fa321f;
    11'b00110100000: data <= 32'hbc6dbc72;
    11'b00110100001: data <= 32'hb551bd1c;
    11'b00110100010: data <= 32'h3aed38d3;
    11'b00110100011: data <= 32'h3c56413a;
    11'b00110100100: data <= 32'h375740e5;
    11'b00110100101: data <= 32'h30c138fb;
    11'b00110100110: data <= 32'h3416b6a4;
    11'b00110100111: data <= 32'hac2d2f07;
    11'b00110101000: data <= 32'hb8d637bd;
    11'b00110101001: data <= 32'ha6b8b829;
    11'b00110101010: data <= 32'h3eeabeda;
    11'b00110101011: data <= 32'h4149bde4;
    11'b00110101100: data <= 32'h3d41b35c;
    11'b00110101101: data <= 32'hba79368a;
    11'b00110101110: data <= 32'hbd692fbe;
    11'b00110101111: data <= 32'hb62ab096;
    11'b00110110000: data <= 32'hacc6b1bb;
    11'b00110110001: data <= 32'hbcdaba09;
    11'b00110110010: data <= 32'hc00fbec1;
    11'b00110110011: data <= 32'hbc21bde8;
    11'b00110110100: data <= 32'h395635ca;
    11'b00110110101: data <= 32'h3c424009;
    11'b00110110110: data <= 32'h2edf3eff;
    11'b00110110111: data <= 32'hb9613737;
    11'b00110111000: data <= 32'hb94834a3;
    11'b00110111001: data <= 32'hb8b23d61;
    11'b00110111010: data <= 32'hb90b3e0e;
    11'b00110111011: data <= 32'h2d63af94;
    11'b00110111100: data <= 32'h3e61bec7;
    11'b00110111101: data <= 32'h40b3bd1b;
    11'b00110111110: data <= 32'h3d8a363c;
    11'b00110111111: data <= 32'h279c3c8f;
    11'b00111000000: data <= 32'h26fb3742;
    11'b00111000001: data <= 32'h3a80b600;
    11'b00111000010: data <= 32'h364bb93a;
    11'b00111000011: data <= 32'hbd61bc2c;
    11'b00111000100: data <= 32'hc052befd;
    11'b00111000101: data <= 32'hba25bedd;
    11'b00111000110: data <= 32'h3c79b789;
    11'b00111000111: data <= 32'h3cb1399d;
    11'b00111001000: data <= 32'hb5fc38bf;
    11'b00111001001: data <= 32'hbdd12c22;
    11'b00111001010: data <= 32'hbd083954;
    11'b00111001011: data <= 32'hbacf3f95;
    11'b00111001100: data <= 32'hbb213ec8;
    11'b00111001101: data <= 32'hb8b8b411;
    11'b00111001110: data <= 32'h382fbe88;
    11'b00111001111: data <= 32'h3db1b94c;
    11'b00111010000: data <= 32'h3cd53d60;
    11'b00111010001: data <= 32'h397c3f99;
    11'b00111010010: data <= 32'h3bd23a0b;
    11'b00111010011: data <= 32'h3daeb444;
    11'b00111010100: data <= 32'h384bb495;
    11'b00111010101: data <= 32'hbce0b559;
    11'b00111010110: data <= 32'hbe63bc97;
    11'b00111010111: data <= 32'h30fcbf3a;
    11'b00111011000: data <= 32'h3f80bd87;
    11'b00111011001: data <= 32'h3d84b858;
    11'b00111011010: data <= 32'hb858b4f1;
    11'b00111011011: data <= 32'hbe02b3be;
    11'b00111011100: data <= 32'hbbc038d4;
    11'b00111011101: data <= 32'hb89b3e40;
    11'b00111011110: data <= 32'hbccb3c0a;
    11'b00111011111: data <= 32'hbea3bac5;
    11'b00111100000: data <= 32'hbae8beac;
    11'b00111100001: data <= 32'h36a2b216;
    11'b00111100010: data <= 32'h3b4a3f48;
    11'b00111100011: data <= 32'h3a914009;
    11'b00111100100: data <= 32'h3c0239ce;
    11'b00111100101: data <= 32'h3c762f60;
    11'b00111100110: data <= 32'h33273a2d;
    11'b00111100111: data <= 32'hbc3d3c14;
    11'b00111101000: data <= 32'hbb27b2b7;
    11'b00111101001: data <= 32'h3ba9beb9;
    11'b00111101010: data <= 32'h409cbf52;
    11'b00111101011: data <= 32'h3decbbe3;
    11'b00111101100: data <= 32'hb41db6ac;
    11'b00111101101: data <= 32'hb945b31f;
    11'b00111101110: data <= 32'h319b34b1;
    11'b00111101111: data <= 32'h315c3a16;
    11'b00111110000: data <= 32'hbd512c7b;
    11'b00111110001: data <= 32'hc0f0bdac;
    11'b00111110010: data <= 32'hbee1bf13;
    11'b00111110011: data <= 32'ha9dfb3cc;
    11'b00111110100: data <= 32'h39d93d6d;
    11'b00111110101: data <= 32'h37993ced;
    11'b00111110110: data <= 32'h342433d9;
    11'b00111110111: data <= 32'h339d37c1;
    11'b00111111000: data <= 32'hb4b73f88;
    11'b00111111001: data <= 32'hbc1c406b;
    11'b00111111010: data <= 32'hb91f37cb;
    11'b00111111011: data <= 32'h3b88bdd6;
    11'b00111111100: data <= 32'h3fc6be7d;
    11'b00111111101: data <= 32'h3d15b778;
    11'b00111111110: data <= 32'h341c339a;
    11'b00111111111: data <= 32'h38bc2e2c;
    11'b01000000000: data <= 32'h3e24285d;
    11'b01000000001: data <= 32'h3ba931fb;
    11'b01000000010: data <= 32'hbcdeb51b;
    11'b01000000011: data <= 32'hc123bdb9;
    11'b01000000100: data <= 32'hbe4ebf0e;
    11'b01000000101: data <= 32'h3498ba2d;
    11'b01000000110: data <= 32'h3a6d317c;
    11'b01000000111: data <= 32'ha34bad70;
    11'b01000001000: data <= 32'hb8a8b7b7;
    11'b01000001001: data <= 32'hb71238ac;
    11'b01000001010: data <= 32'hb84b40c5;
    11'b01000001011: data <= 32'hbc5a4110;
    11'b01000001100: data <= 32'hbc27381a;
    11'b01000001101: data <= 32'h055abd52;
    11'b01000001110: data <= 32'h3aeabc08;
    11'b01000001111: data <= 32'h39f63815;
    11'b01000010000: data <= 32'h38e53c3a;
    11'b01000010001: data <= 32'h3deb364f;
    11'b01000010010: data <= 32'h409ba225;
    11'b01000010011: data <= 32'h3d3b34ff;
    11'b01000010100: data <= 32'hbbe53426;
    11'b01000010101: data <= 32'hc003b993;
    11'b01000010110: data <= 32'hb94abe0b;
    11'b01000010111: data <= 32'h3c4ebd78;
    11'b01000011000: data <= 32'h3c0fbc00;
    11'b01000011001: data <= 32'hb4bfbcaa;
    11'b01000011010: data <= 32'hbaadbc2b;
    11'b01000011011: data <= 32'hb47b3608;
    11'b01000011100: data <= 32'hb0d74019;
    11'b01000011101: data <= 32'hbc493f8b;
    11'b01000011110: data <= 32'hbf29ad06;
    11'b01000011111: data <= 32'hbd37bd7a;
    11'b01000100000: data <= 32'hb562b74a;
    11'b01000100001: data <= 32'h30e13c9f;
    11'b01000100010: data <= 32'h387d3d30;
    11'b01000100011: data <= 32'h3dfc3485;
    11'b01000100100: data <= 32'h40242d02;
    11'b01000100101: data <= 32'h3c243c3f;
    11'b01000100110: data <= 32'hba943e18;
    11'b01000100111: data <= 32'hbcfe3704;
    11'b01000101000: data <= 32'h3471bc3b;
    11'b01000101001: data <= 32'h3e7dbe5e;
    11'b01000101010: data <= 32'h3c40bdb5;
    11'b01000101011: data <= 32'hb43fbd87;
    11'b01000101100: data <= 32'hb488bc72;
    11'b01000101101: data <= 32'h3a232928;
    11'b01000101110: data <= 32'h3a473cd7;
    11'b01000101111: data <= 32'hbada3aba;
    11'b01000110000: data <= 32'hc0b1ba11;
    11'b01000110001: data <= 32'hc046bdc4;
    11'b01000110010: data <= 32'hbb84b4af;
    11'b01000110011: data <= 32'hb1773bb8;
    11'b01000110100: data <= 32'h311038eb;
    11'b01000110101: data <= 32'h39d6b60b;
    11'b01000110110: data <= 32'h3c7e2e3d;
    11'b01000110111: data <= 32'h36cd3f99;
    11'b01000111000: data <= 32'hba42415e;
    11'b01000111001: data <= 32'hba853d3b;
    11'b01000111010: data <= 32'h381ab91a;
    11'b01000111011: data <= 32'h3d7fbd28;
    11'b01000111100: data <= 32'h398dbb26;
    11'b01000111101: data <= 32'hae01b993;
    11'b01000111110: data <= 32'h3979b9d1;
    11'b01000111111: data <= 32'h402fb2de;
    11'b01001000000: data <= 32'h3f1637e0;
    11'b01001000001: data <= 32'hb7fa3316;
    11'b01001000010: data <= 32'hc0a0bb28;
    11'b01001000011: data <= 32'hbfefbd39;
    11'b01001000100: data <= 32'hb8efb7ee;
    11'b01001000101: data <= 32'hac8e2c33;
    11'b01001000110: data <= 32'hb53eb94e;
    11'b01001000111: data <= 32'hb331bd47;
    11'b01001001000: data <= 32'h339eada8;
    11'b01001001001: data <= 32'h2a6d4078;
    11'b01001001010: data <= 32'hb9f741ff;
    11'b01001001011: data <= 32'hbb4e3d8c;
    11'b01001001100: data <= 32'hb08db7d4;
    11'b01001001101: data <= 32'h357bb953;
    11'b01001001110: data <= 32'haaee3185;
    11'b01001001111: data <= 32'haaf234cb;
    11'b01001010000: data <= 32'h3d84b4b4;
    11'b01001010001: data <= 32'h41b9b532;
    11'b01001010010: data <= 32'h40703593;
    11'b01001010011: data <= 32'hb24d3823;
    11'b01001010100: data <= 32'hbee0b32f;
    11'b01001010101: data <= 32'hbbfbbaaf;
    11'b01001010110: data <= 32'h3514ba0e;
    11'b01001010111: data <= 32'h344bbb20;
    11'b01001011000: data <= 32'hb92fbf01;
    11'b01001011001: data <= 32'hb9b5c00a;
    11'b01001011010: data <= 32'h2ff2b6bc;
    11'b01001011011: data <= 32'h35a23f5e;
    11'b01001011100: data <= 32'hb83d4099;
    11'b01001011101: data <= 32'hbd4b397e;
    11'b01001011110: data <= 32'hbcd9b91b;
    11'b01001011111: data <= 32'hbaf2add8;
    11'b01001100000: data <= 32'hba9f3c19;
    11'b01001100001: data <= 32'hb48a3a72;
    11'b01001100010: data <= 32'h3d3fb4d5;
    11'b01001100011: data <= 32'h4130b683;
    11'b01001100100: data <= 32'h3f853a1a;
    11'b01001100101: data <= 32'haf553e22;
    11'b01001100110: data <= 32'hbb8f3b58;
    11'b01001100111: data <= 32'h2fd3b17c;
    11'b01001101000: data <= 32'h3c79ba07;
    11'b01001101001: data <= 32'h36ffbcd4;
    11'b01001101010: data <= 32'hba11bfcf;
    11'b01001101011: data <= 32'hb7bac025;
    11'b01001101100: data <= 32'h3b51b9b5;
    11'b01001101101: data <= 32'h3d243be6;
    11'b01001101110: data <= 32'had8d3c64;
    11'b01001101111: data <= 32'hbe73b36f;
    11'b01001110000: data <= 32'hbfa4bac3;
    11'b01001110001: data <= 32'hbde731e1;
    11'b01001110010: data <= 32'hbcc13c8c;
    11'b01001110011: data <= 32'hb9853635;
    11'b01001110100: data <= 32'h382cbb8b;
    11'b01001110101: data <= 32'h3e0eb8f4;
    11'b01001110110: data <= 32'h3c353d3a;
    11'b01001110111: data <= 32'hb2e44112;
    11'b01001111000: data <= 32'hb6d23f3c;
    11'b01001111001: data <= 32'h3923356f;
    11'b01001111010: data <= 32'h3c90b650;
    11'b01001111011: data <= 32'h2eecb917;
    11'b01001111100: data <= 32'hba7cbca5;
    11'b01001111101: data <= 32'h319fbe03;
    11'b01001111110: data <= 32'h4021baa8;
    11'b01001111111: data <= 32'h409c3292;
    11'b01010000000: data <= 32'h369332c4;
    11'b01010000001: data <= 32'hbde1b92e;
    11'b01010000010: data <= 32'hbecfba33;
    11'b01010000011: data <= 32'hbc4e3208;
    11'b01010000100: data <= 32'hbb94386e;
    11'b01010000101: data <= 32'hbc3ab999;
    11'b01010000110: data <= 32'hb7b4bfb2;
    11'b01010000111: data <= 32'h361bbbde;
    11'b01010001000: data <= 32'h364b3df0;
    11'b01010001001: data <= 32'hb455418f;
    11'b01010001010: data <= 32'hb56b3f5c;
    11'b01010001011: data <= 32'h34e73661;
    11'b01010001100: data <= 32'h35113088;
    11'b01010001101: data <= 32'hb96c3789;
    11'b01010001110: data <= 32'hbbd32b8e;
    11'b01010001111: data <= 32'h3962ba50;
    11'b01010010000: data <= 32'h417eba9a;
    11'b01010010001: data <= 32'h4178ae45;
    11'b01010010010: data <= 32'h396d320a;
    11'b01010010011: data <= 32'hbb61b28f;
    11'b01010010100: data <= 32'hb965b472;
    11'b01010010101: data <= 32'h2b3830df;
    11'b01010010110: data <= 32'hb573b17b;
    11'b01010010111: data <= 32'hbcfbbec0;
    11'b01010011000: data <= 32'hbc6ac146;
    11'b01010011001: data <= 32'ha9e4bd5a;
    11'b01010011010: data <= 32'h37233c61;
    11'b01010011011: data <= 32'haa794012;
    11'b01010011100: data <= 32'hb8273bbf;
    11'b01010011101: data <= 32'hb80c1f16;
    11'b01010011110: data <= 32'hba4038a5;
    11'b01010011111: data <= 32'hbdf53dbf;
    11'b01010100000: data <= 32'hbd233af8;
    11'b01010100001: data <= 32'h3884b838;
    11'b01010100010: data <= 32'h40dcbb11;
    11'b01010100011: data <= 32'h40832de8;
    11'b01010100100: data <= 32'h386c3b6a;
    11'b01010100101: data <= 32'hb4693a75;
    11'b01010100110: data <= 32'h38593714;
    11'b01010100111: data <= 32'h3c9d3483;
    11'b01010101000: data <= 32'h2f3db678;
    11'b01010101001: data <= 32'hbd35bf5b;
    11'b01010101010: data <= 32'hbc55c12d;
    11'b01010101011: data <= 32'h3735bdde;
    11'b01010101100: data <= 32'h3ce83595;
    11'b01010101101: data <= 32'h374539f4;
    11'b01010101110: data <= 32'hb921b383;
    11'b01010101111: data <= 32'hbc50b7e8;
    11'b01010110000: data <= 32'hbd593a35;
    11'b01010110001: data <= 32'hbf2b3ef7;
    11'b01010110010: data <= 32'hbe523a10;
    11'b01010110011: data <= 32'hb093bbee;
    11'b01010110100: data <= 32'h3d15bc9a;
    11'b01010110101: data <= 32'h3ca53717;
    11'b01010110110: data <= 32'h31053f12;
    11'b01010110111: data <= 32'h30973e90;
    11'b01010111000: data <= 32'h3cf83b80;
    11'b01010111001: data <= 32'h3df738b8;
    11'b01010111010: data <= 32'ha1812f73;
    11'b01010111011: data <= 32'hbd92bbd2;
    11'b01010111100: data <= 32'hb90fbf1d;
    11'b01010111101: data <= 32'h3da4bd34;
    11'b01010111110: data <= 32'h405cb523;
    11'b01010111111: data <= 32'h3bc5b4ec;
    11'b01011000000: data <= 32'hb7ddbbcc;
    11'b01011000001: data <= 32'hbb13b943;
    11'b01011000010: data <= 32'hbb023a62;
    11'b01011000011: data <= 32'hbd643d7e;
    11'b01011000100: data <= 32'hbec0af32;
    11'b01011000101: data <= 32'hbc1fbf94;
    11'b01011000110: data <= 32'ha3d8be3d;
    11'b01011000111: data <= 32'h317d387f;
    11'b01011001000: data <= 32'hb12d3ff4;
    11'b01011001001: data <= 32'h331f3e7a;
    11'b01011001010: data <= 32'h3c7e3ab0;
    11'b01011001011: data <= 32'h3b453b3d;
    11'b01011001100: data <= 32'hb99e3c76;
    11'b01011001101: data <= 32'hbe7c3622;
    11'b01011001110: data <= 32'hb394b9df;
    11'b01011001111: data <= 32'h4012bc07;
    11'b01011010000: data <= 32'h4122b8b6;
    11'b01011010001: data <= 32'h3c7fb85d;
    11'b01011010010: data <= 32'haf85ba67;
    11'b01011010011: data <= 32'h2a7fb47c;
    11'b01011010100: data <= 32'h36273aa2;
    11'b01011010101: data <= 32'hb6be3a45;
    11'b01011010110: data <= 32'hbe4ebc0f;
    11'b01011010111: data <= 32'hbe60c124;
    11'b01011011000: data <= 32'hb93cbf63;
    11'b01011011001: data <= 32'hac8f34b3;
    11'b01011011010: data <= 32'hae013d42;
    11'b01011011011: data <= 32'h2eb33912;
    11'b01011011100: data <= 32'h379630af;
    11'b01011011101: data <= 32'hacc23c2e;
    11'b01011011110: data <= 32'hbdee4002;
    11'b01011011111: data <= 32'hbf9d3d9b;
    11'b01011100000: data <= 32'hb468b0e6;
    11'b01011100001: data <= 32'h3f11bb01;
    11'b01011100010: data <= 32'h3ff6b722;
    11'b01011100011: data <= 32'h39d92004;
    11'b01011100100: data <= 32'h33db2c31;
    11'b01011100101: data <= 32'h3cbe3682;
    11'b01011100110: data <= 32'h3eba3bc8;
    11'b01011100111: data <= 32'h35ed383e;
    11'b01011101000: data <= 32'hbda0bcc5;
    11'b01011101001: data <= 32'hbe65c0e3;
    11'b01011101010: data <= 32'hb5b4befd;
    11'b01011101011: data <= 32'h383bb232;
    11'b01011101100: data <= 32'h35d52ec4;
    11'b01011101101: data <= 32'h2635ba1b;
    11'b01011101110: data <= 32'haca5b9a2;
    11'b01011101111: data <= 32'hb9143be2;
    11'b01011110000: data <= 32'hbeec40a0;
    11'b01011110001: data <= 32'hc0093dfd;
    11'b01011110010: data <= 32'hba11b66c;
    11'b01011110011: data <= 32'h397abc4a;
    11'b01011110100: data <= 32'h39afb0dc;
    11'b01011110101: data <= 32'ha4553a42;
    11'b01011110110: data <= 32'h36373b0a;
    11'b01011110111: data <= 32'h3f7c3af2;
    11'b01011111000: data <= 32'h407a3c9a;
    11'b01011111001: data <= 32'h37f43af2;
    11'b01011111010: data <= 32'hbd95b671;
    11'b01011111011: data <= 32'hbcd4bddd;
    11'b01011111100: data <= 32'h3805bcf2;
    11'b01011111101: data <= 32'h3dc0b89c;
    11'b01011111110: data <= 32'h3ae5bb5b;
    11'b01011111111: data <= 32'h2e0dbeee;
    11'b01100000000: data <= 32'ha3f1bc9d;
    11'b01100000001: data <= 32'hb39a3af7;
    11'b01100000010: data <= 32'hbc904000;
    11'b01100000011: data <= 32'hbf373a0a;
    11'b01100000100: data <= 32'hbd6fbceb;
    11'b01100000101: data <= 32'hb884bdde;
    11'b01100000110: data <= 32'hb8221c00;
    11'b01100000111: data <= 32'hb93e3c61;
    11'b01100001000: data <= 32'h34b63b4d;
    11'b01100001001: data <= 32'h3f323934;
    11'b01100001010: data <= 32'h3f3d3cb8;
    11'b01100001011: data <= 32'had913e5e;
    11'b01100001100: data <= 32'hbe6d3b52;
    11'b01100001101: data <= 32'hba75b1d4;
    11'b01100001110: data <= 32'h3cb6b8c4;
    11'b01100001111: data <= 32'h3f76b917;
    11'b01100010000: data <= 32'h3b6ebcc7;
    11'b01100010001: data <= 32'h3345bef4;
    11'b01100010010: data <= 32'h3959bb60;
    11'b01100010011: data <= 32'h3bce3af5;
    11'b01100010100: data <= 32'h24c33db8;
    11'b01100010101: data <= 32'hbd51b12a;
    11'b01100010110: data <= 32'hbebcbfbf;
    11'b01100010111: data <= 32'hbcebbec8;
    11'b01100011000: data <= 32'hbbbcac7d;
    11'b01100011001: data <= 32'hba383922;
    11'b01100011010: data <= 32'h2fc4a631;
    11'b01100011011: data <= 32'h3cbdb420;
    11'b01100011100: data <= 32'h3ac73ba6;
    11'b01100011101: data <= 32'hbb0f4073;
    11'b01100011110: data <= 32'hbf6b3fcc;
    11'b01100011111: data <= 32'hb996390b;
    11'b01100100000: data <= 32'h3c65b341;
    11'b01100100001: data <= 32'h3d5cb67e;
    11'b01100100010: data <= 32'h356cb97d;
    11'b01100100011: data <= 32'h33a2bb6f;
    11'b01100100100: data <= 32'h3e28b3b8;
    11'b01100100101: data <= 32'h40903bfc;
    11'b01100100110: data <= 32'h3c3e3c4a;
    11'b01100100111: data <= 32'hbb06b7f1;
    11'b01100101000: data <= 32'hbe43bf75;
    11'b01100101001: data <= 32'hbbd9bdb6;
    11'b01100101010: data <= 32'hb760b35c;
    11'b01100101011: data <= 32'hb5b6b4e6;
    11'b01100101100: data <= 32'h2841bdb3;
    11'b01100101101: data <= 32'h3895bd7c;
    11'b01100101110: data <= 32'h312b389f;
    11'b01100101111: data <= 32'hbcc240c0;
    11'b01100110000: data <= 32'hbf584030;
    11'b01100110001: data <= 32'hbb16381d;
    11'b01100110010: data <= 32'h3448b584;
    11'b01100110011: data <= 32'h2bceae54;
    11'b01100110100: data <= 32'hb96b2fca;
    11'b01100110101: data <= 32'h28d0a5c0;
    11'b01100110110: data <= 32'h40133481;
    11'b01100110111: data <= 32'h41c63c51;
    11'b01100111000: data <= 32'h3d6d3c9d;
    11'b01100111001: data <= 32'hb9f02b30;
    11'b01100111010: data <= 32'hbc94bb29;
    11'b01100111011: data <= 32'haf33b93c;
    11'b01100111100: data <= 32'h380ab411;
    11'b01100111101: data <= 32'h324cbc7f;
    11'b01100111110: data <= 32'h2923c0e4;
    11'b01100111111: data <= 32'h36abc00d;
    11'b01101000000: data <= 32'h356534a0;
    11'b01101000001: data <= 32'hb8fb4004;
    11'b01101000010: data <= 32'hbd7f3d70;
    11'b01101000011: data <= 32'hbc80b55e;
    11'b01101000100: data <= 32'hba16ba40;
    11'b01101000101: data <= 32'hbce12e17;
    11'b01101000110: data <= 32'hbe3938d8;
    11'b01101000111: data <= 32'hb47532c5;
    11'b01101001000: data <= 32'h3f8a2e8c;
    11'b01101001001: data <= 32'h40f63b1e;
    11'b01101001010: data <= 32'h3a533e1c;
    11'b01101001011: data <= 32'hbbc23c93;
    11'b01101001100: data <= 32'hb9c23712;
    11'b01101001101: data <= 32'h39943414;
    11'b01101001110: data <= 32'h3c73a9f5;
    11'b01101001111: data <= 32'h3513bd2c;
    11'b01101010000: data <= 32'ha12cc0fb;
    11'b01101010001: data <= 32'h3a2ebf6c;
    11'b01101010010: data <= 32'h3d45345b;
    11'b01101010011: data <= 32'h38aa3dab;
    11'b01101010100: data <= 32'hb8e93570;
    11'b01101010101: data <= 32'hbc94bccb;
    11'b01101010110: data <= 32'hbd2ebc4c;
    11'b01101010111: data <= 32'hbee63158;
    11'b01101011000: data <= 32'hbf263737;
    11'b01101011001: data <= 32'hb812b7eb;
    11'b01101011010: data <= 32'h3cfdbab9;
    11'b01101011011: data <= 32'h3dc63608;
    11'b01101011100: data <= 32'hb0623f50;
    11'b01101011101: data <= 32'hbd28400d;
    11'b01101011110: data <= 32'hb7fa3d4b;
    11'b01101011111: data <= 32'h3b133a46;
    11'b01101100000: data <= 32'h3a7f34a5;
    11'b01101100001: data <= 32'hb4a6b9fe;
    11'b01101100010: data <= 32'hb46fbe87;
    11'b01101100011: data <= 32'h3d33bc4c;
    11'b01101100100: data <= 32'h40e83787;
    11'b01101100101: data <= 32'h3ed23bcf;
    11'b01101100110: data <= 32'h29a9b369;
    11'b01101100111: data <= 32'hbaf1bd63;
    11'b01101101000: data <= 32'hbbf4ba79;
    11'b01101101001: data <= 32'hbccb3440;
    11'b01101101010: data <= 32'hbd39b0ed;
    11'b01101101011: data <= 32'hb851bedc;
    11'b01101101100: data <= 32'h3898c014;
    11'b01101101101: data <= 32'h3866b3e3;
    11'b01101101110: data <= 32'hb9483f16;
    11'b01101101111: data <= 32'hbd2e4032;
    11'b01101110000: data <= 32'hb7473cdc;
    11'b01101110001: data <= 32'h3639393b;
    11'b01101110010: data <= 32'hb46e3885;
    11'b01101110011: data <= 32'hbd932eb1;
    11'b01101110100: data <= 32'hba01b863;
    11'b01101110101: data <= 32'h3e35b57f;
    11'b01101110110: data <= 32'h41f038cd;
    11'b01101110111: data <= 32'h40123add;
    11'b01101111000: data <= 32'h331597f1;
    11'b01101111001: data <= 32'hb711b89b;
    11'b01101111010: data <= 32'had6f29db;
    11'b01101111011: data <= 32'had80383e;
    11'b01101111100: data <= 32'hb87bb98e;
    11'b01101111101: data <= 32'hb773c143;
    11'b01101111110: data <= 32'h3409c183;
    11'b01101111111: data <= 32'h36b5b90c;
    11'b01110000000: data <= 32'hb4d33d6b;
    11'b01110000001: data <= 32'hba263d49;
    11'b01110000010: data <= 32'hb6693401;
    11'b01110000011: data <= 32'hb56e2a93;
    11'b01110000100: data <= 32'hbdc73978;
    11'b01110000101: data <= 32'hc0b739c8;
    11'b01110000110: data <= 32'hbcdda701;
    11'b01110000111: data <= 32'h3d37b4d9;
    11'b01110001000: data <= 32'h410835ec;
    11'b01110001001: data <= 32'h3d8c3b92;
    11'b01110001010: data <= 32'hb0613a2c;
    11'b01110001011: data <= 32'hada13918;
    11'b01110001100: data <= 32'h3aad3c3e;
    11'b01110001101: data <= 32'h3a4b3b7d;
    11'b01110001110: data <= 32'hb2c8b9cb;
    11'b01110001111: data <= 32'hb837c13f;
    11'b01110010000: data <= 32'h357ac113;
    11'b01110010001: data <= 32'h3c50b87c;
    11'b01110010010: data <= 32'h3a203a8d;
    11'b01110010011: data <= 32'h2ef132af;
    11'b01110010100: data <= 32'hb1d0bad9;
    11'b01110010101: data <= 32'hb98eb78f;
    11'b01110010110: data <= 32'hbf9239e8;
    11'b01110010111: data <= 32'hc1293a76;
    11'b01110011000: data <= 32'hbda4b698;
    11'b01110011001: data <= 32'h3990bc5c;
    11'b01110011010: data <= 32'h3d96b41d;
    11'b01110011011: data <= 32'h33a93bd5;
    11'b01110011100: data <= 32'hb9763dc0;
    11'b01110011101: data <= 32'h2e023dd5;
    11'b01110011110: data <= 32'h3cf13e7e;
    11'b01110011111: data <= 32'h3a6f3d2d;
    11'b01110100000: data <= 32'hb92bb1b7;
    11'b01110100001: data <= 32'hbb2abec6;
    11'b01110100010: data <= 32'h38b5be41;
    11'b01110100011: data <= 32'h3fe2b0be;
    11'b01110100100: data <= 32'h3f4936eb;
    11'b01110100101: data <= 32'h3ab3b86c;
    11'b01110100110: data <= 32'h31a6bd45;
    11'b01110100111: data <= 32'hb5adb665;
    11'b01110101000: data <= 32'hbd373b58;
    11'b01110101001: data <= 32'hbfc637c9;
    11'b01110101010: data <= 32'hbd00bd78;
    11'b01110101011: data <= 32'h2d5fc06e;
    11'b01110101100: data <= 32'h3557bbd9;
    11'b01110101101: data <= 32'hb8bc3a4a;
    11'b01110101110: data <= 32'hbb353dbc;
    11'b01110101111: data <= 32'h322d3d2d;
    11'b01110110000: data <= 32'h3c113d85;
    11'b01110110001: data <= 32'h9d9b3da9;
    11'b01110110010: data <= 32'hbea738ef;
    11'b01110110011: data <= 32'hbdf4b758;
    11'b01110110100: data <= 32'h3941b845;
    11'b01110110101: data <= 32'h40be32c5;
    11'b01110110110: data <= 32'h40353496;
    11'b01110110111: data <= 32'h3b99b8b9;
    11'b01110111000: data <= 32'h37f9bab7;
    11'b01110111001: data <= 32'h381435a8;
    11'b01110111010: data <= 32'hab763d3f;
    11'b01110111011: data <= 32'hbb513142;
    11'b01110111100: data <= 32'hbb7bc046;
    11'b01110111101: data <= 32'hb3a2c1c7;
    11'b01110111110: data <= 32'haa82bd65;
    11'b01110111111: data <= 32'hb85236b3;
    11'b01111000000: data <= 32'hb7f9396c;
    11'b01111000001: data <= 32'h35fd32d4;
    11'b01111000010: data <= 32'h38423827;
    11'b01111000011: data <= 32'hbc003d2d;
    11'b01111000100: data <= 32'hc12f3cda;
    11'b01111000101: data <= 32'hbfee34ce;
    11'b01111000110: data <= 32'h366eb18d;
    11'b01111000111: data <= 32'h3fa63048;
    11'b01111001000: data <= 32'h3d6a3429;
    11'b01111001001: data <= 32'h35ddacee;
    11'b01111001010: data <= 32'h3905319e;
    11'b01111001011: data <= 32'h3d943d57;
    11'b01111001100: data <= 32'h3c263f25;
    11'b01111001101: data <= 32'hb39e323a;
    11'b01111001110: data <= 32'hba82c032;
    11'b01111001111: data <= 32'hb3bec12c;
    11'b01111010000: data <= 32'h356cbc60;
    11'b01111010001: data <= 32'h34e02d0f;
    11'b01111010010: data <= 32'h3574b661;
    11'b01111010011: data <= 32'h3991bc66;
    11'b01111010100: data <= 32'h3496b55e;
    11'b01111010101: data <= 32'hbd913c8f;
    11'b01111010110: data <= 32'hc1813d77;
    11'b01111010111: data <= 32'hc01431ff;
    11'b01111011000: data <= 32'haa0db9b3;
    11'b01111011001: data <= 32'h3a96b70d;
    11'b01111011010: data <= 32'h22ed316b;
    11'b01111011011: data <= 32'hb80b36fb;
    11'b01111011100: data <= 32'h38a73b55;
    11'b01111011101: data <= 32'h3f5b3f6e;
    11'b01111011110: data <= 32'h3d4c401f;
    11'b01111011111: data <= 32'hb6623901;
    11'b01111100000: data <= 32'hbc6cbcc1;
    11'b01111100001: data <= 32'hb010bdc0;
    11'b01111100010: data <= 32'h3c2cb5e5;
    11'b01111100011: data <= 32'h3d05ac87;
    11'b01111100100: data <= 32'h3c31bcbd;
    11'b01111100101: data <= 32'h3c1abf51;
    11'b01111100110: data <= 32'h387db87a;
    11'b01111100111: data <= 32'hba803cda;
    11'b01111101000: data <= 32'hbfd73caf;
    11'b01111101001: data <= 32'hbe5db870;
    11'b01111101010: data <= 32'hb6c8bed3;
    11'b01111101011: data <= 32'hb403bc9d;
    11'b01111101100: data <= 32'hbc55a9c7;
    11'b01111101101: data <= 32'hbc2c3721;
    11'b01111101110: data <= 32'h38583a00;
    11'b01111101111: data <= 32'h3ef23df4;
    11'b01111110000: data <= 32'h39f93fb8;
    11'b01111110001: data <= 32'hbd093ccc;
    11'b01111110010: data <= 32'hbec12a38;
    11'b01111110011: data <= 32'hafafb0ab;
    11'b01111110100: data <= 32'h3da33545;
    11'b01111110101: data <= 32'h3e14aa38;
    11'b01111110110: data <= 32'h3c43bd4b;
    11'b01111110111: data <= 32'h3c92be65;
    11'b01111111000: data <= 32'h3cec2017;
    11'b01111111001: data <= 32'h36e53e5b;
    11'b01111111010: data <= 32'hb9703b83;
    11'b01111111011: data <= 32'hbb69bcfe;
    11'b01111111100: data <= 32'hb868c0b1;
    11'b01111111101: data <= 32'hb9c5bdd4;
    11'b01111111110: data <= 32'hbd2eb432;
    11'b01111111111: data <= 32'hbadeb0d2;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    