
module memory_rom_24(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3daeb9a3;
    11'b00000000001: data <= 32'h3a09b6cc;
    11'b00000000010: data <= 32'hbb163623;
    11'b00000000011: data <= 32'hbf7faaf8;
    11'b00000000100: data <= 32'hbad7be05;
    11'b00000000101: data <= 32'h3b72c057;
    11'b00000000110: data <= 32'h3c7fbdb6;
    11'b00000000111: data <= 32'hb61bb68a;
    11'b00000001000: data <= 32'hbd672f9f;
    11'b00000001001: data <= 32'hb8fc3996;
    11'b00000001010: data <= 32'h332c3e28;
    11'b00000001011: data <= 32'hb80d3e44;
    11'b00000001100: data <= 32'hbfac330f;
    11'b00000001101: data <= 32'hbf8abc24;
    11'b00000001110: data <= 32'hb2e1b826;
    11'b00000001111: data <= 32'h3d173c38;
    11'b00000010000: data <= 32'h3e063de7;
    11'b00000010001: data <= 32'h3cf43599;
    11'b00000010010: data <= 32'h3cb5b54d;
    11'b00000010011: data <= 32'h3a3638fe;
    11'b00000010100: data <= 32'hb4813e84;
    11'b00000010101: data <= 32'hbaf83988;
    11'b00000010110: data <= 32'ha692be10;
    11'b00000010111: data <= 32'h3cc9c12f;
    11'b00000011000: data <= 32'h3c2dbf0d;
    11'b00000011001: data <= 32'hb25db850;
    11'b00000011010: data <= 32'hb899b054;
    11'b00000011011: data <= 32'h3652a368;
    11'b00000011100: data <= 32'h3a313792;
    11'b00000011101: data <= 32'hba593951;
    11'b00000011110: data <= 32'hc179ad63;
    11'b00000011111: data <= 32'hc146bac7;
    11'b00000100000: data <= 32'hb919b656;
    11'b00000100001: data <= 32'h3b5c397d;
    11'b00000100010: data <= 32'h3abd3a71;
    11'b00000100011: data <= 32'h34772854;
    11'b00000100100: data <= 32'h362a3162;
    11'b00000100101: data <= 32'h38d73eec;
    11'b00000100110: data <= 32'h30334162;
    11'b00000100111: data <= 32'hb6413d23;
    11'b00000101000: data <= 32'h2893bcea;
    11'b00000101001: data <= 32'h3b20c057;
    11'b00000101010: data <= 32'h3b79bc55;
    11'b00000101011: data <= 32'h364921b1;
    11'b00000101100: data <= 32'h3904b224;
    11'b00000101101: data <= 32'h3e51b9a2;
    11'b00000101110: data <= 32'h3d93b5a8;
    11'b00000101111: data <= 32'hb99f33c2;
    11'b00000110000: data <= 32'hc169aa41;
    11'b00000110001: data <= 32'hc0c1bab3;
    11'b00000110010: data <= 32'hb66dbb7a;
    11'b00000110011: data <= 32'h3922b68c;
    11'b00000110100: data <= 32'hac67b4ae;
    11'b00000110101: data <= 32'hba75b777;
    11'b00000110110: data <= 32'hb45b3590;
    11'b00000110111: data <= 32'h383b4049;
    11'b00000111000: data <= 32'h328f41cf;
    11'b00000111001: data <= 32'hb9c33d7f;
    11'b00000111010: data <= 32'hba5bba7b;
    11'b00000111011: data <= 32'h28c9bcc4;
    11'b00000111100: data <= 32'h39492e21;
    11'b00000111101: data <= 32'h3adf3a02;
    11'b00000111110: data <= 32'h3db8b117;
    11'b00000111111: data <= 32'h4068bc04;
    11'b00001000000: data <= 32'h3ef8b5f9;
    11'b00001000001: data <= 32'hb42f39b0;
    11'b00001000010: data <= 32'hbf6b3806;
    11'b00001000011: data <= 32'hbd4aba76;
    11'b00001000100: data <= 32'h340cbe8d;
    11'b00001000101: data <= 32'h382dbdeb;
    11'b00001000110: data <= 32'hb975bcab;
    11'b00001000111: data <= 32'hbd04bb70;
    11'b00001001000: data <= 32'hb25f24ee;
    11'b00001001001: data <= 32'h3a873e56;
    11'b00001001010: data <= 32'h2d524055;
    11'b00001001011: data <= 32'hbe253ba3;
    11'b00001001100: data <= 32'hbfe4b7be;
    11'b00001001101: data <= 32'hbb35b481;
    11'b00001001110: data <= 32'h342c3b82;
    11'b00001001111: data <= 32'h3a3b3c21;
    11'b00001010000: data <= 32'h3d13b461;
    11'b00001010001: data <= 32'h3f88bb22;
    11'b00001010010: data <= 32'h3e8c35d1;
    11'b00001010011: data <= 32'h34483f48;
    11'b00001010100: data <= 32'hb9fe3d66;
    11'b00001010101: data <= 32'hb345b8e0;
    11'b00001010110: data <= 32'h3a1cbfa1;
    11'b00001010111: data <= 32'h375abf09;
    11'b00001011000: data <= 32'hb9edbd0b;
    11'b00001011001: data <= 32'hba5cbc6e;
    11'b00001011010: data <= 32'h3956b91e;
    11'b00001011011: data <= 32'h3ddf36e2;
    11'b00001011100: data <= 32'h28a73c13;
    11'b00001011101: data <= 32'hc054366f;
    11'b00001011110: data <= 32'hc154b56d;
    11'b00001011111: data <= 32'hbd4f2bd1;
    11'b00001100000: data <= 32'hacb63b1c;
    11'b00001100001: data <= 32'h30693841;
    11'b00001100010: data <= 32'h3372b97b;
    11'b00001100011: data <= 32'h3afbb936;
    11'b00001100100: data <= 32'h3ce73d00;
    11'b00001100101: data <= 32'h38f041a2;
    11'b00001100110: data <= 32'hac953fef;
    11'b00001100111: data <= 32'h30f5b480;
    11'b00001101000: data <= 32'h3934bde0;
    11'b00001101001: data <= 32'h3453bc09;
    11'b00001101010: data <= 32'hb6b0b837;
    11'b00001101011: data <= 32'h3139bb91;
    11'b00001101100: data <= 32'h3f20bd06;
    11'b00001101101: data <= 32'h4053b893;
    11'b00001101110: data <= 32'h3323346f;
    11'b00001101111: data <= 32'hc0293306;
    11'b00001110000: data <= 32'hc0afb469;
    11'b00001110001: data <= 32'hbb94b2a7;
    11'b00001110010: data <= 32'hb1582b5d;
    11'b00001110011: data <= 32'hb99db7c5;
    11'b00001110100: data <= 32'hbc0abd24;
    11'b00001110101: data <= 32'hae41b8ee;
    11'b00001110110: data <= 32'h3b483e4c;
    11'b00001110111: data <= 32'h39b941f3;
    11'b00001111000: data <= 32'hb0723fe5;
    11'b00001111001: data <= 32'hb6459b22;
    11'b00001111010: data <= 32'haec6b864;
    11'b00001111011: data <= 32'haf8e34f9;
    11'b00001111100: data <= 32'hb06b381b;
    11'b00001111101: data <= 32'h3ac7b949;
    11'b00001111110: data <= 32'h40b8be35;
    11'b00001111111: data <= 32'h40eababc;
    11'b00010000000: data <= 32'h3896371f;
    11'b00010000001: data <= 32'hbd123934;
    11'b00010000010: data <= 32'hbca3b025;
    11'b00010000011: data <= 32'ha1d3b98d;
    11'b00010000100: data <= 32'ha81ebae9;
    11'b00010000101: data <= 32'hbd29bd4c;
    11'b00010000110: data <= 32'hbec7befb;
    11'b00010000111: data <= 32'hb56ebb45;
    11'b00010001000: data <= 32'h3c2f3c20;
    11'b00010001001: data <= 32'h3996403f;
    11'b00010001010: data <= 32'hb9ba3d32;
    11'b00010001011: data <= 32'hbd922ce7;
    11'b00010001100: data <= 32'hbc0b352a;
    11'b00010001101: data <= 32'hb87a3d84;
    11'b00010001110: data <= 32'hb39e3c7c;
    11'b00010001111: data <= 32'h396db8c3;
    11'b00010010000: data <= 32'h3fcabe19;
    11'b00010010001: data <= 32'h4045b5ac;
    11'b00010010010: data <= 32'h3b043d66;
    11'b00010010011: data <= 32'hb29d3dd5;
    11'b00010010100: data <= 32'h30d930ac;
    11'b00010010101: data <= 32'h3aaebb1e;
    11'b00010010110: data <= 32'h2f43bc70;
    11'b00010010111: data <= 32'hbda6bd64;
    11'b00010011000: data <= 32'hbdf5bf04;
    11'b00010011001: data <= 32'h34c4bd7f;
    11'b00010011010: data <= 32'h3e97ad07;
    11'b00010011011: data <= 32'h3a033a31;
    11'b00010011100: data <= 32'hbce83686;
    11'b00010011101: data <= 32'hc00da15a;
    11'b00010011110: data <= 32'hbd8e39a9;
    11'b00010011111: data <= 32'hba3a3e5a;
    11'b00010100000: data <= 32'hb9d63b03;
    11'b00010100001: data <= 32'hb523bb7b;
    11'b00010100010: data <= 32'h3a03bd95;
    11'b00010100011: data <= 32'h3d92360f;
    11'b00010100100: data <= 32'h3bd54086;
    11'b00010100101: data <= 32'h37e4401f;
    11'b00010100110: data <= 32'h3a5e3697;
    11'b00010100111: data <= 32'h3c06b869;
    11'b00010101000: data <= 32'h25ddb62b;
    11'b00010101001: data <= 32'hbcceb733;
    11'b00010101010: data <= 32'hb9b4bd20;
    11'b00010101011: data <= 32'h3d38bef5;
    11'b00010101100: data <= 32'h40a5bc58;
    11'b00010101101: data <= 32'h3b65b365;
    11'b00010101110: data <= 32'hbcc6ad9f;
    11'b00010101111: data <= 32'hbedbad05;
    11'b00010110000: data <= 32'hbaf6385b;
    11'b00010110001: data <= 32'hb8c13bb3;
    11'b00010110010: data <= 32'hbd50a09a;
    11'b00010110011: data <= 32'hbe3cbe18;
    11'b00010110100: data <= 32'hb7acbd8e;
    11'b00010110101: data <= 32'h39eb39aa;
    11'b00010110110: data <= 32'h3b4840d7;
    11'b00010110111: data <= 32'h38283fc3;
    11'b00010111000: data <= 32'h37a03748;
    11'b00010111001: data <= 32'h369930cb;
    11'b00010111010: data <= 32'hb59e3b68;
    11'b00010111011: data <= 32'hbbdf3abf;
    11'b00010111100: data <= 32'hac34b927;
    11'b00010111101: data <= 32'h3f7bbf59;
    11'b00010111110: data <= 32'h4114bdbc;
    11'b00010111111: data <= 32'h3c5bb4f4;
    11'b00011000000: data <= 32'hb88a309a;
    11'b00011000001: data <= 32'hb85128e8;
    11'b00011000010: data <= 32'h34e930a3;
    11'b00011000011: data <= 32'haeb82f77;
    11'b00011000100: data <= 32'hbecaba93;
    11'b00011000101: data <= 32'hc09cbfbe;
    11'b00011000110: data <= 32'hbbdebe30;
    11'b00011000111: data <= 32'h391c3514;
    11'b00011001000: data <= 32'h3ab43e4f;
    11'b00011001001: data <= 32'h29493c2c;
    11'b00011001010: data <= 32'hb698320e;
    11'b00011001011: data <= 32'hb7333a57;
    11'b00011001100: data <= 32'hba2b4017;
    11'b00011001101: data <= 32'hbc023ee9;
    11'b00011001110: data <= 32'hafacb4da;
    11'b00011001111: data <= 32'h3ddebee5;
    11'b00011010000: data <= 32'h400abc31;
    11'b00011010001: data <= 32'h3c443735;
    11'b00011010010: data <= 32'h343a3b13;
    11'b00011010011: data <= 32'h3a8734ef;
    11'b00011010100: data <= 32'h3dc3ad5f;
    11'b00011010101: data <= 32'h3598b28d;
    11'b00011010110: data <= 32'hbecdbadc;
    11'b00011010111: data <= 32'hc067bf21;
    11'b00011011000: data <= 32'hb82cbee2;
    11'b00011011001: data <= 32'h3c90b893;
    11'b00011011010: data <= 32'h3b1e31fc;
    11'b00011011011: data <= 32'hb769b088;
    11'b00011011100: data <= 32'hbc54b381;
    11'b00011011101: data <= 32'hbab73c1d;
    11'b00011011110: data <= 32'hbaf040b4;
    11'b00011011111: data <= 32'hbcfa3ec0;
    11'b00011100000: data <= 32'hbb50b812;
    11'b00011100001: data <= 32'h33aabe57;
    11'b00011100010: data <= 32'h3be5b59f;
    11'b00011100011: data <= 32'h3a823d75;
    11'b00011100100: data <= 32'h3a543dfc;
    11'b00011100101: data <= 32'h3e3a37d9;
    11'b00011100110: data <= 32'h3f652af7;
    11'b00011100111: data <= 32'h36f23565;
    11'b00011101000: data <= 32'hbddc2c03;
    11'b00011101001: data <= 32'hbdecbc22;
    11'b00011101010: data <= 32'h373fbee6;
    11'b00011101011: data <= 32'h3f45bd8e;
    11'b00011101100: data <= 32'h3c0bbb4d;
    11'b00011101101: data <= 32'hb8a3bb3d;
    11'b00011101110: data <= 32'hbb69b82d;
    11'b00011101111: data <= 32'hb4f43a8e;
    11'b00011110000: data <= 32'hb6f13f33;
    11'b00011110001: data <= 32'hbdf93af3;
    11'b00011110010: data <= 32'hbfcebc56;
    11'b00011110011: data <= 32'hbc55be34;
    11'b00011110100: data <= 32'h29202d63;
    11'b00011110101: data <= 32'h37b13e9a;
    11'b00011110110: data <= 32'h39f43d80;
    11'b00011110111: data <= 32'h3d4d3516;
    11'b00011111000: data <= 32'h3d7036df;
    11'b00011111001: data <= 32'h2e303dc9;
    11'b00011111010: data <= 32'hbcf03dc5;
    11'b00011111011: data <= 32'hba23ad7b;
    11'b00011111100: data <= 32'h3c7cbe14;
    11'b00011111101: data <= 32'h4017be8a;
    11'b00011111110: data <= 32'h3bfcbc5d;
    11'b00011111111: data <= 32'hb3efba91;
    11'b00100000000: data <= 32'h2addb79b;
    11'b00100000001: data <= 32'h3b93369d;
    11'b00100000010: data <= 32'h35f63b61;
    11'b00100000011: data <= 32'hbe20a55d;
    11'b00100000100: data <= 32'hc125be12;
    11'b00100000101: data <= 32'hbec9be4a;
    11'b00100000110: data <= 32'hb40daa56;
    11'b00100000111: data <= 32'h34ba3bee;
    11'b00100001000: data <= 32'h3413368d;
    11'b00100001001: data <= 32'h36fab427;
    11'b00100001010: data <= 32'h373539d3;
    11'b00100001011: data <= 32'hb59d40d9;
    11'b00100001100: data <= 32'hbc9f40e3;
    11'b00100001101: data <= 32'hb8d237d4;
    11'b00100001110: data <= 32'h3b24bcfb;
    11'b00100001111: data <= 32'h3de5bce5;
    11'b00100010000: data <= 32'h3971b5b8;
    11'b00100010001: data <= 32'h339cac76;
    11'b00100010010: data <= 32'h3d06b1d4;
    11'b00100010011: data <= 32'h40692faa;
    11'b00100010100: data <= 32'h3c6436c2;
    11'b00100010101: data <= 32'hbd50b313;
    11'b00100010110: data <= 32'hc0d8bd56;
    11'b00100010111: data <= 32'hbd23bde8;
    11'b00100011000: data <= 32'h32fcb8ce;
    11'b00100011001: data <= 32'h35a5b3a6;
    11'b00100011010: data <= 32'hb4a7bb3e;
    11'b00100011011: data <= 32'hb5ffbbe1;
    11'b00100011100: data <= 32'hadca39bb;
    11'b00100011101: data <= 32'hb70e4155;
    11'b00100011110: data <= 32'hbca840f4;
    11'b00100011111: data <= 32'hbc4d35c4;
    11'b00100100000: data <= 32'hb175bc56;
    11'b00100100001: data <= 32'h34ffb7f6;
    11'b00100100010: data <= 32'h2eae394b;
    11'b00100100011: data <= 32'h37ba3967;
    11'b00100100100: data <= 32'h3fad236f;
    11'b00100100101: data <= 32'h416b2c40;
    11'b00100100110: data <= 32'h3d3b3957;
    11'b00100100111: data <= 32'hbc23383e;
    11'b00100101000: data <= 32'hbeb5b780;
    11'b00100101001: data <= 32'hb393bc99;
    11'b00100101010: data <= 32'h3c05bc70;
    11'b00100101011: data <= 32'h3805bcfe;
    11'b00100101100: data <= 32'hb87bbf2a;
    11'b00100101101: data <= 32'hb7c6bdcc;
    11'b00100101110: data <= 32'h34493686;
    11'b00100101111: data <= 32'h2dab402d;
    11'b00100110000: data <= 32'hbc5b3e76;
    11'b00100110001: data <= 32'hbf2ab4c2;
    11'b00100110010: data <= 32'hbd91bc54;
    11'b00100110011: data <= 32'hba392b5b;
    11'b00100110100: data <= 32'hb74d3cbe;
    11'b00100110101: data <= 32'h34b039d0;
    11'b00100110110: data <= 32'h3ea0b34e;
    11'b00100110111: data <= 32'h406d3069;
    11'b00100111000: data <= 32'h3b643dcf;
    11'b00100111001: data <= 32'hbaa73f31;
    11'b00100111010: data <= 32'hbaf53916;
    11'b00100111011: data <= 32'h3923b963;
    11'b00100111100: data <= 32'h3d9fbcad;
    11'b00100111101: data <= 32'h3724bd8f;
    11'b00100111110: data <= 32'hb807bef1;
    11'b00100111111: data <= 32'h3197bd9b;
    11'b00101000000: data <= 32'h3d9c22c1;
    11'b00101000001: data <= 32'h3c383c8c;
    11'b00101000010: data <= 32'hba9a3858;
    11'b00101000011: data <= 32'hc05fbb35;
    11'b00101000100: data <= 32'hbfd8bc59;
    11'b00101000101: data <= 32'hbc8d3160;
    11'b00101000110: data <= 32'hb98f3aae;
    11'b00101000111: data <= 32'hb2c9aee6;
    11'b00101001000: data <= 32'h39acbbae;
    11'b00101001001: data <= 32'h3c9a2f6f;
    11'b00101001010: data <= 32'h350c4059;
    11'b00101001011: data <= 32'hba114180;
    11'b00101001100: data <= 32'hb7e43d41;
    11'b00101001101: data <= 32'h39aeb499;
    11'b00101001110: data <= 32'h3bd1b9a9;
    11'b00101001111: data <= 32'ha1e0b8de;
    11'b00101010000: data <= 32'hb57dbaef;
    11'b00101010001: data <= 32'h3c6abbbb;
    11'b00101010010: data <= 32'h4136b41e;
    11'b00101010011: data <= 32'h3fa8374b;
    11'b00101010100: data <= 32'hb7472b98;
    11'b00101010101: data <= 32'hbfcabb01;
    11'b00101010110: data <= 32'hbe08bafe;
    11'b00101010111: data <= 32'hb8b7ac09;
    11'b00101011000: data <= 32'hb837af06;
    11'b00101011001: data <= 32'hb9d6bd73;
    11'b00101011010: data <= 32'hb410bf61;
    11'b00101011011: data <= 32'h357baf15;
    11'b00101011100: data <= 32'h2a9d4095;
    11'b00101011101: data <= 32'hb971417e;
    11'b00101011110: data <= 32'hb9483c99;
    11'b00101011111: data <= 32'hab91b238;
    11'b00101100000: data <= 32'haf719444;
    11'b00101100001: data <= 32'hba1c384f;
    11'b00101100010: data <= 32'hb5a73001;
    11'b00101100011: data <= 32'h3e6eb8af;
    11'b00101100100: data <= 32'h4229b5de;
    11'b00101100101: data <= 32'h404536aa;
    11'b00101100110: data <= 32'hb1b83816;
    11'b00101100111: data <= 32'hbcd0adfb;
    11'b00101101000: data <= 32'hb59ab5d9;
    11'b00101101001: data <= 32'h36b7b494;
    11'b00101101010: data <= 32'hb229bb74;
    11'b00101101011: data <= 32'hbc1bc073;
    11'b00101101100: data <= 32'hb8ffc0bc;
    11'b00101101101: data <= 32'h365eb74b;
    11'b00101101110: data <= 32'h37a03ec2;
    11'b00101101111: data <= 32'hb6e63f2a;
    11'b00101110000: data <= 32'hbc4734ce;
    11'b00101110001: data <= 32'hbc45b5e4;
    11'b00101110010: data <= 32'hbcc3387f;
    11'b00101110011: data <= 32'hbdb63d31;
    11'b00101110100: data <= 32'hb91637aa;
    11'b00101110101: data <= 32'h3d2fb99a;
    11'b00101110110: data <= 32'h4103b72f;
    11'b00101110111: data <= 32'h3e623b1b;
    11'b00101111000: data <= 32'hb0353e2e;
    11'b00101111001: data <= 32'hb65b3bf5;
    11'b00101111010: data <= 32'h39f1340d;
    11'b00101111011: data <= 32'h3c7ab25e;
    11'b00101111100: data <= 32'hae42bbfd;
    11'b00101111101: data <= 32'hbc64c03a;
    11'b00101111110: data <= 32'hb460c06b;
    11'b00101111111: data <= 32'h3d21b9cf;
    11'b00110000000: data <= 32'h3dad39f0;
    11'b00110000001: data <= 32'h18453830;
    11'b00110000010: data <= 32'hbd15b8c6;
    11'b00110000011: data <= 32'hbe25b857;
    11'b00110000100: data <= 32'hbe103a31;
    11'b00110000101: data <= 32'hbe713cfe;
    11'b00110000110: data <= 32'hbc3cadc3;
    11'b00110000111: data <= 32'h3593bd94;
    11'b00110001000: data <= 32'h3d15b93a;
    11'b00110001001: data <= 32'h39a53d84;
    11'b00110001010: data <= 32'hb3bf40bd;
    11'b00110001011: data <= 32'h2b133ea0;
    11'b00110001100: data <= 32'h3c68391c;
    11'b00110001101: data <= 32'h3bc5336b;
    11'b00110001110: data <= 32'hb7f9b294;
    11'b00110001111: data <= 32'hbc7dbc61;
    11'b00110010000: data <= 32'h365ebe0f;
    11'b00110010001: data <= 32'h40acba77;
    11'b00110010010: data <= 32'h408e1f45;
    11'b00110010011: data <= 32'h36ccb3bd;
    11'b00110010100: data <= 32'hbc08baf0;
    11'b00110010101: data <= 32'hbc39b698;
    11'b00110010110: data <= 32'hbabd39c1;
    11'b00110010111: data <= 32'hbcde38a1;
    11'b00110011000: data <= 32'hbd95bcb4;
    11'b00110011001: data <= 32'hb937c093;
    11'b00110011010: data <= 32'h322bbbd3;
    11'b00110011011: data <= 32'h30323daf;
    11'b00110011100: data <= 32'hb46b40a4;
    11'b00110011101: data <= 32'h2a6c3d96;
    11'b00110011110: data <= 32'h38f8386a;
    11'b00110011111: data <= 32'h2c493a3e;
    11'b00110100000: data <= 32'hbd0c3bc2;
    11'b00110100001: data <= 32'hbd1130d8;
    11'b00110100010: data <= 32'h3a41ba85;
    11'b00110100011: data <= 32'h4180ba35;
    11'b00110100100: data <= 32'h40ddb192;
    11'b00110100101: data <= 32'h3895ad9f;
    11'b00110100110: data <= 32'hb635b4ca;
    11'b00110100111: data <= 32'h30182e7f;
    11'b00110101000: data <= 32'h36713943;
    11'b00110101001: data <= 32'hb885ad66;
    11'b00110101010: data <= 32'hbe1dbfde;
    11'b00110101011: data <= 32'hbc91c18c;
    11'b00110101100: data <= 32'haaf7bd00;
    11'b00110101101: data <= 32'h35063b3a;
    11'b00110101110: data <= 32'ha9153d5a;
    11'b00110101111: data <= 32'hb1d63554;
    11'b00110110000: data <= 32'hb23f2cb8;
    11'b00110110001: data <= 32'hbb5c3cac;
    11'b00110110010: data <= 32'hbfae3f50;
    11'b00110110011: data <= 32'hbe203a7a;
    11'b00110110100: data <= 32'h3819b946;
    11'b00110110101: data <= 32'h404bba8c;
    11'b00110110110: data <= 32'h3ed22f86;
    11'b00110110111: data <= 32'h357039cb;
    11'b00110111000: data <= 32'h33c03979;
    11'b00110111001: data <= 32'h3d3a39e4;
    11'b00110111010: data <= 32'h3da03a40;
    11'b00110111011: data <= 32'hb19ab0c5;
    11'b00110111100: data <= 32'hbe1ebf4a;
    11'b00110111101: data <= 32'hbbb8c0ed;
    11'b00110111110: data <= 32'h38abbd1a;
    11'b00110111111: data <= 32'h3c842fc7;
    11'b00111000000: data <= 32'h36c09f03;
    11'b00111000001: data <= 32'hb4d0baec;
    11'b00111000010: data <= 32'hb8f3b6a7;
    11'b00111000011: data <= 32'hbcd93d1e;
    11'b00111000100: data <= 32'hbff43fc5;
    11'b00111000101: data <= 32'hbf05380d;
    11'b00111000110: data <= 32'hb4a2bcca;
    11'b00111000111: data <= 32'h3ab8bc33;
    11'b00111001000: data <= 32'h382a37da;
    11'b00111001001: data <= 32'hae483ddc;
    11'b00111001010: data <= 32'h38903d3c;
    11'b00111001011: data <= 32'h3f483c33;
    11'b00111001100: data <= 32'h3e2b3c44;
    11'b00111001101: data <= 32'hb6363830;
    11'b00111001110: data <= 32'hbe47b9ee;
    11'b00111001111: data <= 32'hb6f3bdf6;
    11'b00111010000: data <= 32'h3e13bc1c;
    11'b00111010001: data <= 32'h3fc6b78b;
    11'b00111010010: data <= 32'h3a7dbb57;
    11'b00111010011: data <= 32'hb00ebdc2;
    11'b00111010100: data <= 32'hb338b80e;
    11'b00111010101: data <= 32'hb7c83ce4;
    11'b00111010110: data <= 32'hbd613db7;
    11'b00111010111: data <= 32'hbf19b6df;
    11'b00111011000: data <= 32'hbc8cc012;
    11'b00111011001: data <= 32'hb601bd7c;
    11'b00111011010: data <= 32'hb5fe3889;
    11'b00111011011: data <= 32'hb63c3de0;
    11'b00111011100: data <= 32'h384f3c06;
    11'b00111011101: data <= 32'h3e033a00;
    11'b00111011110: data <= 32'h3a8c3d4c;
    11'b00111011111: data <= 32'hbc533e2f;
    11'b00111100000: data <= 32'hbeee3911;
    11'b00111100001: data <= 32'hac00b756;
    11'b00111100010: data <= 32'h3fd0b9a2;
    11'b00111100011: data <= 32'h4020b8cb;
    11'b00111100100: data <= 32'h3a4cbb78;
    11'b00111100101: data <= 32'h33b9bc56;
    11'b00111100110: data <= 32'h3a83ad9a;
    11'b00111100111: data <= 32'h3b043cc3;
    11'b00111101000: data <= 32'hb5c23a87;
    11'b00111101001: data <= 32'hbe5dbcd6;
    11'b00111101010: data <= 32'hbe30c0fe;
    11'b00111101011: data <= 32'hba5ebe10;
    11'b00111101100: data <= 32'hb704341a;
    11'b00111101101: data <= 32'hb47e38e8;
    11'b00111101110: data <= 32'h3564b149;
    11'b00111101111: data <= 32'h3a2baa9c;
    11'b00111110000: data <= 32'hb01d3d89;
    11'b00111110001: data <= 32'hbee2409b;
    11'b00111110010: data <= 32'hbfa73ddd;
    11'b00111110011: data <= 32'hb185a5c2;
    11'b00111110100: data <= 32'h3dd4b8a2;
    11'b00111110101: data <= 32'h3cf8b540;
    11'b00111110110: data <= 32'h3403b371;
    11'b00111110111: data <= 32'h385db187;
    11'b00111111000: data <= 32'h3f85383f;
    11'b00111111001: data <= 32'h401c3d15;
    11'b00111111010: data <= 32'h356f391d;
    11'b00111111011: data <= 32'hbd88bc9f;
    11'b00111111100: data <= 32'hbd7dc038;
    11'b00111111101: data <= 32'hb4a5bd11;
    11'b00111111110: data <= 32'h3449b2d6;
    11'b00111111111: data <= 32'h30f8b8e9;
    11'b01000000000: data <= 32'h32a7be26;
    11'b01000000001: data <= 32'h3481bafd;
    11'b01000000010: data <= 32'hb7df3cfe;
    11'b01000000011: data <= 32'hbef140cc;
    11'b01000000100: data <= 32'hbf9b3d3f;
    11'b01000000101: data <= 32'hb97db69c;
    11'b01000000110: data <= 32'h3449ba1e;
    11'b01000000111: data <= 32'haf372870;
    11'b01000001000: data <= 32'hb847383f;
    11'b01000001001: data <= 32'h38c53806;
    11'b01000001010: data <= 32'h40b63a80;
    11'b01000001011: data <= 32'h40b63d78;
    11'b01000001100: data <= 32'h350a3c39;
    11'b01000001101: data <= 32'hbd62b210;
    11'b01000001110: data <= 32'hbae3bbcd;
    11'b01000001111: data <= 32'h390cb955;
    11'b01000010000: data <= 32'h3c6fb80e;
    11'b01000010001: data <= 32'h383ebde4;
    11'b01000010010: data <= 32'h33b6c095;
    11'b01000010011: data <= 32'h3750bcc8;
    11'b01000010100: data <= 32'h2fd53c50;
    11'b01000010101: data <= 32'hbb973f9d;
    11'b01000010110: data <= 32'hbe4e36bd;
    11'b01000010111: data <= 32'hbce3bd00;
    11'b01000011000: data <= 32'hbb13bc53;
    11'b01000011001: data <= 32'hbcd232ab;
    11'b01000011010: data <= 32'hbc6639b3;
    11'b01000011011: data <= 32'h369c34e3;
    11'b01000011100: data <= 32'h401a364e;
    11'b01000011101: data <= 32'h3ed33d36;
    11'b01000011110: data <= 32'hb5863f11;
    11'b01000011111: data <= 32'hbe043c74;
    11'b01000100000: data <= 32'hb6d4343c;
    11'b01000100001: data <= 32'h3cd0a812;
    11'b01000100010: data <= 32'h3d4eb718;
    11'b01000100011: data <= 32'h36aabdfb;
    11'b01000100100: data <= 32'h3529c015;
    11'b01000100101: data <= 32'h3ccabac7;
    11'b01000100110: data <= 32'h3da03c20;
    11'b01000100111: data <= 32'h33ec3d05;
    11'b01000101000: data <= 32'hbc35b75f;
    11'b01000101001: data <= 32'hbd9ebf33;
    11'b01000101010: data <= 32'hbd36bca7;
    11'b01000101011: data <= 32'hbda0309a;
    11'b01000101100: data <= 32'hbc6e304f;
    11'b01000101101: data <= 32'h31a9ba42;
    11'b01000101110: data <= 32'h3d37b8e6;
    11'b01000101111: data <= 32'h39863c06;
    11'b01000110000: data <= 32'hbc404089;
    11'b01000110001: data <= 32'hbe983fbd;
    11'b01000110010: data <= 32'hb5513af4;
    11'b01000110011: data <= 32'h3bae3432;
    11'b01000110100: data <= 32'h38beaef0;
    11'b01000110101: data <= 32'hb4f7ba54;
    11'b01000110110: data <= 32'h344fbc64;
    11'b01000110111: data <= 32'h3ff4b159;
    11'b01000111000: data <= 32'h41213c63;
    11'b01000111001: data <= 32'h3c923b50;
    11'b01000111010: data <= 32'hb8fbb914;
    11'b01000111011: data <= 32'hbc84be06;
    11'b01000111100: data <= 32'hba6ab9f8;
    11'b01000111101: data <= 32'hb9a42524;
    11'b01000111110: data <= 32'hb918ba7c;
    11'b01000111111: data <= 32'h29c7c042;
    11'b01001000000: data <= 32'h3981be9b;
    11'b01001000001: data <= 32'h2fff38d3;
    11'b01001000010: data <= 32'hbcb64073;
    11'b01001000011: data <= 32'hbdfd3f27;
    11'b01001000100: data <= 32'hb82a3830;
    11'b01001000101: data <= 32'h2ac02d13;
    11'b01001000110: data <= 32'hb9de341d;
    11'b01001000111: data <= 32'hbd502c31;
    11'b01001001000: data <= 32'h23ceb3e9;
    11'b01001001001: data <= 32'h40953324;
    11'b01001001010: data <= 32'h41c03c5a;
    11'b01001001011: data <= 32'h3cd13c23;
    11'b01001001100: data <= 32'hb84c2ae6;
    11'b01001001101: data <= 32'hb8d0b68a;
    11'b01001001110: data <= 32'h31fb2de8;
    11'b01001001111: data <= 32'h347a2b80;
    11'b01001010000: data <= 32'hb0debde1;
    11'b01001010001: data <= 32'h1ef5c1cc;
    11'b01001010010: data <= 32'h38d0c033;
    11'b01001010011: data <= 32'h37853559;
    11'b01001010100: data <= 32'hb7113ec4;
    11'b01001010101: data <= 32'hbb863acb;
    11'b01001010110: data <= 32'hb9abb6c7;
    11'b01001010111: data <= 32'hbb09b569;
    11'b01001011000: data <= 32'hbf603798;
    11'b01001011001: data <= 32'hc01f378c;
    11'b01001011010: data <= 32'hb51eb1fc;
    11'b01001011011: data <= 32'h3fb3b01a;
    11'b01001011100: data <= 32'h40643a7d;
    11'b01001011101: data <= 32'h37873d93;
    11'b01001011110: data <= 32'hba383c7b;
    11'b01001011111: data <= 32'hb0863ad2;
    11'b01001100000: data <= 32'h3b993b76;
    11'b01001100001: data <= 32'h39ed3537;
    11'b01001100010: data <= 32'hb1c6bd9c;
    11'b01001100011: data <= 32'hae23c144;
    11'b01001100100: data <= 32'h3c00bee2;
    11'b01001100101: data <= 32'h3e073578;
    11'b01001100110: data <= 32'h3a2e3c18;
    11'b01001100111: data <= 32'hb1d2b238;
    11'b01001101000: data <= 32'hb91ebccd;
    11'b01001101001: data <= 32'hbcb9b82c;
    11'b01001101010: data <= 32'hc019387d;
    11'b01001101011: data <= 32'hc02c32f1;
    11'b01001101100: data <= 32'hb851bc15;
    11'b01001101101: data <= 32'h3ca0bc92;
    11'b01001101110: data <= 32'h3c2c343c;
    11'b01001101111: data <= 32'hb74c3e6c;
    11'b01001110000: data <= 32'hbc243f32;
    11'b01001110001: data <= 32'h2ca63dea;
    11'b01001110010: data <= 32'h3c063d30;
    11'b01001110011: data <= 32'h34373988;
    11'b01001110100: data <= 32'hbb36b95e;
    11'b01001110101: data <= 32'hb666be50;
    11'b01001110110: data <= 32'h3de9bad8;
    11'b01001110111: data <= 32'h41003831;
    11'b01001111000: data <= 32'h3ed138bc;
    11'b01001111001: data <= 32'h35ebb929;
    11'b01001111010: data <= 32'hb47dbca9;
    11'b01001111011: data <= 32'hb91bb024;
    11'b01001111100: data <= 32'hbd0e396d;
    11'b01001111101: data <= 32'hbddab670;
    11'b01001111110: data <= 32'hb878c060;
    11'b01001111111: data <= 32'h3793c075;
    11'b01010000000: data <= 32'h3323b4ea;
    11'b01010000001: data <= 32'hbaaa3db4;
    11'b01010000010: data <= 32'hbb763e5f;
    11'b01010000011: data <= 32'h2ed83c4f;
    11'b01010000100: data <= 32'h36dc3c06;
    11'b01010000101: data <= 32'hbaf23bb3;
    11'b01010000110: data <= 32'hbfe33391;
    11'b01010000111: data <= 32'hbae2b7f5;
    11'b01010001000: data <= 32'h3e62b27e;
    11'b01010001001: data <= 32'h417738b8;
    11'b01010001010: data <= 32'h3ef4381d;
    11'b01010001011: data <= 32'h3664b48c;
    11'b01010001100: data <= 32'h31e0b468;
    11'b01010001101: data <= 32'h364a3a14;
    11'b01010001110: data <= 32'hacc23b9a;
    11'b01010001111: data <= 32'hb9c8bab4;
    11'b01010010000: data <= 32'hb7fcc1b9;
    11'b01010010001: data <= 32'h32fbc15b;
    11'b01010010010: data <= 32'h33e3b89a;
    11'b01010010011: data <= 32'hb51f3b51;
    11'b01010010100: data <= 32'hb55c38e4;
    11'b01010010101: data <= 32'h3160aa0a;
    11'b01010010110: data <= 32'hb3f03594;
    11'b01010010111: data <= 32'hbf7d3c44;
    11'b01010011000: data <= 32'hc1773a43;
    11'b01010011001: data <= 32'hbd01b002;
    11'b01010011010: data <= 32'h3cd3b501;
    11'b01010011011: data <= 32'h400234b3;
    11'b01010011100: data <= 32'h3ad938f8;
    11'b01010011101: data <= 32'haae43805;
    11'b01010011110: data <= 32'h38393aed;
    11'b01010011111: data <= 32'h3d173e9f;
    11'b01010100000: data <= 32'h397c3d4f;
    11'b01010100001: data <= 32'hb7e4b99d;
    11'b01010100010: data <= 32'hb8bfc117;
    11'b01010100011: data <= 32'h35f6c05d;
    11'b01010100100: data <= 32'h3be3b642;
    11'b01010100101: data <= 32'h3a1135aa;
    11'b01010100110: data <= 32'h37efb842;
    11'b01010100111: data <= 32'h3653bc6f;
    11'b01010101000: data <= 32'hb6ffaea8;
    11'b01010101001: data <= 32'hc00b3c76;
    11'b01010101010: data <= 32'hc15c3a0a;
    11'b01010101011: data <= 32'hbd5bb935;
    11'b01010101100: data <= 32'h3834bcb0;
    11'b01010101101: data <= 32'h3a1db54b;
    11'b01010101110: data <= 32'hb56e3915;
    11'b01010101111: data <= 32'hb8b03c1d;
    11'b01010110000: data <= 32'h396d3dbb;
    11'b01010110001: data <= 32'h3e253fed;
    11'b01010110010: data <= 32'h382e3e76;
    11'b01010110011: data <= 32'hbc25a7f3;
    11'b01010110100: data <= 32'hbbbfbda3;
    11'b01010110101: data <= 32'h3903bc47;
    11'b01010110110: data <= 32'h3f2a2c1a;
    11'b01010110111: data <= 32'h3e811dc4;
    11'b01010111000: data <= 32'h3c35bcaf;
    11'b01010111001: data <= 32'h39e5bd92;
    11'b01010111010: data <= 32'h2d072d87;
    11'b01010111011: data <= 32'hbca93d27;
    11'b01010111100: data <= 32'hbf5835f1;
    11'b01010111101: data <= 32'hbc64be66;
    11'b01010111110: data <= 32'habeac05f;
    11'b01010111111: data <= 32'hb346bb89;
    11'b01011000000: data <= 32'hbc2936a0;
    11'b01011000001: data <= 32'hb9b03a7c;
    11'b01011000010: data <= 32'h39f73bc3;
    11'b01011000011: data <= 32'h3cca3e08;
    11'b01011000100: data <= 32'hb5e53e9c;
    11'b01011000101: data <= 32'hc00c3a38;
    11'b01011000110: data <= 32'hbdfab184;
    11'b01011000111: data <= 32'h3936add7;
    11'b01011001000: data <= 32'h3fe5361e;
    11'b01011001001: data <= 32'h3e6cad12;
    11'b01011001010: data <= 32'h3b89bc30;
    11'b01011001011: data <= 32'h3c08ba1d;
    11'b01011001100: data <= 32'h3c133b04;
    11'b01011001101: data <= 32'h314c3e90;
    11'b01011001110: data <= 32'hba332c9f;
    11'b01011001111: data <= 32'hba1ec061;
    11'b01011010000: data <= 32'hb4c0c12d;
    11'b01011010001: data <= 32'hb6fbbc78;
    11'b01011010010: data <= 32'hba7b29f0;
    11'b01011010011: data <= 32'hb381ae38;
    11'b01011010100: data <= 32'h3b25b484;
    11'b01011010101: data <= 32'h3986385a;
    11'b01011010110: data <= 32'hbd073de4;
    11'b01011010111: data <= 32'hc17d3d1e;
    11'b01011011000: data <= 32'hbf5a36c9;
    11'b01011011001: data <= 32'h35a02eae;
    11'b01011011010: data <= 32'h3d2e3396;
    11'b01011011011: data <= 32'h38e0aaec;
    11'b01011011100: data <= 32'h3299b74d;
    11'b01011011101: data <= 32'h3c49337d;
    11'b01011011110: data <= 32'h3f583ef2;
    11'b01011011111: data <= 32'h3c8f4008;
    11'b01011100000: data <= 32'hb30f3182;
    11'b01011100001: data <= 32'hb963bf97;
    11'b01011100010: data <= 32'hb2a9bffa;
    11'b01011100011: data <= 32'h2db1b977;
    11'b01011100100: data <= 32'h2e2cb404;
    11'b01011100101: data <= 32'h3878bcaf;
    11'b01011100110: data <= 32'h3ca0be33;
    11'b01011100111: data <= 32'h3821b3e9;
    11'b01011101000: data <= 32'hbda23d35;
    11'b01011101001: data <= 32'hc1393d2d;
    11'b01011101010: data <= 32'hbede2fee;
    11'b01011101011: data <= 32'hae07b86b;
    11'b01011101100: data <= 32'h2fddb568;
    11'b01011101101: data <= 32'hba42aeaf;
    11'b01011101110: data <= 32'hb9601ece;
    11'b01011101111: data <= 32'h3bcc3a3c;
    11'b01011110000: data <= 32'h403d4003;
    11'b01011110001: data <= 32'h3cd64049;
    11'b01011110010: data <= 32'hb83b3929;
    11'b01011110011: data <= 32'hbbd0ba98;
    11'b01011110100: data <= 32'ha85db98e;
    11'b01011110101: data <= 32'h3a542f78;
    11'b01011110110: data <= 32'h3b56b558;
    11'b01011110111: data <= 32'h3c50bf3e;
    11'b01011111000: data <= 32'h3d8fc024;
    11'b01011111001: data <= 32'h3b06b52b;
    11'b01011111010: data <= 32'hb8d93d7e;
    11'b01011111011: data <= 32'hbe653bf2;
    11'b01011111100: data <= 32'hbc92b982;
    11'b01011111101: data <= 32'hb685bdf8;
    11'b01011111110: data <= 32'hbad6bb6b;
    11'b01011111111: data <= 32'hbee7b44f;
    11'b01100000000: data <= 32'hbc60aeb6;
    11'b01100000001: data <= 32'h3b4235c1;
    11'b01100000010: data <= 32'h3f6d3d8b;
    11'b01100000011: data <= 32'h37b23f7c;
    11'b01100000100: data <= 32'hbda83cba;
    11'b01100000101: data <= 32'hbdf13638;
    11'b01100000110: data <= 32'h1a23383e;
    11'b01100000111: data <= 32'h3c1f3a17;
    11'b01100001000: data <= 32'h3b6cb3f8;
    11'b01100001001: data <= 32'h3ad0bf03;
    11'b01100001010: data <= 32'h3d8fbe82;
    11'b01100001011: data <= 32'h3e3e355d;
    11'b01100001100: data <= 32'h398e3ed3;
    11'b01100001101: data <= 32'hb4a739b9;
    11'b01100001110: data <= 32'hb75abd2b;
    11'b01100001111: data <= 32'hb708bfa6;
    11'b01100010000: data <= 32'hbc79bc10;
    11'b01100010001: data <= 32'hbed0b69c;
    11'b01100010010: data <= 32'hba48ba42;
    11'b01100010011: data <= 32'h3c17badd;
    11'b01100010100: data <= 32'h3d9431e7;
    11'b01100010101: data <= 32'hb6253d50;
    11'b01100010110: data <= 32'hc0473dcf;
    11'b01100010111: data <= 32'hbf163c1c;
    11'b01100011000: data <= 32'hafe23ba7;
    11'b01100011001: data <= 32'h38643a9a;
    11'b01100011010: data <= 32'ha852b16a;
    11'b01100011011: data <= 32'haec6bce4;
    11'b01100011100: data <= 32'h3c5fb980;
    11'b01100011101: data <= 32'h40423cba;
    11'b01100011110: data <= 32'h3ecc4018;
    11'b01100011111: data <= 32'h381d3986;
    11'b01100100000: data <= 32'haf5dbca4;
    11'b01100100001: data <= 32'hb43ebd68;
    11'b01100100010: data <= 32'hb94db621;
    11'b01100100011: data <= 32'hbb1fb5d9;
    11'b01100100100: data <= 32'ha66ebe68;
    11'b01100100101: data <= 32'h3d15c04b;
    11'b01100100110: data <= 32'h3c91bafc;
    11'b01100100111: data <= 32'hb9473ae9;
    11'b01100101000: data <= 32'hc0143d62;
    11'b01100101001: data <= 32'hbded3a64;
    11'b01100101010: data <= 32'hb40636db;
    11'b01100101011: data <= 32'hb5fe3501;
    11'b01100101100: data <= 32'hbdc4b2d0;
    11'b01100101101: data <= 32'hbd09b9c5;
    11'b01100101110: data <= 32'h395aaa91;
    11'b01100101111: data <= 32'h40833df5;
    11'b01100110000: data <= 32'h3f5a4014;
    11'b01100110001: data <= 32'h35e83b0e;
    11'b01100110010: data <= 32'hb512b52a;
    11'b01100110011: data <= 32'had21a93a;
    11'b01100110100: data <= 32'h29b7398d;
    11'b01100110101: data <= 32'ha2f9ae4e;
    11'b01100110110: data <= 32'h3842c01d;
    11'b01100110111: data <= 32'h3da0c178;
    11'b01100111000: data <= 32'h3d0ebc95;
    11'b01100111001: data <= 32'hacde3a4e;
    11'b01100111010: data <= 32'hbc183c12;
    11'b01100111011: data <= 32'hb9171d8c;
    11'b01100111100: data <= 32'hb281b840;
    11'b01100111101: data <= 32'hbc98b4ef;
    11'b01100111110: data <= 32'hc0e6b50c;
    11'b01100111111: data <= 32'hbfa4b91e;
    11'b01101000000: data <= 32'h3689b45e;
    11'b01101000001: data <= 32'h3fc53b04;
    11'b01101000010: data <= 32'h3c943e10;
    11'b01101000011: data <= 32'hb7fb3c3b;
    11'b01101000100: data <= 32'hbabf3966;
    11'b01101000101: data <= 32'h9f783d01;
    11'b01101000110: data <= 32'h36eb3e65;
    11'b01101000111: data <= 32'h317a3334;
    11'b01101001000: data <= 32'h353dbfaf;
    11'b01101001001: data <= 32'h3cbcc0ae;
    11'b01101001010: data <= 32'h3e66b856;
    11'b01101001011: data <= 32'h3c023c75;
    11'b01101001100: data <= 32'h359839c1;
    11'b01101001101: data <= 32'h3551b9a6;
    11'b01101001110: data <= 32'h29e7bc66;
    11'b01101001111: data <= 32'hbd3bb6eb;
    11'b01101010000: data <= 32'hc0fbb463;
    11'b01101010001: data <= 32'hbecabbf8;
    11'b01101010010: data <= 32'h37c2bd13;
    11'b01101010011: data <= 32'h3ddbb623;
    11'b01101010100: data <= 32'h32963962;
    11'b01101010101: data <= 32'hbd623c0b;
    11'b01101010110: data <= 32'hbcb23cbc;
    11'b01101010111: data <= 32'h22823f03;
    11'b01101011000: data <= 32'h33963f37;
    11'b01101011001: data <= 32'hb8983625;
    11'b01101011010: data <= 32'hb96bbd7c;
    11'b01101011011: data <= 32'h38b0bd6a;
    11'b01101011100: data <= 32'h3f4f3669;
    11'b01101011101: data <= 32'h3f6d3e05;
    11'b01101011110: data <= 32'h3cf838ac;
    11'b01101011111: data <= 32'h3aecba98;
    11'b01101100000: data <= 32'h358db9f9;
    11'b01101100001: data <= 32'hba92336e;
    11'b01101100010: data <= 32'hbea22bf0;
    11'b01101100011: data <= 32'hbafbbddd;
    11'b01101100100: data <= 32'h3a40c0c7;
    11'b01101100101: data <= 32'h3c86be26;
    11'b01101100110: data <= 32'hb491a65b;
    11'b01101100111: data <= 32'hbdc839d2;
    11'b01101101000: data <= 32'hbaf73b42;
    11'b01101101001: data <= 32'h30d13cee;
    11'b01101101010: data <= 32'hb5713d11;
    11'b01101101011: data <= 32'hbf3734de;
    11'b01101101100: data <= 32'hbfbaba83;
    11'b01101101101: data <= 32'haed2b848;
    11'b01101101110: data <= 32'h3eeb3b2c;
    11'b01101101111: data <= 32'h3fb53e06;
    11'b01101110000: data <= 32'h3c87384e;
    11'b01101110001: data <= 32'h397db522;
    11'b01101110010: data <= 32'h382a3619;
    11'b01101110011: data <= 32'hacc33da4;
    11'b01101110100: data <= 32'hb90e38fb;
    11'b01101110101: data <= 32'hb066bea1;
    11'b01101110110: data <= 32'h3b97c1c8;
    11'b01101110111: data <= 32'h3c35bf7a;
    11'b01101111000: data <= 32'ha4b3b19a;
    11'b01101111001: data <= 32'hb8f035fb;
    11'b01101111010: data <= 32'h2c712d28;
    11'b01101111011: data <= 32'h380b30f9;
    11'b01101111100: data <= 32'hba9337c5;
    11'b01101111101: data <= 32'hc16c30de;
    11'b01101111110: data <= 32'hc154b889;
    11'b01101111111: data <= 32'hb7ebb764;
    11'b01110000000: data <= 32'h3d6337ab;
    11'b01110000001: data <= 32'h3ccb3b39;
    11'b01110000010: data <= 32'h31b6367d;
    11'b01110000011: data <= 32'h270235d5;
    11'b01110000100: data <= 32'h38493e3e;
    11'b01110000101: data <= 32'h371c40d7;
    11'b01110000110: data <= 32'hb1a23c80;
    11'b01110000111: data <= 32'hb080bda0;
    11'b01110001000: data <= 32'h395cc0e8;
    11'b01110001001: data <= 32'h3c5cbcd9;
    11'b01110001010: data <= 32'h39e533ec;
    11'b01110001011: data <= 32'h3912301d;
    11'b01110001100: data <= 32'h3ca5b9e0;
    11'b01110001101: data <= 32'h3bd9b943;
    11'b01110001110: data <= 32'hba9530f7;
    11'b01110001111: data <= 32'hc168330b;
    11'b01110010000: data <= 32'hc0deb92f;
    11'b01110010001: data <= 32'hb5d9bc87;
    11'b01110010010: data <= 32'h3b3eb92d;
    11'b01110010011: data <= 32'h318eacb5;
    11'b01110010100: data <= 32'hbb192e05;
    11'b01110010101: data <= 32'hb8123967;
    11'b01110010110: data <= 32'h386f4004;
    11'b01110010111: data <= 32'h37ec4149;
    11'b01110011000: data <= 32'hb8cb3d20;
    11'b01110011001: data <= 32'hbbf9baf2;
    11'b01110011010: data <= 32'hab9ebd94;
    11'b01110011011: data <= 32'h3c1aacf2;
    11'b01110011100: data <= 32'h3d6e3ab2;
    11'b01110011101: data <= 32'h3ddf248b;
    11'b01110011110: data <= 32'h3f03bc46;
    11'b01110011111: data <= 32'h3d58b8f0;
    11'b01110100000: data <= 32'hb50c393f;
    11'b01110100001: data <= 32'hbf3a3966;
    11'b01110100010: data <= 32'hbdc8ba82;
    11'b01110100011: data <= 32'h2f5fbff8;
    11'b01110100100: data <= 32'h38e5bef2;
    11'b01110100101: data <= 32'hb80cbaed;
    11'b01110100110: data <= 32'hbd29b4d7;
    11'b01110100111: data <= 32'hb6293575;
    11'b01110101000: data <= 32'h3a503dbb;
    11'b01110101001: data <= 32'h330f3feb;
    11'b01110101010: data <= 32'hbe343c2b;
    11'b01110101011: data <= 32'hc05bb5b8;
    11'b01110101100: data <= 32'hbb00b695;
    11'b01110101101: data <= 32'h3a1339b0;
    11'b01110101110: data <= 32'h3d523c22;
    11'b01110101111: data <= 32'h3d3cae54;
    11'b01110110000: data <= 32'h3df5badd;
    11'b01110110001: data <= 32'h3d8d330a;
    11'b01110110010: data <= 32'h36353f01;
    11'b01110110011: data <= 32'hb9183d81;
    11'b01110110100: data <= 32'hb6e4ba54;
    11'b01110110101: data <= 32'h37e1c0b7;
    11'b01110110110: data <= 32'h37d4c00d;
    11'b01110110111: data <= 32'hb823bbd5;
    11'b01110111000: data <= 32'hba15b8ab;
    11'b01110111001: data <= 32'h3755b74d;
    11'b01110111010: data <= 32'h3d2c336c;
    11'b01110111011: data <= 32'ha2e43b81;
    11'b01110111100: data <= 32'hc095395f;
    11'b01110111101: data <= 32'hc1bfae20;
    11'b01110111110: data <= 32'hbd18acf4;
    11'b01110111111: data <= 32'h364938cf;
    11'b01111000000: data <= 32'h38db385e;
    11'b01111000001: data <= 32'h33f7b60e;
    11'b01111000010: data <= 32'h38c8b717;
    11'b01111000011: data <= 32'h3cc03cd3;
    11'b01111000100: data <= 32'h3b304175;
    11'b01111000101: data <= 32'h2ba43fbc;
    11'b01111000110: data <= 32'haf99b801;
    11'b01111000111: data <= 32'h35b1bf97;
    11'b01111001000: data <= 32'h364cbd1c;
    11'b01111001001: data <= 32'ha9f7b5bc;
    11'b01111001010: data <= 32'h3468b90b;
    11'b01111001011: data <= 32'h3e15bd00;
    11'b01111001100: data <= 32'h3f75ba6a;
    11'b01111001101: data <= 32'h2d1c349f;
    11'b01111001110: data <= 32'hc076388f;
    11'b01111001111: data <= 32'hc122ac2c;
    11'b01111010000: data <= 32'hbbe9b74f;
    11'b01111010001: data <= 32'h2fbfb49b;
    11'b01111010010: data <= 32'hb648b657;
    11'b01111010011: data <= 32'hbc13ba8b;
    11'b01111010100: data <= 32'hb417b468;
    11'b01111010101: data <= 32'h3c0c3e4f;
    11'b01111010110: data <= 32'h3c2241cb;
    11'b01111010111: data <= 32'hacce3fee;
    11'b01111011000: data <= 32'hb9baadec;
    11'b01111011001: data <= 32'hb53abadc;
    11'b01111011010: data <= 32'h31c72993;
    11'b01111011011: data <= 32'h36363850;
    11'b01111011100: data <= 32'h3c09b83e;
    11'b01111011101: data <= 32'h4027be90;
    11'b01111011110: data <= 32'h4054bc2c;
    11'b01111011111: data <= 32'h38063814;
    11'b01111100000: data <= 32'hbd5f3ba4;
    11'b01111100001: data <= 32'hbda6acd6;
    11'b01111100010: data <= 32'hb2e5bc64;
    11'b01111100011: data <= 32'h29c1bd01;
    11'b01111100100: data <= 32'hbc6fbcaf;
    11'b01111100101: data <= 32'hbec8bcdb;
    11'b01111100110: data <= 32'hb6e3b89d;
    11'b01111100111: data <= 32'h3c993bfb;
    11'b01111101000: data <= 32'h3b43402c;
    11'b01111101001: data <= 32'hba443de8;
    11'b01111101010: data <= 32'hbefd328d;
    11'b01111101011: data <= 32'hbc8c30c0;
    11'b01111101100: data <= 32'hb0583c66;
    11'b01111101101: data <= 32'h35753c35;
    11'b01111101110: data <= 32'h3aa3b829;
    11'b01111101111: data <= 32'h3ec9be44;
    11'b01111110000: data <= 32'h3ff3b770;
    11'b01111110001: data <= 32'h3c083db9;
    11'b01111110010: data <= 32'hb11c3e9c;
    11'b01111110011: data <= 32'hb06528c7;
    11'b01111110100: data <= 32'h37e0bd92;
    11'b01111110101: data <= 32'h2d02be04;
    11'b01111110110: data <= 32'hbcf5bccb;
    11'b01111110111: data <= 32'hbdbfbd44;
    11'b01111111000: data <= 32'h32cdbcd0;
    11'b01111111001: data <= 32'h3e92b2cb;
    11'b01111111010: data <= 32'h3a573a61;
    11'b01111111011: data <= 32'hbda43a25;
    11'b01111111100: data <= 32'hc0c7348e;
    11'b01111111101: data <= 32'hbdeb38ac;
    11'b01111111110: data <= 32'hb6103d15;
    11'b01111111111: data <= 32'hb3f83a58;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    