
module memory_rom_54(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3caebc3c;
    11'b00000000001: data <= 32'h392bb971;
    11'b00000000010: data <= 32'hb95638a4;
    11'b00000000011: data <= 32'hbf2a384e;
    11'b00000000100: data <= 32'hbd42bc70;
    11'b00000000101: data <= 32'h329dc0aa;
    11'b00000000110: data <= 32'h3987bf03;
    11'b00000000111: data <= 32'hb6afb572;
    11'b00000001000: data <= 32'hbd0a37b4;
    11'b00000001001: data <= 32'hb7633aa0;
    11'b00000001010: data <= 32'h391a3d87;
    11'b00000001011: data <= 32'h28f53ea2;
    11'b00000001100: data <= 32'hbed23a99;
    11'b00000001101: data <= 32'hc048b695;
    11'b00000001110: data <= 32'hb761b78a;
    11'b00000001111: data <= 32'h3dd938c5;
    11'b00000010000: data <= 32'h3f883c02;
    11'b00000010001: data <= 32'h3d4028bd;
    11'b00000010010: data <= 32'h3c23b94d;
    11'b00000010011: data <= 32'h3b8434cc;
    11'b00000010100: data <= 32'h33d63e76;
    11'b00000010101: data <= 32'hb8e83c00;
    11'b00000010110: data <= 32'hb7e8bd55;
    11'b00000010111: data <= 32'h35e4c1a1;
    11'b00000011000: data <= 32'h3826c020;
    11'b00000011001: data <= 32'hb4e2b81f;
    11'b00000011010: data <= 32'hb8e228cb;
    11'b00000011011: data <= 32'h351fb004;
    11'b00000011100: data <= 32'h3b28325e;
    11'b00000011101: data <= 32'hb7703ac5;
    11'b00000011110: data <= 32'hc12739e1;
    11'b00000011111: data <= 32'hc1a7a60a;
    11'b00000100000: data <= 32'hbab5b2d0;
    11'b00000100001: data <= 32'h3c2135d9;
    11'b00000100010: data <= 32'h3c4a385c;
    11'b00000100011: data <= 32'h34cba5b5;
    11'b00000100100: data <= 32'h363421c1;
    11'b00000100101: data <= 32'h3c3a3d9e;
    11'b00000100110: data <= 32'h3b754112;
    11'b00000100111: data <= 32'h28473dcc;
    11'b00000101000: data <= 32'hb541bc50;
    11'b00000101001: data <= 32'h3263c0ac;
    11'b00000101010: data <= 32'h38abbd84;
    11'b00000101011: data <= 32'h363cb024;
    11'b00000101100: data <= 32'h3825b52f;
    11'b00000101101: data <= 32'h3d1ebc71;
    11'b00000101110: data <= 32'h3d1dba4c;
    11'b00000101111: data <= 32'hb7db3630;
    11'b00000110000: data <= 32'hc11839fd;
    11'b00000110001: data <= 32'hc128ac96;
    11'b00000110010: data <= 32'hb9f7ba28;
    11'b00000110011: data <= 32'h37cbb8c6;
    11'b00000110100: data <= 32'hae36b443;
    11'b00000110101: data <= 32'hbb36b319;
    11'b00000110110: data <= 32'hb33935b4;
    11'b00000110111: data <= 32'h3c533f50;
    11'b00000111000: data <= 32'h3c4c4175;
    11'b00000111001: data <= 32'hb36c3e7a;
    11'b00000111010: data <= 32'hbbf6b77c;
    11'b00000111011: data <= 32'hb5b7bcb0;
    11'b00000111100: data <= 32'h3903b100;
    11'b00000111101: data <= 32'h3c1e37c1;
    11'b00000111110: data <= 32'h3d36b7e7;
    11'b00000111111: data <= 32'h3f38be51;
    11'b00001000000: data <= 32'h3e6ebb72;
    11'b00001000001: data <= 32'h2a053991;
    11'b00001000010: data <= 32'hbe5a3c32;
    11'b00001000011: data <= 32'hbe2fb505;
    11'b00001000100: data <= 32'hb481be72;
    11'b00001000101: data <= 32'h2e6ebe60;
    11'b00001000110: data <= 32'hbb76bb96;
    11'b00001000111: data <= 32'hbdf3b860;
    11'b00001001000: data <= 32'hb45527e1;
    11'b00001001001: data <= 32'h3cd13ce4;
    11'b00001001010: data <= 32'h3a334017;
    11'b00001001011: data <= 32'hbc743daa;
    11'b00001001100: data <= 32'hc01330ac;
    11'b00001001101: data <= 32'hbc15a8fb;
    11'b00001001110: data <= 32'h377d3a53;
    11'b00001001111: data <= 32'h3c253a73;
    11'b00001010000: data <= 32'h3c81b86f;
    11'b00001010001: data <= 32'h3e1abd9d;
    11'b00001010010: data <= 32'h3ec1b2ec;
    11'b00001010011: data <= 32'h3ab53e73;
    11'b00001010100: data <= 32'hb4ba3e49;
    11'b00001010101: data <= 32'hb6a5b69d;
    11'b00001010110: data <= 32'h314fc007;
    11'b00001010111: data <= 32'ha68abf6c;
    11'b00001011000: data <= 32'hbc21bc17;
    11'b00001011001: data <= 32'hbc7cbaa0;
    11'b00001011010: data <= 32'h35f0ba90;
    11'b00001011011: data <= 32'h3e1aabeb;
    11'b00001011100: data <= 32'h36e33b7a;
    11'b00001011101: data <= 32'hbf793c1c;
    11'b00001011110: data <= 32'hc1593762;
    11'b00001011111: data <= 32'hbd5d36bd;
    11'b00001100000: data <= 32'h30a63ae5;
    11'b00001100001: data <= 32'h34d53822;
    11'b00001100010: data <= 32'h25a9b963;
    11'b00001100011: data <= 32'h38d0bb50;
    11'b00001100100: data <= 32'h3e0839ee;
    11'b00001100101: data <= 32'h3dbb40f7;
    11'b00001100110: data <= 32'h38544002;
    11'b00001100111: data <= 32'h2c71b2b7;
    11'b00001101000: data <= 32'h324ebe52;
    11'b00001101001: data <= 32'h9d8bbc5d;
    11'b00001101010: data <= 32'hb850b63b;
    11'b00001101011: data <= 32'hb162bb3f;
    11'b00001101100: data <= 32'h3d1cbecf;
    11'b00001101101: data <= 32'h3fb8bce7;
    11'b00001101110: data <= 32'h367f3095;
    11'b00001101111: data <= 32'hbf693a76;
    11'b00001110000: data <= 32'hc0b736f4;
    11'b00001110001: data <= 32'hbc272ce9;
    11'b00001110010: data <= 32'hb0a02eb1;
    11'b00001110011: data <= 32'hba1eb368;
    11'b00001110100: data <= 32'hbd62bb5f;
    11'b00001110101: data <= 32'hb59bb8f4;
    11'b00001110110: data <= 32'h3d133c9a;
    11'b00001110111: data <= 32'h3e47413e;
    11'b00001111000: data <= 32'h37df4004;
    11'b00001111001: data <= 32'hb5c931db;
    11'b00001111010: data <= 32'hb467b815;
    11'b00001111011: data <= 32'ha6fa349d;
    11'b00001111100: data <= 32'h1f44387f;
    11'b00001111101: data <= 32'h3895ba55;
    11'b00001111110: data <= 32'h3f0fc048;
    11'b00001111111: data <= 32'h4048be58;
    11'b00010000000: data <= 32'h3a2a31fa;
    11'b00010000001: data <= 32'hbbcc3bf2;
    11'b00010000010: data <= 32'hbcb9342c;
    11'b00010000011: data <= 32'hb3e0b918;
    11'b00010000100: data <= 32'hb393ba8f;
    11'b00010000101: data <= 32'hbe35bb17;
    11'b00010000110: data <= 32'hc04cbcb7;
    11'b00010000111: data <= 32'hb983ba91;
    11'b00010001000: data <= 32'h3cf738e2;
    11'b00010001001: data <= 32'h3d523f3f;
    11'b00010001010: data <= 32'hb37d3dfd;
    11'b00010001011: data <= 32'hbd333807;
    11'b00010001100: data <= 32'hbb533881;
    11'b00010001101: data <= 32'hb13e3dcf;
    11'b00010001110: data <= 32'h2d993cd1;
    11'b00010001111: data <= 32'h3720b955;
    11'b00010010000: data <= 32'h3d86c005;
    11'b00010010001: data <= 32'h3fcabc2f;
    11'b00010010010: data <= 32'h3d203bbe;
    11'b00010010011: data <= 32'h34053df3;
    11'b00010010100: data <= 32'h31593192;
    11'b00010010101: data <= 32'h385bbc41;
    11'b00010010110: data <= 32'hb093bc72;
    11'b00010010111: data <= 32'hbeb9bb0f;
    11'b00010011000: data <= 32'hbfe6bceb;
    11'b00010011001: data <= 32'hb2edbdab;
    11'b00010011010: data <= 32'h3e15b8d7;
    11'b00010011011: data <= 32'h3c1637d7;
    11'b00010011100: data <= 32'hbbc53a03;
    11'b00010011101: data <= 32'hbfca388d;
    11'b00010011110: data <= 32'hbcba3c25;
    11'b00010011111: data <= 32'hb4e73ef0;
    11'b00010100000: data <= 32'hb6d73c7c;
    11'b00010100001: data <= 32'hb8bcb9c3;
    11'b00010100010: data <= 32'h3426be49;
    11'b00010100011: data <= 32'h3da0b08d;
    11'b00010100100: data <= 32'h3e6b3f50;
    11'b00010100101: data <= 32'h3c583f8d;
    11'b00010100110: data <= 32'h3b0833e9;
    11'b00010100111: data <= 32'h3a96ba78;
    11'b00010101000: data <= 32'ha6f2b68d;
    11'b00010101001: data <= 32'hbcf9ac95;
    11'b00010101010: data <= 32'hbc6ebbb0;
    11'b00010101011: data <= 32'h3943c009;
    11'b00010101100: data <= 32'h3fa1bf05;
    11'b00010101101: data <= 32'h3b4db856;
    11'b00010101110: data <= 32'hbc6033be;
    11'b00010101111: data <= 32'hbebf368e;
    11'b00010110000: data <= 32'hb9d239fb;
    11'b00010110001: data <= 32'hb4663c61;
    11'b00010110010: data <= 32'hbcde36f0;
    11'b00010110011: data <= 32'hbfbfbbab;
    11'b00010110100: data <= 32'hbb88bced;
    11'b00010110101: data <= 32'h3abf35e0;
    11'b00010110110: data <= 32'h3e48400a;
    11'b00010110111: data <= 32'h3c593f13;
    11'b00010111000: data <= 32'h38c935aa;
    11'b00010111001: data <= 32'h372e962f;
    11'b00010111010: data <= 32'ha8873b8b;
    11'b00010111011: data <= 32'hb97d3c85;
    11'b00010111100: data <= 32'hb4d8b7f3;
    11'b00010111101: data <= 32'h3cc5c081;
    11'b00010111110: data <= 32'h400ec050;
    11'b00010111111: data <= 32'h3c21b96f;
    11'b00011000000: data <= 32'hb7563492;
    11'b00011000001: data <= 32'hb8533296;
    11'b00011000010: data <= 32'h34f52a26;
    11'b00011000011: data <= 32'h9ce03099;
    11'b00011000100: data <= 32'hbf1ab42e;
    11'b00011000101: data <= 32'hc18cbca2;
    11'b00011000110: data <= 32'hbdf5bcf0;
    11'b00011000111: data <= 32'h390329d3;
    11'b00011001000: data <= 32'h3d183cfb;
    11'b00011001001: data <= 32'h363e3c1b;
    11'b00011001010: data <= 32'hb54834fa;
    11'b00011001011: data <= 32'hb2ec3aa1;
    11'b00011001100: data <= 32'hb0834046;
    11'b00011001101: data <= 32'hb7434004;
    11'b00011001110: data <= 32'hb3a2b05b;
    11'b00011001111: data <= 32'h3ad4c011;
    11'b00011010000: data <= 32'h3e83be9e;
    11'b00011010001: data <= 32'h3cc42ae8;
    11'b00011010010: data <= 32'h38243a3d;
    11'b00011010011: data <= 32'h3aae2ea7;
    11'b00011010100: data <= 32'h3d70b7cf;
    11'b00011010101: data <= 32'h35e2b4f7;
    11'b00011010110: data <= 32'hbf23b500;
    11'b00011010111: data <= 32'hc14abc25;
    11'b00011011000: data <= 32'hbc68be02;
    11'b00011011001: data <= 32'h3afbbb5d;
    11'b00011011010: data <= 32'h3ba2ae5b;
    11'b00011011011: data <= 32'hb6bc1d20;
    11'b00011011100: data <= 32'hbc702bc7;
    11'b00011011101: data <= 32'hb85b3c9d;
    11'b00011011110: data <= 32'hb0c240f1;
    11'b00011011111: data <= 32'hb965401a;
    11'b00011100000: data <= 32'hbc20af79;
    11'b00011100001: data <= 32'hb480be4d;
    11'b00011100010: data <= 32'h3a75b9a3;
    11'b00011100011: data <= 32'h3caf3c11;
    11'b00011100100: data <= 32'h3cb63cf9;
    11'b00011100101: data <= 32'h3e6c2d02;
    11'b00011100110: data <= 32'h3f3ab7d0;
    11'b00011100111: data <= 32'h38d4311e;
    11'b00011101000: data <= 32'hbd4237fa;
    11'b00011101001: data <= 32'hbf04b7f2;
    11'b00011101010: data <= 32'hb107befb;
    11'b00011101011: data <= 32'h3d45bf80;
    11'b00011101100: data <= 32'h3a35bcc9;
    11'b00011101101: data <= 32'hba15b9b9;
    11'b00011101110: data <= 32'hbc44b450;
    11'b00011101111: data <= 32'haeb93a7d;
    11'b00011110000: data <= 32'h303d3f52;
    11'b00011110001: data <= 32'hbc6e3d50;
    11'b00011110010: data <= 32'hc056b66b;
    11'b00011110011: data <= 32'hbe32bcc3;
    11'b00011110100: data <= 32'h9ba6a32d;
    11'b00011110101: data <= 32'h3b523da4;
    11'b00011110110: data <= 32'h3c683ca0;
    11'b00011110111: data <= 32'h3d62a89e;
    11'b00011111000: data <= 32'h3dc4a637;
    11'b00011111001: data <= 32'h38943d30;
    11'b00011111010: data <= 32'hb9cf3f11;
    11'b00011111011: data <= 32'hba6833b9;
    11'b00011111100: data <= 32'h3886bedb;
    11'b00011111101: data <= 32'h3df5c059;
    11'b00011111110: data <= 32'h39aabd7f;
    11'b00011111111: data <= 32'hb729b9d9;
    11'b00100000000: data <= 32'hb065b7c8;
    11'b00100000001: data <= 32'h3bf02d85;
    11'b00100000010: data <= 32'h39873a19;
    11'b00100000011: data <= 32'hbd77376e;
    11'b00100000100: data <= 32'hc1c3b956;
    11'b00100000101: data <= 32'hc050bc29;
    11'b00100000110: data <= 32'hb54da8a1;
    11'b00100000111: data <= 32'h387b3ad9;
    11'b00100001000: data <= 32'h360135dc;
    11'b00100001001: data <= 32'h354cb5ed;
    11'b00100001010: data <= 32'h391137c2;
    11'b00100001011: data <= 32'h364440b4;
    11'b00100001100: data <= 32'hb6034171;
    11'b00100001101: data <= 32'hb76a3a1b;
    11'b00100001110: data <= 32'h372ebd8c;
    11'b00100001111: data <= 32'h3c3ebe86;
    11'b00100010000: data <= 32'h38acb8ac;
    11'b00100010001: data <= 32'h3244b01a;
    11'b00100010010: data <= 32'h3c58b822;
    11'b00100010011: data <= 32'h4044b84f;
    11'b00100010100: data <= 32'h3d152c09;
    11'b00100010101: data <= 32'hbce1320f;
    11'b00100010110: data <= 32'hc164b856;
    11'b00100010111: data <= 32'hbef7bc2e;
    11'b00100011000: data <= 32'ha501b954;
    11'b00100011001: data <= 32'h34bab536;
    11'b00100011010: data <= 32'hb80aba0d;
    11'b00100011011: data <= 32'hb951baf0;
    11'b00100011100: data <= 32'h2d5a38e0;
    11'b00100011101: data <= 32'h35c0413c;
    11'b00100011110: data <= 32'hb5cc4188;
    11'b00100011111: data <= 32'hbb673a20;
    11'b00100100000: data <= 32'hb814bba8;
    11'b00100100001: data <= 32'h3069b8fb;
    11'b00100100010: data <= 32'h349b388a;
    11'b00100100011: data <= 32'h38f33861;
    11'b00100100100: data <= 32'h3f1eb7e9;
    11'b00100100101: data <= 32'h413cb9ec;
    11'b00100100110: data <= 32'h3e2c32cf;
    11'b00100100111: data <= 32'hb9f13a7c;
    11'b00100101000: data <= 32'hbf032da9;
    11'b00100101001: data <= 32'hb915bbf9;
    11'b00100101010: data <= 32'h38fbbd68;
    11'b00100101011: data <= 32'h31c8bd57;
    11'b00100101100: data <= 32'hbc0fbe2f;
    11'b00100101101: data <= 32'hbb6cbd2b;
    11'b00100101110: data <= 32'h351e330c;
    11'b00100101111: data <= 32'h39b03fb4;
    11'b00100110000: data <= 32'hb8073fa8;
    11'b00100110001: data <= 32'hbf1534f0;
    11'b00100110010: data <= 32'hbeb8b920;
    11'b00100110011: data <= 32'hba2932d1;
    11'b00100110100: data <= 32'hafa43d02;
    11'b00100110101: data <= 32'h37373969;
    11'b00100110110: data <= 32'h3de0b93a;
    11'b00100110111: data <= 32'h4051b876;
    11'b00100111000: data <= 32'h3d7f3c30;
    11'b00100111001: data <= 32'hb3073fde;
    11'b00100111010: data <= 32'hb9663b88;
    11'b00100111011: data <= 32'h35d2ba1f;
    11'b00100111100: data <= 32'h3c15be11;
    11'b00100111101: data <= 32'h2e1cbddb;
    11'b00100111110: data <= 32'hbbbbbe0c;
    11'b00100111111: data <= 32'hb4efbdab;
    11'b00101000000: data <= 32'h3d2bb742;
    11'b00101000001: data <= 32'h3d923a00;
    11'b00101000010: data <= 32'hb8333a55;
    11'b00101000011: data <= 32'hc09fb221;
    11'b00101000100: data <= 32'hc078b801;
    11'b00101000101: data <= 32'hbc5e36f6;
    11'b00101000110: data <= 32'hb7023c0c;
    11'b00101000111: data <= 32'hb3fa2745;
    11'b00101001000: data <= 32'h35cbbc6e;
    11'b00101001001: data <= 32'h3c77b4f6;
    11'b00101001010: data <= 32'h3bb03f97;
    11'b00101001011: data <= 32'h2e3e41bd;
    11'b00101001100: data <= 32'haf523dff;
    11'b00101001101: data <= 32'h3884b6a5;
    11'b00101001110: data <= 32'h3a0bbbbd;
    11'b00101001111: data <= 32'hb062b8be;
    11'b00101010000: data <= 32'hb8c9b9a9;
    11'b00101010001: data <= 32'h3980bcea;
    11'b00101010010: data <= 32'h40c2bc1e;
    11'b00101010011: data <= 32'h4017b0d1;
    11'b00101010100: data <= 32'hb4c63249;
    11'b00101010101: data <= 32'hc02bb417;
    11'b00101010110: data <= 32'hbf00b6af;
    11'b00101010111: data <= 32'hb8f22d7e;
    11'b00101011000: data <= 32'hb81a2d06;
    11'b00101011001: data <= 32'hbc4dbc24;
    11'b00101011010: data <= 32'hba84bed6;
    11'b00101011011: data <= 32'h33ffb50f;
    11'b00101011100: data <= 32'h39b8402d;
    11'b00101011101: data <= 32'h317941b5;
    11'b00101011110: data <= 32'hb4c63d89;
    11'b00101011111: data <= 32'hb003b056;
    11'b00101100000: data <= 32'hae2d9e1f;
    11'b00101100001: data <= 32'hb87939c7;
    11'b00101100010: data <= 32'hb59c346a;
    11'b00101100011: data <= 32'h3d1bbbcd;
    11'b00101100100: data <= 32'h41a2bd0c;
    11'b00101100101: data <= 32'h407fb451;
    11'b00101100110: data <= 32'h2cd4383c;
    11'b00101100111: data <= 32'hbcb1348a;
    11'b00101101000: data <= 32'hb7f0b382;
    11'b00101101001: data <= 32'h350eb637;
    11'b00101101010: data <= 32'hb636ba64;
    11'b00101101011: data <= 32'hbe5ebf2c;
    11'b00101101100: data <= 32'hbd57c03b;
    11'b00101101101: data <= 32'h31ccb93c;
    11'b00101101110: data <= 32'h3b953da4;
    11'b00101101111: data <= 32'h311c3f7c;
    11'b00101110000: data <= 32'hbb403945;
    11'b00101110001: data <= 32'hbc8aab13;
    11'b00101110010: data <= 32'hbbda3a8f;
    11'b00101110011: data <= 32'hbbfc3e9d;
    11'b00101110100: data <= 32'hb82c39cb;
    11'b00101110101: data <= 32'h3badbbe2;
    11'b00101110110: data <= 32'h407fbcc6;
    11'b00101110111: data <= 32'h3f6134f9;
    11'b00101111000: data <= 32'h36083e00;
    11'b00101111001: data <= 32'haf4f3c75;
    11'b00101111010: data <= 32'h39ea2c82;
    11'b00101111011: data <= 32'h3c2db7f1;
    11'b00101111100: data <= 32'hb4b9bb32;
    11'b00101111101: data <= 32'hbe8dbeb1;
    11'b00101111110: data <= 32'hbbd2c01a;
    11'b00101111111: data <= 32'h3b89bc88;
    11'b00110000000: data <= 32'h3e65341c;
    11'b00110000001: data <= 32'h33b73830;
    11'b00110000010: data <= 32'hbd5eb1bb;
    11'b00110000011: data <= 32'hbe90af9f;
    11'b00110000100: data <= 32'hbcf93c76;
    11'b00110000101: data <= 32'hbcb83eb9;
    11'b00110000110: data <= 32'hbc423504;
    11'b00110000111: data <= 32'hb011bd93;
    11'b00110001000: data <= 32'h3bf8bc44;
    11'b00110001001: data <= 32'h3c623c12;
    11'b00110001010: data <= 32'h378840a8;
    11'b00110001011: data <= 32'h38023e8b;
    11'b00110001100: data <= 32'h3cdb356d;
    11'b00110001101: data <= 32'h3c2eab88;
    11'b00110001110: data <= 32'hb756a967;
    11'b00110001111: data <= 32'hbd96b972;
    11'b00110010000: data <= 32'hb0febe2b;
    11'b00110010001: data <= 32'h3fbdbde6;
    11'b00110010010: data <= 32'h4077b973;
    11'b00110010011: data <= 32'h3708b597;
    11'b00110010100: data <= 32'hbcb6b850;
    11'b00110010101: data <= 32'hbca3b053;
    11'b00110010110: data <= 32'hb8de3b23;
    11'b00110010111: data <= 32'hbbb23b95;
    11'b00110011000: data <= 32'hbea4b913;
    11'b00110011001: data <= 32'hbd50bff5;
    11'b00110011010: data <= 32'hb0c5bc5c;
    11'b00110011011: data <= 32'h38363ce6;
    11'b00110011100: data <= 32'h3695409e;
    11'b00110011101: data <= 32'h36f63d8f;
    11'b00110011110: data <= 32'h39fc35dd;
    11'b00110011111: data <= 32'h35613985;
    11'b00110100000: data <= 32'hbb083d28;
    11'b00110100001: data <= 32'hbcd2389c;
    11'b00110100010: data <= 32'h3686bb8e;
    11'b00110100011: data <= 32'h40b7be2b;
    11'b00110100100: data <= 32'h40adbb3f;
    11'b00110100101: data <= 32'h38ddb435;
    11'b00110100110: data <= 32'hb73fb1a3;
    11'b00110100111: data <= 32'h2eec28ec;
    11'b00110101000: data <= 32'h38b53807;
    11'b00110101001: data <= 32'hb7c53048;
    11'b00110101010: data <= 32'hbff2bd79;
    11'b00110101011: data <= 32'hbfc2c0a9;
    11'b00110101100: data <= 32'hb7bebd19;
    11'b00110101101: data <= 32'h385a399c;
    11'b00110101110: data <= 32'h35ef3d41;
    11'b00110101111: data <= 32'hac5b36ae;
    11'b00110110000: data <= 32'hb12a2e53;
    11'b00110110001: data <= 32'hb81c3d3d;
    11'b00110110010: data <= 32'hbd23409a;
    11'b00110110011: data <= 32'hbd193d3a;
    11'b00110110100: data <= 32'h32bfb99b;
    11'b00110110101: data <= 32'h3f1fbdab;
    11'b00110110110: data <= 32'h3ed9b708;
    11'b00110110111: data <= 32'h389e3895;
    11'b00110111000: data <= 32'h365838ce;
    11'b00110111001: data <= 32'h3dab355b;
    11'b00110111010: data <= 32'h3e743589;
    11'b00110111011: data <= 32'hae99aa6f;
    11'b00110111100: data <= 32'hbfc6bcfb;
    11'b00110111101: data <= 32'hbeccc027;
    11'b00110111110: data <= 32'h2f03bdcb;
    11'b00110111111: data <= 32'h3c75b3e4;
    11'b00111000000: data <= 32'h3749ae91;
    11'b00111000001: data <= 32'hb811b9cf;
    11'b00111000010: data <= 32'hb9b8b490;
    11'b00111000011: data <= 32'hba393df4;
    11'b00111000100: data <= 32'hbd4640e3;
    11'b00111000101: data <= 32'hbe353c61;
    11'b00111000110: data <= 32'hb975bbf6;
    11'b00111000111: data <= 32'h377bbd2b;
    11'b00111001000: data <= 32'h393e33a0;
    11'b00111001001: data <= 32'h353f3da7;
    11'b00111001010: data <= 32'h3af43c81;
    11'b00111001011: data <= 32'h400437f4;
    11'b00111001100: data <= 32'h3f613885;
    11'b00111001101: data <= 32'haf52390c;
    11'b00111001110: data <= 32'hbec7b27e;
    11'b00111001111: data <= 32'hbb76bd14;
    11'b00111010000: data <= 32'h3c53bdbf;
    11'b00111010001: data <= 32'h3effbc17;
    11'b00111010010: data <= 32'h38adbc60;
    11'b00111010011: data <= 32'hb81cbd66;
    11'b00111010100: data <= 32'hb62bb7ee;
    11'b00111010101: data <= 32'haebc3cf6;
    11'b00111010110: data <= 32'hba9a3f26;
    11'b00111010111: data <= 32'hbf313278;
    11'b00111011000: data <= 32'hbed5be53;
    11'b00111011001: data <= 32'hba5dbd1b;
    11'b00111011010: data <= 32'hb2ae388a;
    11'b00111011011: data <= 32'h27933e16;
    11'b00111011100: data <= 32'h3a0d3ad8;
    11'b00111011101: data <= 32'h3e8b3481;
    11'b00111011110: data <= 32'h3ce93bda;
    11'b00111011111: data <= 32'hb8123f22;
    11'b00111100000: data <= 32'hbdf13cac;
    11'b00111100001: data <= 32'hb49ab5b0;
    11'b00111100010: data <= 32'h3e6ebce4;
    11'b00111100011: data <= 32'h3f62bcb3;
    11'b00111100100: data <= 32'h3863bc77;
    11'b00111100101: data <= 32'haddebc7c;
    11'b00111100110: data <= 32'h39a5b600;
    11'b00111100111: data <= 32'h3ccc3ac4;
    11'b00111101000: data <= 32'ha52f3b6e;
    11'b00111101001: data <= 32'hbf3eb8e8;
    11'b00111101010: data <= 32'hc072bfb8;
    11'b00111101011: data <= 32'hbd03bd30;
    11'b00111101100: data <= 32'hb5eb3500;
    11'b00111101101: data <= 32'hae83398f;
    11'b00111101110: data <= 32'h33feb2dc;
    11'b00111101111: data <= 32'h39b9b505;
    11'b00111110000: data <= 32'h352a3d14;
    11'b00111110001: data <= 32'hbb74415c;
    11'b00111110010: data <= 32'hbdbb4011;
    11'b00111110011: data <= 32'hb40c2f2a;
    11'b00111110100: data <= 32'h3cc4bbb1;
    11'b00111110101: data <= 32'h3c8bb994;
    11'b00111110110: data <= 32'h3278b4cf;
    11'b00111110111: data <= 32'h36b6b525;
    11'b00111111000: data <= 32'h3f8dab92;
    11'b00111111001: data <= 32'h40bc38d4;
    11'b00111111010: data <= 32'h39023868;
    11'b00111111011: data <= 32'hbe58b926;
    11'b00111111100: data <= 32'hbfd4be74;
    11'b00111111101: data <= 32'hb9a8bcb6;
    11'b00111111110: data <= 32'h31e1b4d1;
    11'b00111111111: data <= 32'h9f37b8b4;
    11'b01000000000: data <= 32'hb3ddbe0a;
    11'b01000000001: data <= 32'h1f05bbf8;
    11'b01000000010: data <= 32'had833ce6;
    11'b01000000011: data <= 32'hbb6f4190;
    11'b01000000100: data <= 32'hbdcc3f94;
    11'b01000000101: data <= 32'hba97afc8;
    11'b01000000110: data <= 32'h2473ba99;
    11'b01000000111: data <= 32'haccb2423;
    11'b01000001000: data <= 32'hb5f13945;
    11'b01000001001: data <= 32'h390f355d;
    11'b01000001010: data <= 32'h40d92df5;
    11'b01000001011: data <= 32'h416638d1;
    11'b01000001100: data <= 32'h39cc3b71;
    11'b01000001101: data <= 32'hbd2d3411;
    11'b01000001110: data <= 32'hbca7b947;
    11'b01000001111: data <= 32'h3597ba9e;
    11'b01000010000: data <= 32'h3b74ba51;
    11'b01000010001: data <= 32'h3037be0e;
    11'b01000010010: data <= 32'hb6e1c085;
    11'b01000010011: data <= 32'h2bc6bd78;
    11'b01000010100: data <= 32'h36fb3b2b;
    11'b01000010101: data <= 32'hb4e94033;
    11'b01000010110: data <= 32'hbd6d3b97;
    11'b01000010111: data <= 32'hbe2cba5f;
    11'b01000011000: data <= 32'hbcafbaa2;
    11'b01000011001: data <= 32'hbc5e37cd;
    11'b01000011010: data <= 32'hbb0f3c0e;
    11'b01000011011: data <= 32'h36633303;
    11'b01000011100: data <= 32'h400eb33e;
    11'b01000011101: data <= 32'h40203990;
    11'b01000011110: data <= 32'h345f3f12;
    11'b01000011111: data <= 32'hbc6c3e2a;
    11'b01000100000: data <= 32'hb68136d6;
    11'b01000100001: data <= 32'h3c62b5a8;
    11'b01000100010: data <= 32'h3cbcba3e;
    11'b01000100011: data <= 32'h2527be0c;
    11'b01000100100: data <= 32'hb4e4c01a;
    11'b01000100101: data <= 32'h3ab6bcec;
    11'b01000100110: data <= 32'h3e97381b;
    11'b01000100111: data <= 32'h396f3c9c;
    11'b01000101000: data <= 32'hbc49abb6;
    11'b01000101001: data <= 32'hbf6fbd34;
    11'b01000101010: data <= 32'hbe68ba6b;
    11'b01000101011: data <= 32'hbd413800;
    11'b01000101100: data <= 32'hbc3137de;
    11'b01000101101: data <= 32'haf66b9fb;
    11'b01000101110: data <= 32'h3c27bc02;
    11'b01000101111: data <= 32'h3bf3394d;
    11'b01000110000: data <= 32'hb4d940dd;
    11'b01000110001: data <= 32'hbc2040c0;
    11'b01000110010: data <= 32'hb0533bf5;
    11'b01000110011: data <= 32'h3bca8f90;
    11'b01000110100: data <= 32'h38b8b43c;
    11'b01000110101: data <= 32'hb7efb922;
    11'b01000110110: data <= 32'hb007bc7b;
    11'b01000110111: data <= 32'h3f11ba30;
    11'b01000111000: data <= 32'h41913457;
    11'b01000111001: data <= 32'h3dd9388f;
    11'b01000111010: data <= 32'hb997b5fc;
    11'b01000111011: data <= 32'hbe12bc77;
    11'b01000111100: data <= 32'hbc0db844;
    11'b01000111101: data <= 32'hb95832f2;
    11'b01000111110: data <= 32'hbab3b82d;
    11'b01000111111: data <= 32'hb8cac003;
    11'b01001000000: data <= 32'h30f2bf66;
    11'b01001000001: data <= 32'h350436aa;
    11'b01001000010: data <= 32'hb72f40d9;
    11'b01001000011: data <= 32'hbb684068;
    11'b01001000100: data <= 32'hb62b39b5;
    11'b01001000101: data <= 32'h2d082b5c;
    11'b01001000110: data <= 32'hb8a336fe;
    11'b01001000111: data <= 32'hbd073774;
    11'b01001001000: data <= 32'hb102b2b4;
    11'b01001001001: data <= 32'h4053b755;
    11'b01001001010: data <= 32'h422e31bd;
    11'b01001001011: data <= 32'h3e3c392b;
    11'b01001001100: data <= 32'hb7063394;
    11'b01001001101: data <= 32'hb9ccb2e2;
    11'b01001001110: data <= 32'h316e2468;
    11'b01001001111: data <= 32'h34fb1f2d;
    11'b01001010000: data <= 32'hb83abd1f;
    11'b01001010001: data <= 32'hbabdc17d;
    11'b01001010010: data <= 32'hac9dc089;
    11'b01001010011: data <= 32'h38592c61;
    11'b01001010100: data <= 32'h2e7a3ee5;
    11'b01001010101: data <= 32'hb9143c9a;
    11'b01001010110: data <= 32'hba6bb144;
    11'b01001010111: data <= 32'hbb5aaf42;
    11'b01001011000: data <= 32'hbe613b8d;
    11'b01001011001: data <= 32'hbf743c4e;
    11'b01001011010: data <= 32'hb76da7cd;
    11'b01001011011: data <= 32'h3ee6b974;
    11'b01001011100: data <= 32'h40bb2da8;
    11'b01001011101: data <= 32'h3b823cac;
    11'b01001011110: data <= 32'hb66e3d3f;
    11'b01001011111: data <= 32'h2abd3b00;
    11'b01001100000: data <= 32'h3c9a390b;
    11'b01001100001: data <= 32'h3ade30a1;
    11'b01001100010: data <= 32'hb828bcdc;
    11'b01001100011: data <= 32'hbb07c0f0;
    11'b01001100100: data <= 32'h363ac002;
    11'b01001100101: data <= 32'h3e18b202;
    11'b01001100110: data <= 32'h3c5a3a1c;
    11'b01001100111: data <= 32'hb1a4aca9;
    11'b01001101000: data <= 32'hbb82bbb0;
    11'b01001101001: data <= 32'hbd0cb353;
    11'b01001101010: data <= 32'hbf1a3c5c;
    11'b01001101011: data <= 32'hbfd23aee;
    11'b01001101100: data <= 32'hbb1bba00;
    11'b01001101101: data <= 32'h39c7bdca;
    11'b01001101110: data <= 32'h3c68b06d;
    11'b01001101111: data <= 32'h2d063e73;
    11'b01001110000: data <= 32'hb7cf4012;
    11'b01001110001: data <= 32'h36e93db5;
    11'b01001110010: data <= 32'h3d533bba;
    11'b01001110011: data <= 32'h383638ec;
    11'b01001110100: data <= 32'hbc09b539;
    11'b01001110101: data <= 32'hbb33bd79;
    11'b01001110110: data <= 32'h3c44bd20;
    11'b01001110111: data <= 32'h410eb42a;
    11'b01001111000: data <= 32'h3f802e1e;
    11'b01001111001: data <= 32'h3389b974;
    11'b01001111010: data <= 32'hb8bbbc38;
    11'b01001111011: data <= 32'hb928a0b2;
    11'b01001111100: data <= 32'hbbe73c05;
    11'b01001111101: data <= 32'hbe072fe3;
    11'b01001111110: data <= 32'hbcd0bf71;
    11'b01001111111: data <= 32'hb344c0a1;
    11'b01010000000: data <= 32'h305ab791;
    11'b01010000001: data <= 32'hb5d13e30;
    11'b01010000010: data <= 32'hb7593f49;
    11'b01010000011: data <= 32'h35e83c22;
    11'b01010000100: data <= 32'h39c73a9f;
    11'b01010000101: data <= 32'hb7993ca8;
    11'b01010000110: data <= 32'hbf313aaa;
    11'b01010000111: data <= 32'hbc3eb1eb;
    11'b01010001000: data <= 32'h3d6fb941;
    11'b01010001001: data <= 32'h418fb3d4;
    11'b01010001010: data <= 32'h3f92149b;
    11'b01010001011: data <= 32'h3598b5e6;
    11'b01010001100: data <= 32'h2ce9b582;
    11'b01010001101: data <= 32'h38a9388c;
    11'b01010001110: data <= 32'h33eb3ba9;
    11'b01010001111: data <= 32'hbb14b7da;
    11'b01010010000: data <= 32'hbd40c111;
    11'b01010010001: data <= 32'hb8d5c15f;
    11'b01010010010: data <= 32'h2b9ab9d7;
    11'b01010010011: data <= 32'ha7d73b7b;
    11'b01010010100: data <= 32'hb0e339cd;
    11'b01010010101: data <= 32'h305dad0b;
    11'b01010010110: data <= 32'hae2335a1;
    11'b01010010111: data <= 32'hbda93e14;
    11'b01010011000: data <= 32'hc0c83e4c;
    11'b01010011001: data <= 32'hbd5634e4;
    11'b01010011010: data <= 32'h3bc2b912;
    11'b01010011011: data <= 32'h4006b541;
    11'b01010011100: data <= 32'h3c413544;
    11'b01010011101: data <= 32'h2e7b37f0;
    11'b01010011110: data <= 32'h39953943;
    11'b01010011111: data <= 32'h3eb63ccb;
    11'b01010100000: data <= 32'h3c6f3c76;
    11'b01010100001: data <= 32'hb8d0b6ef;
    11'b01010100010: data <= 32'hbd40c06e;
    11'b01010100011: data <= 32'hb561c07f;
    11'b01010100100: data <= 32'h3a6cb9da;
    11'b01010100101: data <= 32'h3acb3002;
    11'b01010100110: data <= 32'h3578b8cf;
    11'b01010100111: data <= 32'h2c8cbcc1;
    11'b01010101000: data <= 32'hb684abcb;
    11'b01010101001: data <= 32'hbe3a3e67;
    11'b01010101010: data <= 32'hc0b23e33;
    11'b01010101011: data <= 32'hbe2db0ef;
    11'b01010101100: data <= 32'h2e9fbd11;
    11'b01010101101: data <= 32'h393ab8c9;
    11'b01010101110: data <= 32'haea9394a;
    11'b01010101111: data <= 32'hb4c63c99;
    11'b01010110000: data <= 32'h3be23cb0;
    11'b01010110001: data <= 32'h40123dc5;
    11'b01010110010: data <= 32'h3c393db1;
    11'b01010110011: data <= 32'hbb6e356e;
    11'b01010110100: data <= 32'hbd7cbc1d;
    11'b01010110101: data <= 32'h3268bcea;
    11'b01010110110: data <= 32'h3eceb7bb;
    11'b01010110111: data <= 32'h3e64b6e4;
    11'b01010111000: data <= 32'h39a6bd85;
    11'b01010111001: data <= 32'h34fabe54;
    11'b01010111010: data <= 32'h2fd1a8a3;
    11'b01010111011: data <= 32'hb98f3e27;
    11'b01010111100: data <= 32'hbe833bbc;
    11'b01010111101: data <= 32'hbe2cbc81;
    11'b01010111110: data <= 32'hb9c3c02d;
    11'b01010111111: data <= 32'hb79cbb60;
    11'b01011000000: data <= 32'hbaee392d;
    11'b01011000001: data <= 32'hb8003bef;
    11'b01011000010: data <= 32'h3b6739be;
    11'b01011000011: data <= 32'h3e663c45;
    11'b01011000100: data <= 32'h331d3eb5;
    11'b01011000101: data <= 32'hbea53d79;
    11'b01011000110: data <= 32'hbe3234f8;
    11'b01011000111: data <= 32'h37e5b44e;
    11'b01011001000: data <= 32'h3feab278;
    11'b01011001001: data <= 32'h3e43b808;
    11'b01011001010: data <= 32'h3900bcff;
    11'b01011001011: data <= 32'h39bebc48;
    11'b01011001100: data <= 32'h3ce33776;
    11'b01011001101: data <= 32'h397d3e19;
    11'b01011001110: data <= 32'hb94e3649;
    11'b01011001111: data <= 32'hbd6fbf2f;
    11'b01011010000: data <= 32'hbc34c0d9;
    11'b01011010001: data <= 32'hb9eebc1e;
    11'b01011010010: data <= 32'hba223411;
    11'b01011010011: data <= 32'hb4bd2165;
    11'b01011010100: data <= 32'h39e0b83b;
    11'b01011010101: data <= 32'h3adc3410;
    11'b01011010110: data <= 32'hb97f3ee1;
    11'b01011010111: data <= 32'hc0764014;
    11'b01011011000: data <= 32'hbedf3bf4;
    11'b01011011001: data <= 32'h34722606;
    11'b01011011010: data <= 32'h3d3db0b2;
    11'b01011011011: data <= 32'h38f0b2df;
    11'b01011011100: data <= 32'h2b17b7dc;
    11'b01011011101: data <= 32'h3c17b019;
    11'b01011011110: data <= 32'h40773c51;
    11'b01011011111: data <= 32'h3ef73e7e;
    11'b01011100000: data <= 32'hacfe352f;
    11'b01011100001: data <= 32'hbcb6be3f;
    11'b01011100010: data <= 32'hba79bf8a;
    11'b01011100011: data <= 32'hb02ab9e2;
    11'b01011100100: data <= 32'h2511b3f3;
    11'b01011100101: data <= 32'h31c2bce6;
    11'b01011100110: data <= 32'h392dbf56;
    11'b01011100111: data <= 32'h3771b7cd;
    11'b01011101000: data <= 32'hbb2e3e52;
    11'b01011101001: data <= 32'hc037400c;
    11'b01011101010: data <= 32'hbead3981;
    11'b01011101011: data <= 32'hb4cfb7a8;
    11'b01011101100: data <= 32'h2999b626;
    11'b01011101101: data <= 32'hb9f72f17;
    11'b01011101110: data <= 32'hb98a325e;
    11'b01011101111: data <= 32'h3c3b3703;
    11'b01011110000: data <= 32'h412a3d15;
    11'b01011110001: data <= 32'h3f723edd;
    11'b01011110010: data <= 32'hb3773ab1;
    11'b01011110011: data <= 32'hbcb8b77b;
    11'b01011110100: data <= 32'hb4b8b96a;
    11'b01011110101: data <= 32'h3a1fb022;
    11'b01011110110: data <= 32'h3a65b837;
    11'b01011110111: data <= 32'h381ebfec;
    11'b01011111000: data <= 32'h39c6c0d6;
    11'b01011111001: data <= 32'h3a26b96a;
    11'b01011111010: data <= 32'hb0103db8;
    11'b01011111011: data <= 32'hbcdb3ddf;
    11'b01011111100: data <= 32'hbd40b3ea;
    11'b01011111101: data <= 32'hbaa6bd3b;
    11'b01011111110: data <= 32'hbc35b98f;
    11'b01011111111: data <= 32'hbede32e1;
    11'b01100000000: data <= 32'hbc9b3350;
    11'b01100000001: data <= 32'h3afa2cac;
    11'b01100000010: data <= 32'h405839f8;
    11'b01100000011: data <= 32'h3c623e86;
    11'b01100000100: data <= 32'hbb8d3e44;
    11'b01100000101: data <= 32'hbd673aa3;
    11'b01100000110: data <= 32'h2ce5380f;
    11'b01100000111: data <= 32'h3cc43734;
    11'b01100001000: data <= 32'h3ad4b6ff;
    11'b01100001001: data <= 32'h3506bf7e;
    11'b01100001010: data <= 32'h3a91c003;
    11'b01100001011: data <= 32'h3e4fb364;
    11'b01100001100: data <= 32'h3cd13d9f;
    11'b01100001101: data <= 32'ha4903ac8;
    11'b01100001110: data <= 32'hba5cbc1e;
    11'b01100001111: data <= 32'hbbb2bee5;
    11'b01100010000: data <= 32'hbd58b9b4;
    11'b01100010001: data <= 32'hbf012dd2;
    11'b01100010010: data <= 32'hbc2fb7a6;
    11'b01100010011: data <= 32'h3943bc78;
    11'b01100010100: data <= 32'h3da1b4c0;
    11'b01100010101: data <= 32'h2edb3d46;
    11'b01100010110: data <= 32'hbe584004;
    11'b01100010111: data <= 32'hbdd63e1b;
    11'b01100011000: data <= 32'h2d9f3bbf;
    11'b01100011001: data <= 32'h3a33393b;
    11'b01100011010: data <= 32'ha835ae7f;
    11'b01100011011: data <= 32'hb795bc70;
    11'b01100011100: data <= 32'h3a1bbc13;
    11'b01100011101: data <= 32'h40ac371a;
    11'b01100011110: data <= 32'h40883de1;
    11'b01100011111: data <= 32'h3a2338bf;
    11'b01100100000: data <= 32'hb6a0bc19;
    11'b01100100001: data <= 32'hb923bd03;
    11'b01100100010: data <= 32'hb9ddb312;
    11'b01100100011: data <= 32'hbba7ab2f;
    11'b01100100100: data <= 32'hb839bdcc;
    11'b01100100101: data <= 32'h3871c0d9;
    11'b01100100110: data <= 32'h3af3bd0e;
    11'b01100100111: data <= 32'hb4f13b70;
    11'b01100101000: data <= 32'hbe2b3f83;
    11'b01100101001: data <= 32'hbcf53cf1;
    11'b01100101010: data <= 32'hb0dd37ff;
    11'b01100101011: data <= 32'hb3343680;
    11'b01100101100: data <= 32'hbd943368;
    11'b01100101101: data <= 32'hbdddb4f2;
    11'b01100101110: data <= 32'h380fb458;
    11'b01100101111: data <= 32'h411339cc;
    11'b01100110000: data <= 32'h40d13db3;
    11'b01100110001: data <= 32'h39813a57;
    11'b01100110010: data <= 32'hb625b233;
    11'b01100110011: data <= 32'haf65aa8f;
    11'b01100110100: data <= 32'h33c33920;
    11'b01100110101: data <= 32'ha63aa263;
    11'b01100110110: data <= 32'hae37c00f;
    11'b01100110111: data <= 32'h383ac213;
    11'b01100111000: data <= 32'h3b21be4b;
    11'b01100111001: data <= 32'h327e3996;
    11'b01100111010: data <= 32'hb9553d2d;
    11'b01100111011: data <= 32'hb90733d3;
    11'b01100111100: data <= 32'hb570b734;
    11'b01100111101: data <= 32'hbc7f16fe;
    11'b01100111110: data <= 32'hc0ce3679;
    11'b01100111111: data <= 32'hc02da860;
    11'b01101000000: data <= 32'h3216b62c;
    11'b01101000001: data <= 32'h4027338b;
    11'b01101000010: data <= 32'h3e6c3c64;
    11'b01101000011: data <= 32'haee53caf;
    11'b01101000100: data <= 32'hb9163b20;
    11'b01101000101: data <= 32'h34d13cb4;
    11'b01101000110: data <= 32'h3b083db2;
    11'b01101000111: data <= 32'h3450342a;
    11'b01101001000: data <= 32'hb3bfbf66;
    11'b01101001001: data <= 32'h3694c137;
    11'b01101001010: data <= 32'h3d68bc54;
    11'b01101001011: data <= 32'h3d3c39dd;
    11'b01101001100: data <= 32'h38973922;
    11'b01101001101: data <= 32'h3013b9bc;
    11'b01101001110: data <= 32'hb3a7bc5e;
    11'b01101001111: data <= 32'hbd3faddf;
    11'b01101010000: data <= 32'hc0e1376e;
    11'b01101010001: data <= 32'hbfefb683;
    11'b01101010010: data <= 32'h191abd5e;
    11'b01101010011: data <= 32'h3d23bac4;
    11'b01101010100: data <= 32'h37733835;
    11'b01101010101: data <= 32'hbbae3d5b;
    11'b01101010110: data <= 32'hbaae3dde;
    11'b01101010111: data <= 32'h37683ea6;
    11'b01101011000: data <= 32'h3a343eba;
    11'b01101011001: data <= 32'hb60b38e4;
    11'b01101011010: data <= 32'hbc39bc3a;
    11'b01101011011: data <= 32'h2d81bdfb;
    11'b01101011100: data <= 32'h3f3ab2f4;
    11'b01101011101: data <= 32'h40763b2d;
    11'b01101011110: data <= 32'h3d9e3446;
    11'b01101011111: data <= 32'h38f1bc02;
    11'b01101100000: data <= 32'h30a6baea;
    11'b01101100001: data <= 32'hb95e3687;
    11'b01101100010: data <= 32'hbe3238a4;
    11'b01101100011: data <= 32'hbd38bc3c;
    11'b01101100100: data <= 32'h14f2c0fc;
    11'b01101100101: data <= 32'h3939bf7f;
    11'b01101100110: data <= 32'hb305a604;
    11'b01101100111: data <= 32'hbca83c5e;
    11'b01101101000: data <= 32'hb90b3c81;
    11'b01101101001: data <= 32'h37893c83;
    11'b01101101010: data <= 32'h2e8d3d3f;
    11'b01101101011: data <= 32'hbe463ad3;
    11'b01101101100: data <= 32'hc03db1dd;
    11'b01101101101: data <= 32'hb5f9b802;
    11'b01101101110: data <= 32'h3f5f350b;
    11'b01101101111: data <= 32'h409d3b26;
    11'b01101110000: data <= 32'h3d2a33ae;
    11'b01101110001: data <= 32'h389ab7fe;
    11'b01101110010: data <= 32'h38d730e9;
    11'b01101110011: data <= 32'h35d03d60;
    11'b01101110100: data <= 32'hb64f3adf;
    11'b01101110101: data <= 32'hb8fcbdbb;
    11'b01101110110: data <= 32'h2951c20c;
    11'b01101110111: data <= 32'h379bc05c;
    11'b01101111000: data <= 32'ha82db39b;
    11'b01101111001: data <= 32'hb7ca3851;
    11'b01101111010: data <= 32'h2a5f2d3d;
    11'b01101111011: data <= 32'h3851a455;
    11'b01101111100: data <= 32'hb8753958;
    11'b01101111101: data <= 32'hc0f83b82;
    11'b01101111110: data <= 32'hc18a3433;
    11'b01101111111: data <= 32'hb9d6b4bf;
    11'b01110000000: data <= 32'h3d7d2981;
    11'b01110000001: data <= 32'h3dcd381c;
    11'b01110000010: data <= 32'h354a35a5;
    11'b01110000011: data <= 32'h2ec23519;
    11'b01110000100: data <= 32'h3b653d1f;
    11'b01110000101: data <= 32'h3c94405f;
    11'b01110000110: data <= 32'h32a73ce8;
    11'b01110000111: data <= 32'hb842bcca;
    11'b01110001000: data <= 32'hae98c114;
    11'b01110001001: data <= 32'h3961be3a;
    11'b01110001010: data <= 32'h3a4aa463;
    11'b01110001011: data <= 32'h3921a4b5;
    11'b01110001100: data <= 32'h3b1abc03;
    11'b01110001101: data <= 32'h3a4cbba3;
    11'b01110001110: data <= 32'hb930352b;
    11'b01110001111: data <= 32'hc0f03bf8;
    11'b01110010000: data <= 32'hc124307b;
    11'b01110010001: data <= 32'hba2fbb9c;
    11'b01110010010: data <= 32'h3948bb46;
    11'b01110010011: data <= 32'h326ab0e9;
    11'b01110010100: data <= 32'hba6d3547;
    11'b01110010101: data <= 32'hb5ac3a14;
    11'b01110010110: data <= 32'h3c383edb;
    11'b01110010111: data <= 32'h3d1740c8;
    11'b01110011000: data <= 32'hb01f3def;
    11'b01110011001: data <= 32'hbcc8b76c;
    11'b01110011010: data <= 32'hb830bd51;
    11'b01110011011: data <= 32'h3b3db6de;
    11'b01110011100: data <= 32'h3e25368e;
    11'b01110011101: data <= 32'h3dadb56f;
    11'b01110011110: data <= 32'h3d7dbe02;
    11'b01110011111: data <= 32'h3c8abc2c;
    11'b01110100000: data <= 32'ha8ed3930;
    11'b01110100001: data <= 32'hbdf63cc8;
    11'b01110100010: data <= 32'hbe9db451;
    11'b01110100011: data <= 32'hb826bf99;
    11'b01110100100: data <= 32'h2e36bf86;
    11'b01110100101: data <= 32'hb974b9e7;
    11'b01110100110: data <= 32'hbd512ba6;
    11'b01110100111: data <= 32'hb59736a7;
    11'b01110101000: data <= 32'h3c833c6a;
    11'b01110101001: data <= 32'h3acb3f47;
    11'b01110101010: data <= 32'hbc5f3df5;
    11'b01110101011: data <= 32'hc0633552;
    11'b01110101100: data <= 32'hbc33b0e3;
    11'b01110101101: data <= 32'h3ae536e4;
    11'b01110101110: data <= 32'h3e4b390f;
    11'b01110101111: data <= 32'h3cf8b686;
    11'b01110110000: data <= 32'h3caebd00;
    11'b01110110001: data <= 32'h3d92b463;
    11'b01110110010: data <= 32'h3b5d3e08;
    11'b01110110011: data <= 32'hb1673e41;
    11'b01110110100: data <= 32'hb929b824;
    11'b01110110101: data <= 32'hb34fc0b8;
    11'b01110110110: data <= 32'hae18c045;
    11'b01110110111: data <= 32'hb9f3baba;
    11'b01110111000: data <= 32'hbb62b563;
    11'b01110111001: data <= 32'h338db883;
    11'b01110111010: data <= 32'h3d30b222;
    11'b01110111011: data <= 32'h35a53adc;
    11'b01110111100: data <= 32'hbfa23d3c;
    11'b01110111101: data <= 32'hc19b3a24;
    11'b01110111110: data <= 32'hbd6034bc;
    11'b01110111111: data <= 32'h37eb373c;
    11'b01111000000: data <= 32'h3a1b35fa;
    11'b01111000001: data <= 32'h30b1b659;
    11'b01111000010: data <= 32'h3671b8ff;
    11'b01111000011: data <= 32'h3dc539cc;
    11'b01111000100: data <= 32'h3eae40a2;
    11'b01111000101: data <= 32'h395d3faa;
    11'b01111000110: data <= 32'hb39eb557;
    11'b01111000111: data <= 32'hb304bf98;
    11'b01111001000: data <= 32'h211cbd93;
    11'b01111001001: data <= 32'hb07cb5a5;
    11'b01111001010: data <= 32'h2a74b918;
    11'b01111001011: data <= 32'h3c2fbe6d;
    11'b01111001100: data <= 32'h3e4abd6e;
    11'b01111001101: data <= 32'h342f31b7;
    11'b01111001110: data <= 32'hbf933cb6;
    11'b01111001111: data <= 32'hc10439c0;
    11'b01111010000: data <= 32'hbca2b016;
    11'b01111010001: data <= 32'h249cb50a;
    11'b01111010010: data <= 32'hb70fb42f;
    11'b01111010011: data <= 32'hbcd3b7b8;
    11'b01111010100: data <= 32'hb671b36a;
    11'b01111010101: data <= 32'h3d6b3c90;
    11'b01111010110: data <= 32'h3f6640e7;
    11'b01111010111: data <= 32'h389a3ff6;
    11'b01111011000: data <= 32'hb9793251;
    11'b01111011001: data <= 32'hb8bbb9d7;
    11'b01111011010: data <= 32'h30ffab39;
    11'b01111011011: data <= 32'h382636c1;
    11'b01111011100: data <= 32'h3a51b9bb;
    11'b01111011101: data <= 32'h3defc046;
    11'b01111011110: data <= 32'h3f2abec8;
    11'b01111011111: data <= 32'h39ab3413;
    11'b01111100000: data <= 32'hbb9f3d36;
    11'b01111100001: data <= 32'hbd953679;
    11'b01111100010: data <= 32'hb880bb94;
    11'b01111100011: data <= 32'hb4a7bce6;
    11'b01111100100: data <= 32'hbd5bba8f;
    11'b01111100101: data <= 32'hbff4b96b;
    11'b01111100110: data <= 32'hb96eb754;
    11'b01111100111: data <= 32'h3d4a387f;
    11'b01111101000: data <= 32'h3e153ed3;
    11'b01111101001: data <= 32'hb3683eb2;
    11'b01111101010: data <= 32'hbe6239e5;
    11'b01111101011: data <= 32'hbc6a3739;
    11'b01111101100: data <= 32'h30773c43;
    11'b01111101101: data <= 32'h39033ba8;
    11'b01111101110: data <= 32'h3918b92b;
    11'b01111101111: data <= 32'h3c8ebfe4;
    11'b01111110000: data <= 32'h3f0abc6f;
    11'b01111110001: data <= 32'h3dad3bfc;
    11'b01111110010: data <= 32'h35dc3ea4;
    11'b01111110011: data <= 32'hafcb316f;
    11'b01111110100: data <= 32'h2c49bdbd;
    11'b01111110101: data <= 32'hb4fbbdf9;
    11'b01111110110: data <= 32'hbdecba82;
    11'b01111110111: data <= 32'hbf28baa1;
    11'b01111111000: data <= 32'hb3bebcd7;
    11'b01111111001: data <= 32'h3de5b9cd;
    11'b01111111010: data <= 32'h3c4437be;
    11'b01111111011: data <= 32'hbc223c8b;
    11'b01111111100: data <= 32'hc06a3bc4;
    11'b01111111101: data <= 32'hbd493bc2;
    11'b01111111110: data <= 32'ha8273d47;
    11'b01111111111: data <= 32'h232c3b15;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    