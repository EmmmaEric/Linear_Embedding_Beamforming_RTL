
    module interp_rom_3(
    CLK, rst,
    Addr, CEB, Q
    );

    input CLK, rst;
    input [9:0] Addr;
    input CEB;		
    output [20:0] Q;

    (*rom_style = "block" *) reg [20:0] data;

    always @(posedge CLK) begin
    if (rst) begin
        data <= 20'd0;
    end else begin
    if (CEB)
    case(Addr)
            10'b00000000: data <= 20'b00100000000000000000;
        10'b00000001: data <= 20'b00100000000010000000;
        10'b00000010: data <= 20'b00100000000010000000;
        10'b00000011: data <= 20'b00100000000000000000;
        10'b00000100: data <= 20'b00000000000000000000;
        10'b00000101: data <= 20'b00000000000000000000;
        10'b00000110: data <= 20'b00000000000000000000;
        10'b00000111: data <= 20'b00100000000010000000;
        10'b00001000: data <= 20'b00100000000010000000;
        10'b00001001: data <= 20'b00000000000010000000;
        10'b00001010: data <= 20'b00000000000010000000;
        10'b00001011: data <= 20'b00100000000010000000;
        10'b00001100: data <= 20'b00100000000010000000;
        10'b00001101: data <= 20'b00100000000000000000;
        10'b00001110: data <= 20'b00100000000010000000;
        10'b00001111: data <= 20'b00100000000000000000;
        10'b00010000: data <= 20'b00000000000010000000;
        10'b00010001: data <= 20'b00100000000010000000;
        10'b00010010: data <= 20'b00100000000000000000;
        10'b00010011: data <= 20'b00000000000000000000;
        10'b00010100: data <= 20'b00000000000000000000;
        10'b00010101: data <= 20'b00000000000010000000;
        10'b00010110: data <= 20'b00100000000010000000;
        10'b00010111: data <= 20'b00100000000000000000;
        10'b00011000: data <= 20'b00000000000010000000;
        10'b00011001: data <= 20'b00100000000010000000;
        10'b00011010: data <= 20'b00100000000010000000;
        10'b00011011: data <= 20'b00100000000000000000;
        10'b00011100: data <= 20'b00000000000000000000;
        10'b00011101: data <= 20'b00000000000010000000;
        10'b00011110: data <= 20'b00000000000000000000;
        10'b00011111: data <= 20'b00000000000010000000;
        10'b00100000: data <= 20'b00000000000000000000;
        10'b00100001: data <= 20'b00000000000000000000;
        10'b00100010: data <= 20'b00000000000010000000;
        10'b00100011: data <= 20'b00100000000000000000;
        10'b00100100: data <= 20'b00000000000000000000;
        10'b00100101: data <= 20'b00000000000000000000;
        10'b00100110: data <= 20'b00100000000010000000;
        10'b00100111: data <= 20'b00100000000010000000;
        10'b00101000: data <= 20'b00000000000010000000;
        10'b00101001: data <= 20'b00000000000010000000;
        10'b00101010: data <= 20'b00000000000000000000;
        10'b00101011: data <= 20'b00000000000010000000;
        10'b00101100: data <= 20'b00100000000000000000;
        10'b00101101: data <= 20'b00000000000010000000;
        10'b00101110: data <= 20'b00100000000010000000;
        10'b00101111: data <= 20'b00000000010000000001;
        10'b00110000: data <= 20'b00000000000010000000;
        10'b00110001: data <= 20'b00100000000010000000;
        10'b00110010: data <= 20'b00100000000000000000;
        10'b00110011: data <= 20'b00100000000010000000;
        10'b00110100: data <= 20'b00000000000010000000;
        10'b00110101: data <= 20'b00100000000000000000;
        10'b00110110: data <= 20'b00000000000000000000;
        10'b00110111: data <= 20'b00100000000010000000;
        10'b00111000: data <= 20'b00000000000010000000;
        10'b00111001: data <= 20'b00000000000010000000;
        10'b00111010: data <= 20'b00100000000010000000;
        10'b00111011: data <= 20'b00100000000010000000;
        10'b00111100: data <= 20'b00100000000000000000;
        10'b00111101: data <= 20'b00100000000000000000;
        10'b00111110: data <= 20'b00000000000010000000;
        10'b00111111: data <= 20'b00100000000010000000;
        10'b01000000: data <= 20'b00100000000010000000;
        10'b01000001: data <= 20'b00100000000000000000;
        10'b01000010: data <= 20'b00000000000000000000;
        10'b01000011: data <= 20'b00000000000000000000;
        10'b01000100: data <= 20'b00100000000010000000;
        10'b01000101: data <= 20'b00100000000010000000;
        10'b01000110: data <= 20'b00100000000000000000;
        10'b01000111: data <= 20'b00100000000010000000;
        10'b01001000: data <= 20'b00100000000010000000;
        10'b01001001: data <= 20'b00000000000010000000;
        10'b01001010: data <= 20'b00100000000000000000;
        10'b01001011: data <= 20'b00000000000000000000;
        10'b01001100: data <= 20'b00000000000010000001;
        10'b01001101: data <= 20'b00000000000000000000;
        10'b01001110: data <= 20'b00000000000000000000;
        10'b01001111: data <= 20'b00000000000010000000;
        10'b01010000: data <= 20'b00000000000000000000;
        10'b01010001: data <= 20'b00000000000010000000;
        10'b01010010: data <= 20'b00000000000010000000;
        10'b01010011: data <= 20'b00100000000000000000;
        10'b01010100: data <= 20'b00100000000010000000;
        10'b01010101: data <= 20'b00100000000010000000;
        10'b01010110: data <= 20'b00000000000000000000;
        10'b01010111: data <= 20'b00000000000000000000;
        10'b01011000: data <= 20'b00000000000000000000;
        10'b01011001: data <= 20'b00100000000010000000;
        10'b01011010: data <= 20'b00100000000010000000;
        10'b01011011: data <= 20'b00000000000010000000;
        10'b01011100: data <= 20'b00100000000000000000;
        10'b01011101: data <= 20'b00000000000000000000;
        10'b01011110: data <= 20'b00100000000010000000;
        10'b01011111: data <= 20'b00000000000010000000;
        10'b01100000: data <= 20'b00100000000000000000;
        10'b01100001: data <= 20'b00000000000010000000;
        10'b01100010: data <= 20'b00000000000010000000;
        10'b01100011: data <= 20'b00100000000000000000;
        10'b01100100: data <= 20'b00100000000010000000;
        10'b01100101: data <= 20'b00000000000010000000;
        10'b01100110: data <= 20'b00100000010000000000;
        10'b01100111: data <= 20'b00100000000000000001;
        10'b01101000: data <= 20'b00000000000010000000;
        10'b01101001: data <= 20'b00000000000010000000;
        10'b01101010: data <= 20'b00000000000000000000;
        10'b01101011: data <= 20'b00100000000010000000;
        10'b01101100: data <= 20'b00100000000000000000;
        10'b01101101: data <= 20'b00100000000010000000;
        10'b01101110: data <= 20'b00000000000010000000;
        10'b01101111: data <= 20'b00100000000000000000;
        10'b01110000: data <= 20'b00000000000010000000;
        10'b01110001: data <= 20'b00100000000010000000;
        10'b01110010: data <= 20'b00100000000000000000;
        10'b01110011: data <= 20'b00100000000010000000;
        10'b01110100: data <= 20'b00000000000000000000;
        10'b01110101: data <= 20'b00000000000000000000;
        10'b01110110: data <= 20'b00000000000000000000;
        10'b01110111: data <= 20'b00000000000010000000;
        10'b01111000: data <= 20'b00100000000000000000;
        10'b01111001: data <= 20'b00000000000010000000;
        10'b01111010: data <= 20'b00100000000000000000;
        10'b01111011: data <= 20'b00000000000010000000;
        10'b01111100: data <= 20'b00100000000000000000;
        10'b01111101: data <= 20'b00100000000000000000;
        10'b01111110: data <= 20'b00000000000010000000;
        10'b01111111: data <= 20'b00100000000010000000;
        10'b10000000: data <= 20'b00100000000010000000;
        10'b10000001: data <= 20'b00100000000000000000;
        10'b10000010: data <= 20'b00000000000000000000;
        10'b10000011: data <= 20'b00100000000000000000;
        10'b10000100: data <= 20'b00000000010000000000;
        10'b10000101: data <= 20'b00100000000000000000;
        10'b10000110: data <= 20'b00000000000000000000;
        10'b10000111: data <= 20'b00000000000010000000;
        10'b10001000: data <= 20'b00000000000000000000;
        10'b10001001: data <= 20'b00000000000000000000;
        10'b10001010: data <= 20'b00100000000010000000;
        10'b10001011: data <= 20'b00100000000010000000;
        10'b10001100: data <= 20'b00100000010010000000;
        10'b10001101: data <= 20'b00000000000010000000;
        10'b10001110: data <= 20'b00000000000010000000;
        10'b10001111: data <= 20'b00100000000010000000;
        10'b10010000: data <= 20'b00100000000010000000;
        10'b10010001: data <= 20'b00000000000000000000;
        10'b10010010: data <= 20'b00100000000010000000;
        10'b10010011: data <= 20'b00000000000010000000;
        10'b10010100: data <= 20'b00100000000000000000;
        10'b10010101: data <= 20'b00000000000010000000;
        10'b10010110: data <= 20'b00000000000010000000;
        10'b10010111: data <= 20'b00100000000010000000;
        10'b10011000: data <= 20'b00100000000000000000;
        10'b10011001: data <= 20'b00000000000000000000;
        10'b10011010: data <= 20'b00000000000010000000;
        10'b10011011: data <= 20'b00100000000010000000;
        10'b10011100: data <= 20'b00100000000000000000;
        10'b10011101: data <= 20'b00000000000000000000;
        10'b10011110: data <= 20'b00000000000010000000;
        10'b10011111: data <= 20'b00100000000000000000;
        10'b10100000: data <= 20'b00000000000010000000;
        10'b10100001: data <= 20'b00100000000000000000;
        10'b10100010: data <= 20'b00000000000000000000;
        10'b10100011: data <= 20'b00100000000010000000;
        10'b10100100: data <= 20'b00100000000010000000;
        10'b10100101: data <= 20'b00100000000000000000;
        10'b10100110: data <= 20'b00100000000010000000;
        10'b10100111: data <= 20'b00000000000000000000;
        10'b10101000: data <= 20'b00100000000010000000;
        10'b10101001: data <= 20'b00000000000010000000;
        10'b10101010: data <= 20'b00100000000010000000;
        10'b10101011: data <= 20'b00000000000010000000;
        10'b10101100: data <= 20'b00100000000010000000;
        10'b10101101: data <= 20'b00000000000010000000;
        10'b10101110: data <= 20'b00100000000010000000;
        10'b10101111: data <= 20'b00000000000010000000;
        10'b10110000: data <= 20'b00000000010010000000;
        10'b10110001: data <= 20'b00000000000000000000;
        10'b10110010: data <= 20'b00100000000000000000;
        10'b10110011: data <= 20'b00000000000010000000;
        10'b10110100: data <= 20'b00000000000000000000;
        10'b10110101: data <= 20'b00100000000000000000;
        10'b10110110: data <= 20'b00000000000010000000;
        10'b10110111: data <= 20'b00000000000010000000;
        10'b10111000: data <= 20'b00100000000000000000;
        10'b10111001: data <= 20'b00100000000000000000;
        10'b10111010: data <= 20'b00100000000010000010;
        10'b10111011: data <= 20'b00000000000000000000;
        10'b10111100: data <= 20'b00100000000000000000;
        10'b10111101: data <= 20'b00000000000000000000;
        10'b10111110: data <= 20'b00000000000010000000;
        10'b10111111: data <= 20'b00100000000000000000;
        10'b11000000: data <= 20'b00000000000010000000;
        10'b11000001: data <= 20'b00000000000000000000;
        10'b11000010: data <= 20'b00100000000000000000;
        10'b11000011: data <= 20'b00000000000000000000;
        10'b11000100: data <= 20'b00000000000010000000;
        10'b11000101: data <= 20'b00000000000010000000;
        10'b11000110: data <= 20'b00100000000010000000;
        10'b11000111: data <= 20'b00100000000000000000;
        10'b11001000: data <= 20'b00100000000010000000;
        10'b11001001: data <= 20'b00000000000010000000;
        10'b11001010: data <= 20'b00100000000000000000;
        10'b11001011: data <= 20'b00000000000010000000;
        10'b11001100: data <= 20'b00100000000010000000;
        10'b11001101: data <= 20'b00000000000010000000;
        10'b11001110: data <= 20'b00100000000000000000;
        10'b11001111: data <= 20'b00100000000000000000;
        10'b11010000: data <= 20'b00100000000010000000;
        10'b11010001: data <= 20'b00000000000000000001;
        10'b11010010: data <= 20'b00000000000010000000;
        10'b11010011: data <= 20'b00000000000000000000;
        10'b11010100: data <= 20'b00100000000000000000;
        10'b11010101: data <= 20'b00000000000010000000;
        10'b11010110: data <= 20'b00000000000010000000;
        10'b11010111: data <= 20'b00000000000000000000;
        10'b11011000: data <= 20'b00000000000010000000;
        10'b11011001: data <= 20'b00000000000000000000;
        10'b11011010: data <= 20'b00100000000010000000;
        10'b11011011: data <= 20'b00100000000010000000;
        10'b11011100: data <= 20'b00100000000000000000;
        10'b11011101: data <= 20'b00000000000000000000;
        10'b11011110: data <= 20'b00000000000010000000;
        10'b11011111: data <= 20'b00000000000000000000;
        10'b11100000: data <= 20'b00000000000010000000;
        10'b11100001: data <= 20'b00000000000000000000;
        10'b11100010: data <= 20'b00100000000000000000;
        10'b11100011: data <= 20'b00100000000010000000;
        10'b11100100: data <= 20'b00000000000000000000;
        10'b11100101: data <= 20'b00000000000000000000;
        10'b11100110: data <= 20'b00000000000010000000;
        10'b11100111: data <= 20'b00100000000000000000;
        10'b11101000: data <= 20'b00000000000010000000;
        10'b11101001: data <= 20'b00100000000010000000;
        10'b11101010: data <= 20'b00100000000000000000;
        10'b11101011: data <= 20'b00000000000000000000;
        10'b11101100: data <= 20'b00100000000010000000;
        10'b11101101: data <= 20'b00100000000010000000;
        10'b11101110: data <= 20'b00000000000010000001;
        10'b11101111: data <= 20'b00100000000010000000;
        10'b11110000: data <= 20'b00100000000010000000;
        10'b11110001: data <= 20'b00100000000000000000;
        10'b11110010: data <= 20'b00000000000010000000;
        10'b11110011: data <= 20'b00100000000010000000;
        10'b11110100: data <= 20'b00100000000000000000;
        10'b11110101: data <= 20'b00000000000000000000;
        10'b11110110: data <= 20'b00100000000010000000;
        10'b11110111: data <= 20'b00000000000000000000;
        10'b11111000: data <= 20'b00000000100010000000;
        10'b11111001: data <= 20'b00000000000000000000;
        10'b11111010: data <= 20'b00000000000010000000;
        10'b11111011: data <= 20'b00000000000000000000;
        10'b11111100: data <= 20'b00100000000000000000;
        10'b11111101: data <= 20'b00000000000010000000;
        10'b11111110: data <= 20'b00100000000010000000;
        10'b11111111: data <= 20'b00100000000000000000;
        10'b100000000: data <= 20'b00100000000000000000;
        10'b100000001: data <= 20'b00100000000000000000;
        10'b100000010: data <= 20'b00100000000010000000;
        10'b100000011: data <= 20'b00100000000010000000;
        10'b100000100: data <= 20'b00100000000000000000;
        10'b100000101: data <= 20'b00100000000000000000;
        10'b100000110: data <= 20'b00000000000000000000;
        10'b100000111: data <= 20'b00000000000000000000;
        10'b100001000: data <= 20'b00100000000010000000;
        10'b100001001: data <= 20'b00100000000010000000;
        10'b100001010: data <= 20'b00000000000010000000;
        10'b100001011: data <= 20'b00100000000000000000;
        10'b100001100: data <= 20'b00000000000010000000;
        10'b100001101: data <= 20'b00000000000010000000;
        10'b100001110: data <= 20'b00000000000010000000;
        10'b100001111: data <= 20'b00000000000000000000;
        10'b100010000: data <= 20'b00000000000010000000;
        10'b100010001: data <= 20'b00100000000010000000;
        10'b100010010: data <= 20'b00000000000000000000;
        10'b100010011: data <= 20'b00000000000010000000;
        10'b100010100: data <= 20'b00100000010000000000;
        10'b100010101: data <= 20'b00100000000000000000;
        10'b100010110: data <= 20'b00000000000000000000;
        10'b100010111: data <= 20'b00000000000000000000;
        10'b100011000: data <= 20'b00000000000000000000;
        10'b100011001: data <= 20'b00000000000000000000;
        10'b100011010: data <= 20'b00000000000010000000;
        10'b100011011: data <= 20'b00100000000010000000;
        10'b100011100: data <= 20'b00100000000010000000;
        10'b100011101: data <= 20'b00100000000010000000;
        10'b100011110: data <= 20'b00100000000000000000;
        10'b100011111: data <= 20'b00000000000010000000;
        10'b100100000: data <= 20'b00000000000010000000;
        10'b100100001: data <= 20'b00100000000000000000;
        10'b100100010: data <= 20'b00000000000010000000;
        10'b100100011: data <= 20'b00000000000010000000;
        10'b100100100: data <= 20'b00000000000010000000;
        10'b100100101: data <= 20'b00100000010000000001;
        10'b100100110: data <= 20'b00000000000010000000;
        10'b100100111: data <= 20'b00000000000010000000;
        10'b100101000: data <= 20'b00100000000010000000;
        10'b100101001: data <= 20'b00100000000000000000;
        10'b100101010: data <= 20'b00000000000010000000;
        10'b100101011: data <= 20'b00100000000010000000;
        10'b100101100: data <= 20'b00000000000010000000;
        10'b100101101: data <= 20'b00000000000010000000;
        10'b100101110: data <= 20'b00100000000010000000;
        10'b100101111: data <= 20'b00100000000010000000;
        10'b100110000: data <= 20'b00100000000010000000;
        10'b100110001: data <= 20'b00000000000000000000;
        10'b100110010: data <= 20'b00000000000010000000;
        10'b100110011: data <= 20'b00000000000010000000;
        10'b100110100: data <= 20'b00100000000000000000;
        10'b100110101: data <= 20'b00100000000010000000;
        10'b100110110: data <= 20'b00100000000010000000;
        10'b100110111: data <= 20'b00100000000000000000;
        10'b100111000: data <= 20'b00000000000000000000;
        10'b100111001: data <= 20'b00000000000000000000;
        10'b100111010: data <= 20'b00000000000010000000;
        10'b100111011: data <= 20'b00000000000000000000;
        10'b100111100: data <= 20'b00100000000000000000;
        10'b100111101: data <= 20'b00000000000000000000;
        10'b100111110: data <= 20'b00000000000000000000;
        10'b100111111: data <= 20'b00000000000000000000;
        10'b101000000: data <= 20'b00100000000010000000;
        10'b101000001: data <= 20'b00100000000010000000;
        10'b101000010: data <= 20'b00100000000010000000;
        10'b101000011: data <= 20'b00100000000010000000;
        10'b101000100: data <= 20'b00000000000000000000;
        10'b101000101: data <= 20'b00100000000010000000;
        10'b101000110: data <= 20'b00000000000010000000;
        10'b101000111: data <= 20'b00000000000010000000;
        10'b101001000: data <= 20'b00000000000000000000;
        10'b101001001: data <= 20'b00000000000000000000;
        10'b101001010: data <= 20'b00000000000010000000;
        10'b101001011: data <= 20'b00000000000010000000;
        10'b101001100: data <= 20'b00100000000000000000;
        10'b101001101: data <= 20'b00100000000010000001;
        10'b101001110: data <= 20'b00100000000000000000;
        10'b101001111: data <= 20'b00000000000000000000;
        10'b101010000: data <= 20'b00000000000000000000;
        10'b101010001: data <= 20'b00100000000000000000;
        10'b101010010: data <= 20'b00100000000000000000;
        10'b101010011: data <= 20'b00000000000010000000;
        10'b101010100: data <= 20'b00100000000010000000;
        10'b101010101: data <= 20'b00100000000010000000;
        10'b101010110: data <= 20'b00100000000000000000;
        10'b101010111: data <= 20'b00100000000000000000;
        10'b101011000: data <= 20'b00100000000010000000;
        10'b101011001: data <= 20'b00000000000010000000;
        10'b101011010: data <= 20'b00000000000000000000;
        10'b101011011: data <= 20'b00100000000010000000;
        10'b101011100: data <= 20'b00100000000000000000;
        10'b101011101: data <= 20'b00100000000000000000;
        10'b101011110: data <= 20'b00100000000010000000;
        10'b101011111: data <= 20'b00000000010010000000;
        10'b101100000: data <= 20'b00000000000000000000;
        10'b101100001: data <= 20'b00000000000010000000;
        10'b101100010: data <= 20'b00000000000010000000;
        10'b101100011: data <= 20'b00100000000010000000;
        10'b101100100: data <= 20'b00000000000000000000;
        10'b101100101: data <= 20'b00100000000010000000;
        10'b101100110: data <= 20'b00000000000010000000;
        10'b101100111: data <= 20'b00100000000010000000;
        10'b101101000: data <= 20'b00100000000010000000;
        10'b101101001: data <= 20'b00100000000000000000;
        10'b101101010: data <= 20'b00000000000000000000;
        10'b101101011: data <= 20'b00000000000010000000;
        10'b101101100: data <= 20'b00100000000010000000;
        10'b101101101: data <= 20'b00100000000010000001;
        10'b101101110: data <= 20'b00100000000010000000;
        10'b101101111: data <= 20'b00100000000010000000;
        10'b101110000: data <= 20'b00000000000010000000;
        10'b101110001: data <= 20'b00000000000000000000;
        10'b101110010: data <= 20'b00000000000000000000;
        10'b101110011: data <= 20'b00000000000010000000;
        10'b101110100: data <= 20'b00000000000010000000;
        10'b101110101: data <= 20'b00000000000010000000;
        10'b101110110: data <= 20'b00100000000000000000;
        10'b101110111: data <= 20'b00100000000000000000;
        10'b101111000: data <= 20'b00100000000000000000;
        10'b101111001: data <= 20'b00000000000000000000;
        10'b101111010: data <= 20'b00100000000010000000;
        10'b101111011: data <= 20'b00000000000000000000;
        10'b101111100: data <= 20'b00000000000010000000;
        10'b101111101: data <= 20'b00100000000000000000;
        10'b101111110: data <= 20'b00000000000000000000;
        10'b101111111: data <= 20'b00000000000010000000;
        10'b110000000: data <= 20'b00100000000000000000;
        10'b110000001: data <= 20'b00100000000000000000;
        10'b110000010: data <= 20'b00100000000000000000;
        10'b110000011: data <= 20'b00100000000000000000;
        10'b110000100: data <= 20'b00100000000010000000;
        10'b110000101: data <= 20'b00100000000010000000;
        10'b110000110: data <= 20'b00000000000000000000;
        10'b110000111: data <= 20'b00100000000010000000;
        10'b110001000: data <= 20'b00100000000010000000;
        10'b110001001: data <= 20'b00100000000010000000;
        10'b110001010: data <= 20'b00000000000000000000;
        10'b110001011: data <= 20'b00100000000000000000;
        10'b110001100: data <= 20'b00000000000000000000;
        10'b110001101: data <= 20'b00100000000010000000;
        10'b110001110: data <= 20'b00100000000010000000;
        10'b110001111: data <= 20'b00000000000000000000;
        10'b110010000: data <= 20'b00000000000010000000;
        10'b110010001: data <= 20'b00000000000000000000;
        10'b110010010: data <= 20'b00000000000000000000;
        10'b110010011: data <= 20'b00100000000000000000;
        10'b110010100: data <= 20'b00000000000010000000;
        10'b110010101: data <= 20'b00000000000010000000;
        10'b110010110: data <= 20'b00000000000000000000;
        10'b110010111: data <= 20'b00000000000000000000;
        10'b110011000: data <= 20'b00100000000010000000;
        10'b110011001: data <= 20'b00000000000000000000;
        10'b110011010: data <= 20'b00100000000000000000;
        10'b110011011: data <= 20'b00000000000010000000;
        10'b110011100: data <= 20'b00000000000010000001;
        10'b110011101: data <= 20'b00000000000010000000;
        10'b110011110: data <= 20'b00100000000010000000;
        10'b110011111: data <= 20'b00100000000000000000;
        10'b110100000: data <= 20'b00000000000010000000;
        10'b110100001: data <= 20'b00100000000000000000;
        10'b110100010: data <= 20'b00000000000010000000;
        10'b110100011: data <= 20'b00000000000000000000;
        10'b110100100: data <= 20'b00100000000010000000;
        10'b110100101: data <= 20'b00000000000010000000;
        10'b110100110: data <= 20'b00100000000010000000;
        10'b110100111: data <= 20'b00000000000010000000;
        10'b110101000: data <= 20'b00000000000010000000;
        10'b110101001: data <= 20'b00100000000000000000;
        10'b110101010: data <= 20'b00000000000000000000;
        10'b110101011: data <= 20'b00100000000010000000;
        10'b110101100: data <= 20'b00100000000010000000;
        10'b110101101: data <= 20'b00000000000010000000;
        10'b110101110: data <= 20'b00000000000010000000;
        10'b110101111: data <= 20'b00000000000000000000;
        10'b110110000: data <= 20'b00000000000000000000;
        10'b110110001: data <= 20'b00000000000010000000;
        10'b110110010: data <= 20'b00100000000010000000;
        10'b110110011: data <= 20'b00100000000010000000;
        10'b110110100: data <= 20'b00000000000000000000;
        10'b110110101: data <= 20'b00100000000000000000;
        10'b110110110: data <= 20'b00000000000010000000;
        10'b110110111: data <= 20'b00000000000000000000;
        10'b110111000: data <= 20'b00100000000000000000;
        10'b110111001: data <= 20'b00000000000000000000;
        10'b110111010: data <= 20'b00000000000010000000;
        10'b110111011: data <= 20'b00100000000000000000;
        10'b110111100: data <= 20'b00100000000000000000;
        10'b110111101: data <= 20'b00000000000010000000;
        10'b110111110: data <= 20'b00100000000000000000;
        10'b110111111: data <= 20'b00000000000010000000;
        10'b111000000: data <= 20'b00000000000000000000;
        10'b111000001: data <= 20'b00000000000000000000;
        10'b111000010: data <= 20'b00100000000010000000;
        10'b111000011: data <= 20'b00100000000000000000;
        10'b111000100: data <= 20'b00000000000000000000;
        10'b111000101: data <= 20'b00100000000000000000;
        10'b111000110: data <= 20'b00100000000010000000;
        10'b111000111: data <= 20'b00100000000010000000;
        10'b111001000: data <= 20'b00000000000010000000;
        10'b111001001: data <= 20'b00000000000000000000;
        10'b111001010: data <= 20'b00000000000000000000;
        10'b111001011: data <= 20'b00000000000000000000;
        10'b111001100: data <= 20'b00100000000000000001;
        10'b111001101: data <= 20'b00100000000010000000;
        10'b111001110: data <= 20'b00000000000010000000;
        10'b111001111: data <= 20'b00000000000010000000;
        10'b111010000: data <= 20'b00000000000010000000;
        10'b111010001: data <= 20'b00100000000010000000;
        10'b111010010: data <= 20'b00100000000000000000;
        10'b111010011: data <= 20'b00000000000000000000;
        10'b111010100: data <= 20'b00100000000000000000;
        10'b111010101: data <= 20'b00000000000010000000;
        10'b111010110: data <= 20'b00000000000010000000;
        10'b111010111: data <= 20'b00100000000000000000;
        10'b111011000: data <= 20'b00100000000010000000;
        10'b111011001: data <= 20'b00100000000010000000;
        10'b111011010: data <= 20'b00100000000000000000;
        10'b111011011: data <= 20'b00000000000000000000;
        10'b111011100: data <= 20'b00100000000010000000;
        10'b111011101: data <= 20'b00000000000000000000;
        10'b111011110: data <= 20'b00000000000000000000;
        10'b111011111: data <= 20'b00100000000000000000;
        10'b111100000: data <= 20'b00000000000010000000;
        10'b111100001: data <= 20'b00100001010010000000;
        10'b111100010: data <= 20'b00100000000010000000;
        10'b111100011: data <= 20'b00100000000010000000;
        10'b111100100: data <= 20'b00100000000000000000;
        10'b111100101: data <= 20'b00100000000010000000;
        10'b111100110: data <= 20'b00100000000000000000;
        10'b111100111: data <= 20'b00000000000000000000;
        10'b111101000: data <= 20'b00000000000010000000;
        10'b111101001: data <= 20'b00000000000010000000;
        10'b111101010: data <= 20'b00100000000010000000;
        10'b111101011: data <= 20'b00100000000000000000;
        10'b111101100: data <= 20'b00000000000010000000;
        10'b111101101: data <= 20'b00100000000010000000;
        10'b111101110: data <= 20'b00000000000010000000;
        10'b111101111: data <= 20'b00100000000000000000;
        10'b111110000: data <= 20'b00000000000010000000;
        10'b111110001: data <= 20'b00100000000010000000;
        10'b111110010: data <= 20'b00000000000000000000;
        10'b111110011: data <= 20'b00100000000010000000;
        10'b111110100: data <= 20'b00000000000000000000;
        10'b111110101: data <= 20'b00100000000000000000;
        10'b111110110: data <= 20'b00100000000010000000;
        10'b111110111: data <= 20'b00000000000010000000;
        10'b111111000: data <= 20'b00000000000000000000;
        10'b111111001: data <= 20'b00100000000000000000;
        10'b111111010: data <= 20'b00000000000000000000;
        10'b111111011: data <= 20'b00100000000000000000;
        10'b111111100: data <= 20'b00000000000000000000;
        10'b111111101: data <= 20'b00000000000000000000;
        10'b111111110: data <= 20'b00100000000010000000;
        10'b111111111: data <= 20'b00100000000000000000;
        10'b1000000000: data <= 20'b00000000000000000000;
        10'b1000000001: data <= 20'b00000000000000000000;
        10'b1000000010: data <= 20'b00000000000010000000;
        10'b1000000011: data <= 20'b00100000000010000000;
        10'b1000000100: data <= 20'b00100000000010000000;
        10'b1000000101: data <= 20'b00000000000000000000;
        10'b1000000110: data <= 20'b00000000000000000000;
        10'b1000000111: data <= 20'b00100000100000000000;
        10'b1000001000: data <= 20'b00100000000000000000;
        10'b1000001001: data <= 20'b00000000000010000000;
        10'b1000001010: data <= 20'b00100000000010000000;
        10'b1000001011: data <= 20'b00000000000000000000;
        10'b1000001100: data <= 20'b00100000000000000000;
        10'b1000001101: data <= 20'b00100000000000000000;
        10'b1000001110: data <= 20'b00000000000010000000;
        10'b1000001111: data <= 20'b00100000000010000000;
        10'b1000010000: data <= 20'b00000000000010000000;
        10'b1000010001: data <= 20'b00100000000010000000;
        10'b1000010010: data <= 20'b00000000000000000000;
        10'b1000010011: data <= 20'b00100000000000000000;
        10'b1000010100: data <= 20'b00100000000000000000;
        10'b1000010101: data <= 20'b00000000000000000000;
        10'b1000010110: data <= 20'b00000000000000000000;
        10'b1000010111: data <= 20'b00000000000000000000;
        10'b1000011000: data <= 20'b00000000000010000000;
        10'b1000011001: data <= 20'b00000000000000000000;
        10'b1000011010: data <= 20'b00000000000000000000;
        10'b1000011011: data <= 20'b00100000000010000000;
        10'b1000011100: data <= 20'b00100000010010000001;
        10'b1000011101: data <= 20'b00000000000000000000;
        10'b1000011110: data <= 20'b00100000000000000000;
        10'b1000011111: data <= 20'b00000000000000000000;
        10'b1000100000: data <= 20'b00000000000010000000;
        10'b1000100001: data <= 20'b00100000000010000000;
        10'b1000100010: data <= 20'b00000000000000000000;
        10'b1000100011: data <= 20'b00000000010010000001;
        10'b1000100100: data <= 20'b00000000000000000000;
        10'b1000100101: data <= 20'b00100000000010000000;
        10'b1000100110: data <= 20'b00000000000010000000;
        10'b1000100111: data <= 20'b00100000000010000000;
        10'b1000101000: data <= 20'b00100000000010000000;
        10'b1000101001: data <= 20'b00100000000010000000;
        10'b1000101010: data <= 20'b00000000000000000000;
        10'b1000101011: data <= 20'b00000000000010000000;
        10'b1000101100: data <= 20'b00000000000010000000;
        10'b1000101101: data <= 20'b00100000000000000000;
        10'b1000101110: data <= 20'b00000000000000000000;
        10'b1000101111: data <= 20'b00100000000010000000;
        10'b1000110000: data <= 20'b00000000000010000000;
        10'b1000110001: data <= 20'b00000000000000000000;
        10'b1000110010: data <= 20'b00000000000000000000;
        10'b1000110011: data <= 20'b00000000000000000000;
        10'b1000110100: data <= 20'b00000000000000000000;
        10'b1000110101: data <= 20'b00000000000000000000;
        10'b1000110110: data <= 20'b00000000000010000000;
        10'b1000110111: data <= 20'b00100000000010000000;
        10'b1000111000: data <= 20'b00100000000000000000;
        10'b1000111001: data <= 20'b00000000000010000000;
        10'b1000111010: data <= 20'b00100000000010000000;
        10'b1000111011: data <= 20'b00100000000000000000;
        10'b1000111100: data <= 20'b00000000000000000000;
        10'b1000111101: data <= 20'b00000000000010000000;
        10'b1000111110: data <= 20'b00000000000000000000;
        10'b1000111111: data <= 20'b00000000000010000000;
        10'b1001000000: data <= 20'b00100000000010000000;
        10'b1001000001: data <= 20'b00000000000000000000;
        10'b1001000010: data <= 20'b00000000000010000000;
        10'b1001000011: data <= 20'b00000000000010000000;
        10'b1001000100: data <= 20'b00100000000000000000;
        10'b1001000101: data <= 20'b00100000000010000000;
        10'b1001000110: data <= 20'b00000000000000000000;
        10'b1001000111: data <= 20'b00100000000000000000;
        10'b1001001000: data <= 20'b00000000000000000000;
        10'b1001001001: data <= 20'b00100000000010000000;
        10'b1001001010: data <= 20'b00100000000000000000;
        10'b1001001011: data <= 20'b00000000000010000000;
        10'b1001001100: data <= 20'b00000000000010000000;
        10'b1001001101: data <= 20'b00100000000000000000;
        10'b1001001110: data <= 20'b00000000000000000000;
        10'b1001001111: data <= 20'b00000000000000000000;
        10'b1001010000: data <= 20'b00000000000000000000;
        10'b1001010001: data <= 20'b00000000000000000000;
        10'b1001010010: data <= 20'b00000000000010000000;
        10'b1001010011: data <= 20'b00000000000010000000;
        10'b1001010100: data <= 20'b00100000000000000000;
        10'b1001010101: data <= 20'b00100000000000000000;
        10'b1001010110: data <= 20'b00100000000010000000;
        10'b1001010111: data <= 20'b00000000000010000000;
        10'b1001011000: data <= 20'b00100000000000000000;
        10'b1001011001: data <= 20'b00100000000010000000;
        10'b1001011010: data <= 20'b00000000000010000000;
        10'b1001011011: data <= 20'b00100000000000000000;
        10'b1001011100: data <= 20'b00000000000010000000;
        10'b1001011101: data <= 20'b00100000000010000000;
        10'b1001011110: data <= 20'b00000000000000000000;
        10'b1001011111: data <= 20'b00100000000010000000;
        10'b1001100000: data <= 20'b00000000000010000000;
        10'b1001100001: data <= 20'b00100000000010000000;
        10'b1001100010: data <= 20'b00100000000000000000;
        10'b1001100011: data <= 20'b00100000000000000000;
        10'b1001100100: data <= 20'b00000000000000000000;
        10'b1001100101: data <= 20'b00000000000000000000;
        10'b1001100110: data <= 20'b00000000000000000000;
        10'b1001100111: data <= 20'b00000000000000000000;
        10'b1001101000: data <= 20'b00100000000010000000;
        10'b1001101001: data <= 20'b00100000000010000000;
        10'b1001101010: data <= 20'b00100000000000000000;
        10'b1001101011: data <= 20'b00000000000010000000;
        10'b1001101100: data <= 20'b00100000000000000000;
        10'b1001101101: data <= 20'b00100000000010000000;
        10'b1001101110: data <= 20'b00000000000010000000;
        10'b1001101111: data <= 20'b00100000000000000000;
        10'b1001110000: data <= 20'b00100000000010000000;
        10'b1001110001: data <= 20'b00100000000000000000;
        10'b1001110010: data <= 20'b00100000000000000000;
        10'b1001110011: data <= 20'b00000000000000000000;
        10'b1001110100: data <= 20'b00100000000010000000;
        10'b1001110101: data <= 20'b00000000000000000000;
        10'b1001110110: data <= 20'b00100000000010000000;
        10'b1001110111: data <= 20'b00100000000000000000;
        10'b1001111000: data <= 20'b00100000000000000000;
        10'b1001111001: data <= 20'b00000000000000000000;
        10'b1001111010: data <= 20'b00100000000000000000;
        10'b1001111011: data <= 20'b00000000000000000000;
        10'b1001111100: data <= 20'b00100000000010000000;
        10'b1001111101: data <= 20'b00000000000000000000;
        10'b1001111110: data <= 20'b00100000000000000000;
        10'b1001111111: data <= 20'b00000000000000000000;
        10'b1010000000: data <= 20'b00100000000000000000;
        10'b1010000001: data <= 20'b00100000000010000000;
        10'b1010000010: data <= 20'b00100000000010000000;
        10'b1010000011: data <= 20'b00100000000010000000;
        10'b1010000100: data <= 20'b00100000000000000000;
        10'b1010000101: data <= 20'b00100000000000000000;
        10'b1010000110: data <= 20'b00000000000010000000;
        10'b1010000111: data <= 20'b00100000000010000000;
        10'b1010001000: data <= 20'b00000000000010000000;
        10'b1010001001: data <= 20'b00100000000000000000;
        10'b1010001010: data <= 20'b00000000000000000000;
        10'b1010001011: data <= 20'b00100000000010000000;
        10'b1010001100: data <= 20'b00100000000010000000;
        10'b1010001101: data <= 20'b00100000000010000000;
        10'b1010001110: data <= 20'b00100000000000000000;
        10'b1010001111: data <= 20'b00000000000000000000;
        10'b1010010000: data <= 20'b00100000000010000000;
        10'b1010010001: data <= 20'b00100000000000000000;
        10'b1010010010: data <= 20'b00000000000000000000;
        10'b1010010011: data <= 20'b00100000000000000000;
        10'b1010010100: data <= 20'b00100000000000000000;
        10'b1010010101: data <= 20'b00100000110000000010;
        10'b1010010110: data <= 20'b00000000000010000000;
        10'b1010010111: data <= 20'b00100000000000000000;
        10'b1010011000: data <= 20'b00000000000000000000;
        10'b1010011001: data <= 20'b00000000000010000000;
        10'b1010011010: data <= 20'b00000000010010000000;
        10'b1010011011: data <= 20'b00000000000000000000;
        10'b1010011100: data <= 20'b00100000000010000000;
        10'b1010011101: data <= 20'b00100000000000000000;
        10'b1010011110: data <= 20'b00000000000010000000;
        10'b1010011111: data <= 20'b00100000000000000000;
        10'b1010100000: data <= 20'b00100000000010000000;
        10'b1010100001: data <= 20'b00000000000010000000;
        10'b1010100010: data <= 20'b00100000000000000000;
        10'b1010100011: data <= 20'b00100000000010000000;
        10'b1010100100: data <= 20'b00000000000000000000;
        10'b1010100101: data <= 20'b00000000000000000000;
        10'b1010100110: data <= 20'b00100000000000000000;
        10'b1010100111: data <= 20'b00000000000010000000;
        10'b1010101000: data <= 20'b00100000000000000000;
        10'b1010101001: data <= 20'b00100000000000000000;
        10'b1010101010: data <= 20'b00100000000000000000;
        10'b1010101011: data <= 20'b00100000010000000000;
        10'b1010101100: data <= 20'b00000000000010000000;
        10'b1010101101: data <= 20'b00000000000010000000;
        10'b1010101110: data <= 20'b00000000000010000000;
        10'b1010101111: data <= 20'b00100000000000000000;
        10'b1010110000: data <= 20'b00100000000010000000;
        10'b1010110001: data <= 20'b00100000000010000000;
        10'b1010110010: data <= 20'b00100000000010000000;
        10'b1010110011: data <= 20'b00000000000010000000;
        10'b1010110100: data <= 20'b00000000000010000000;
        10'b1010110101: data <= 20'b00100000000010000000;
        10'b1010110110: data <= 20'b00100000000010000000;
        10'b1010110111: data <= 20'b00000000000010000000;
        10'b1010111000: data <= 20'b00000000000000000000;
        10'b1010111001: data <= 20'b00000000000000000000;
        10'b1010111010: data <= 20'b00100000000010000000;
        10'b1010111011: data <= 20'b00000000000010000000;
        10'b1010111100: data <= 20'b00100000000010000000;
        10'b1010111101: data <= 20'b00000000000000000000;
        10'b1010111110: data <= 20'b00100000000000000000;
        10'b1010111111: data <= 20'b00000000000000000000;
        10'b1011000000: data <= 20'b00000000000000000000;
        10'b1011000001: data <= 20'b00000000000010000000;
        10'b1011000010: data <= 20'b00000000000010000000;
        10'b1011000011: data <= 20'b00100000000000000000;
        10'b1011000100: data <= 20'b00000000000010000000;
        10'b1011000101: data <= 20'b00000000000010000000;
        10'b1011000110: data <= 20'b00000000000010000000;
        10'b1011000111: data <= 20'b00100000000000000000;
        10'b1011001000: data <= 20'b00100000000010000000;
        10'b1011001001: data <= 20'b00000000000010000000;
        10'b1011001010: data <= 20'b00000000000000000000;
        10'b1011001011: data <= 20'b00100000000000000000;
        10'b1011001100: data <= 20'b00000000000000000000;
        10'b1011001101: data <= 20'b00000000000010000000;
        10'b1011001110: data <= 20'b00000000000010000000;
        10'b1011001111: data <= 20'b00100000000000000000;
        10'b1011010000: data <= 20'b00100000000010000000;
        10'b1011010001: data <= 20'b00000000000010000000;
        10'b1011010010: data <= 20'b00100000000010000000;
        10'b1011010011: data <= 20'b00000000000000000000;
        10'b1011010100: data <= 20'b00100000000010000000;
        10'b1011010101: data <= 20'b00000000000010000000;
        10'b1011010110: data <= 20'b00000000000000000000;
        10'b1011010111: data <= 20'b00000000000010000000;
        10'b1011011000: data <= 20'b00100000000000000000;
        10'b1011011001: data <= 20'b00000000000010000000;
        10'b1011011010: data <= 20'b00100000000010000000;
        10'b1011011011: data <= 20'b00000000000010000000;
        10'b1011011100: data <= 20'b00100000000010000000;
        10'b1011011101: data <= 20'b00000000000000000000;
        10'b1011011110: data <= 20'b00000000000000000000;
        10'b1011011111: data <= 20'b00100000000010000000;
        10'b1011100000: data <= 20'b00100000000010000000;
        10'b1011100001: data <= 20'b00000000000010000000;
        10'b1011100010: data <= 20'b00100000000010000000;
        10'b1011100011: data <= 20'b00000000000000000000;
        10'b1011100100: data <= 20'b00000000000010000000;
        10'b1011100101: data <= 20'b00100000000000000000;
        10'b1011100110: data <= 20'b00000000000000000000;
        10'b1011100111: data <= 20'b00000000000010000000;
        10'b1011101000: data <= 20'b00100000000010000000;
        10'b1011101001: data <= 20'b00100000000010000000;
        10'b1011101010: data <= 20'b00000000000010000000;
        10'b1011101011: data <= 20'b00000000000000000000;
        10'b1011101100: data <= 20'b00000000000010000000;
        10'b1011101101: data <= 20'b00000000000000000000;
        10'b1011101110: data <= 20'b00000000000000000000;
        10'b1011101111: data <= 20'b00100000000000000000;
        10'b1011110000: data <= 20'b00000000000000000000;
        10'b1011110001: data <= 20'b00100000000000000000;
        10'b1011110010: data <= 20'b00100000010010000000;
        10'b1011110011: data <= 20'b00000000000010000000;
        10'b1011110100: data <= 20'b00100000000010000000;
        10'b1011110101: data <= 20'b00000000000010000000;
        10'b1011110110: data <= 20'b00000000000000000000;
        10'b1011110111: data <= 20'b00000000000010000000;
        10'b1011111000: data <= 20'b00100000000000000000;
        10'b1011111001: data <= 20'b00000000000000000000;
        10'b1011111010: data <= 20'b00100000000000000000;
        10'b1011111011: data <= 20'b00000000000000000000;
        10'b1011111100: data <= 20'b00100000000010000000;
        10'b1011111101: data <= 20'b00000000000000000000;
        10'b1011111110: data <= 20'b00000000000000000000;
        10'b1011111111: data <= 20'b00100000000000000000;
        10'b1100000000: data <= 20'b00100000000000000000;
        10'b1100000001: data <= 20'b00100000000010000000;
        10'b1100000010: data <= 20'b00000000000000000000;
        10'b1100000011: data <= 20'b00100000000010000000;
        10'b1100000100: data <= 20'b00100000000000000000;
        10'b1100000101: data <= 20'b00100000000000000000;
        10'b1100000110: data <= 20'b00000000000010000000;
        10'b1100000111: data <= 20'b00000000000010000000;
        10'b1100001000: data <= 20'b00000000000000000000;
        10'b1100001001: data <= 20'b00100000000000000000;
        10'b1100001010: data <= 20'b00000000000010000000;
        10'b1100001011: data <= 20'b00000000000000000000;
        10'b1100001100: data <= 20'b00000000000010000000;
        10'b1100001101: data <= 20'b00000000000000000000;
        10'b1100001110: data <= 20'b00100000000010000000;
        10'b1100001111: data <= 20'b00000000000010000000;
        10'b1100010000: data <= 20'b00100000000000000000;
        10'b1100010001: data <= 20'b00100000000010000000;
        10'b1100010010: data <= 20'b00000000000000000000;
        10'b1100010011: data <= 20'b00000000000000000000;
        10'b1100010100: data <= 20'b00100000000010000000;
        10'b1100010101: data <= 20'b00000000000010000000;
        10'b1100010110: data <= 20'b00100000000000000000;
        10'b1100010111: data <= 20'b00100000000010000000;
        10'b1100011000: data <= 20'b00100000000010000000;
        10'b1100011001: data <= 20'b00000000000010000000;
        10'b1100011010: data <= 20'b00000000000010000000;
        10'b1100011011: data <= 20'b00100000000010000000;
        10'b1100011100: data <= 20'b00000000000000000000;
        10'b1100011101: data <= 20'b00000000000000000000;
        10'b1100011110: data <= 20'b00000000000000000000;
        10'b1100011111: data <= 20'b00000000000010000000;
        10'b1100100000: data <= 20'b00100000000000000000;
        10'b1100100001: data <= 20'b00100000000000000000;
        10'b1100100010: data <= 20'b00100000000010000000;
        10'b1100100011: data <= 20'b00000000000010000000;
        10'b1100100100: data <= 20'b00000000000010000000;
        10'b1100100101: data <= 20'b00000000000000000000;
        10'b1100100110: data <= 20'b00000000000000000000;
        10'b1100100111: data <= 20'b00000000000000000000;
        10'b1100101000: data <= 20'b00100000000000000000;
        10'b1100101001: data <= 20'b00000000000010000000;
        10'b1100101010: data <= 20'b00000000000000000000;
        10'b1100101011: data <= 20'b00100000000000000000;
        10'b1100101100: data <= 20'b00100000000010000000;
        10'b1100101101: data <= 20'b00100000000010000000;
        10'b1100101110: data <= 20'b00100000000010000000;
        10'b1100101111: data <= 20'b00100000000000000000;
        10'b1100110000: data <= 20'b00000000000010000000;
        10'b1100110001: data <= 20'b00100000000000000000;
        10'b1100110010: data <= 20'b00100000000000000000;
        10'b1100110011: data <= 20'b00100000000010000000;
        10'b1100110100: data <= 20'b00000000000010000000;
        10'b1100110101: data <= 20'b00000000000010000000;
        10'b1100110110: data <= 20'b00100000000000000000;
        10'b1100110111: data <= 20'b00100000000010000000;
        10'b1100111000: data <= 20'b00000000000010000000;
        10'b1100111001: data <= 20'b00100000000010000000;
        10'b1100111010: data <= 20'b00000000000010000000;
        10'b1100111011: data <= 20'b00100000000010000000;
        10'b1100111100: data <= 20'b00000000000010000000;
        10'b1100111101: data <= 20'b00000000000010000000;
        10'b1100111110: data <= 20'b00100000000000000000;
        10'b1100111111: data <= 20'b00000000000010000000;
        10'b1101000000: data <= 20'b00000000000000000000;
        10'b1101000001: data <= 20'b00000000000010000000;
        10'b1101000010: data <= 20'b00000000000010000000;
        10'b1101000011: data <= 20'b00000000000010000000;
        10'b1101000100: data <= 20'b00000000000010000000;
        10'b1101000101: data <= 20'b00100000000010000000;
        10'b1101000110: data <= 20'b00000000000010000000;
        10'b1101000111: data <= 20'b00100000000010000000;
        10'b1101001000: data <= 20'b00100000000010000000;
        10'b1101001001: data <= 20'b00000000000000000000;
        10'b1101001010: data <= 20'b00100000000010000000;
        10'b1101001011: data <= 20'b00000000000000000000;
        10'b1101001100: data <= 20'b00100000000010000000;
        10'b1101001101: data <= 20'b00100000000000000000;
        10'b1101001110: data <= 20'b00100000000010000000;
        10'b1101001111: data <= 20'b00100000000010000000;
        10'b1101010000: data <= 20'b00100000000000000000;
        10'b1101010001: data <= 20'b00000000000010000000;
        10'b1101010010: data <= 20'b00000000000010000000;
        10'b1101010011: data <= 20'b00100000000000000000;
        10'b1101010100: data <= 20'b00100000000010000000;
        10'b1101010101: data <= 20'b00000000000000000000;
        10'b1101010110: data <= 20'b00100000000010000000;
        10'b1101010111: data <= 20'b00100000000010000000;
        10'b1101011000: data <= 20'b00000000000000000000;
        10'b1101011001: data <= 20'b00000000000010000000;
        10'b1101011010: data <= 20'b00100000000010000000;
        10'b1101011011: data <= 20'b00100000000010000000;
        10'b1101011100: data <= 20'b00000000000010000000;
        10'b1101011101: data <= 20'b00000000000000000000;
        10'b1101011110: data <= 20'b00100000000010000000;
        10'b1101011111: data <= 20'b00100000000010000000;
        10'b1101100000: data <= 20'b00000000000000000000;
        10'b1101100001: data <= 20'b00000000000000000000;
        10'b1101100010: data <= 20'b00000000000010000000;
        10'b1101100011: data <= 20'b00000000000010000000;
        10'b1101100100: data <= 20'b00000000000000000000;
        10'b1101100101: data <= 20'b00000000000010000000;
        10'b1101100110: data <= 20'b00000000000000000000;
        10'b1101100111: data <= 20'b00100000000000000000;
        10'b1101101000: data <= 20'b00000000010010000000;
        10'b1101101001: data <= 20'b00100000000000000000;
        10'b1101101010: data <= 20'b00000000000000000000;
        10'b1101101011: data <= 20'b00100000000000000000;
        10'b1101101100: data <= 20'b00000000000010000000;
        10'b1101101101: data <= 20'b00000000000010000000;
        10'b1101101110: data <= 20'b00100000000010000000;
        10'b1101101111: data <= 20'b00100000000010000000;
        10'b1101110000: data <= 20'b00100000000010000000;
        10'b1101110001: data <= 20'b00000000000000000000;
        10'b1101110010: data <= 20'b00000000000010000000;
        10'b1101110011: data <= 20'b00100000000000000000;
        10'b1101110100: data <= 20'b00100000000000000000;
        10'b1101110101: data <= 20'b00100000000010000000;
        10'b1101110110: data <= 20'b00100000000010000000;
        10'b1101110111: data <= 20'b00100000000000000000;
        10'b1101111000: data <= 20'b00100000000000000000;
        10'b1101111001: data <= 20'b00000000000010000000;
        10'b1101111010: data <= 20'b00000000010010000001;
        10'b1101111011: data <= 20'b00000000000010000000;
        10'b1101111100: data <= 20'b00100000000010000000;
        10'b1101111101: data <= 20'b00000000000000000000;
        10'b1101111110: data <= 20'b00000000000000000000;
        10'b1101111111: data <= 20'b00000000000000000000;
        10'b1110000000: data <= 20'b00100000000010000000;
        10'b1110000001: data <= 20'b00000000000010000000;
        10'b1110000010: data <= 20'b00100000000000000000;
        10'b1110000011: data <= 20'b00000000000000000000;
        10'b1110000100: data <= 20'b00000000000010000000;
        10'b1110000101: data <= 20'b00000000000010000000;
        10'b1110000110: data <= 20'b00000000000010000000;
        10'b1110000111: data <= 20'b00100000000000000000;
        10'b1110001000: data <= 20'b00000000000010000000;
        10'b1110001001: data <= 20'b00000000000010000000;
        10'b1110001010: data <= 20'b00000000000010000000;
        10'b1110001011: data <= 20'b00000000000010000000;
        10'b1110001100: data <= 20'b00100000000010000000;
        10'b1110001101: data <= 20'b00100000000010000000;
        10'b1110001110: data <= 20'b00000000000010000000;
        10'b1110001111: data <= 20'b00100000000000000000;
        10'b1110010000: data <= 20'b00000000000000000000;
        10'b1110010001: data <= 20'b00000000000010000000;
        10'b1110010010: data <= 20'b00000000000000000000;
        10'b1110010011: data <= 20'b00000000000000000000;
        10'b1110010100: data <= 20'b00000000000010000000;
        10'b1110010101: data <= 20'b00000000000010000000;
        10'b1110010110: data <= 20'b00000000000010000000;
        10'b1110010111: data <= 20'b00100000000000000000;
        10'b1110011000: data <= 20'b00000000000010000000;
        10'b1110011001: data <= 20'b00100000000000000000;
        10'b1110011010: data <= 20'b00000000000010000000;
        10'b1110011011: data <= 20'b00000000000010000000;
        10'b1110011100: data <= 20'b00000000000000000000;
        10'b1110011101: data <= 20'b00000000000010000000;
        10'b1110011110: data <= 20'b00100000000000000000;
        10'b1110011111: data <= 20'b00100000000000000000;
        10'b1110100000: data <= 20'b00000000000010000000;
        10'b1110100001: data <= 20'b00000000000000000000;
        10'b1110100010: data <= 20'b00100000000000000000;
        10'b1110100011: data <= 20'b00000000000010000000;
        10'b1110100100: data <= 20'b00000000000000000000;
        10'b1110100101: data <= 20'b00100000000010000000;
        10'b1110100110: data <= 20'b00100000000000000000;
        10'b1110100111: data <= 20'b00100000000010000000;
        10'b1110101000: data <= 20'b00100000000010000000;
        10'b1110101001: data <= 20'b00000000000010000000;
        10'b1110101010: data <= 20'b00100000000010000000;
        10'b1110101011: data <= 20'b00000000000000000000;
        10'b1110101100: data <= 20'b00000000000000000000;
        10'b1110101101: data <= 20'b00100000000000000000;
        10'b1110101110: data <= 20'b00100000000000000000;
        10'b1110101111: data <= 20'b00100000000000000000;
        10'b1110110000: data <= 20'b00000000000000000000;
        10'b1110110001: data <= 20'b00000000000010000000;
        10'b1110110010: data <= 20'b00000000000000000000;
        10'b1110110011: data <= 20'b00100000000000000000;
        10'b1110110100: data <= 20'b00100000000000000000;
        10'b1110110101: data <= 20'b00000000000000000000;
        10'b1110110110: data <= 20'b00000000000010000000;
        10'b1110110111: data <= 20'b00100000000010000000;
        10'b1110111000: data <= 20'b00100000000000000000;
        10'b1110111001: data <= 20'b00100000000000000000;
        10'b1110111010: data <= 20'b00100000000010000000;
        10'b1110111011: data <= 20'b00000000000000000000;
        10'b1110111100: data <= 20'b00100000000010000000;
        10'b1110111101: data <= 20'b00100000000010000000;
        10'b1110111110: data <= 20'b00100000000010000000;
        10'b1110111111: data <= 20'b00000000000000000000;
        10'b1111000000: data <= 20'b00100000000010000000;
        10'b1111000001: data <= 20'b00000000000000000000;
        10'b1111000010: data <= 20'b00000000000010000000;
        10'b1111000011: data <= 20'b00100000000010000000;
        10'b1111000100: data <= 20'b00100000000000000000;
        10'b1111000101: data <= 20'b00000000000010000000;
        10'b1111000110: data <= 20'b00100000000010000000;
        10'b1111000111: data <= 20'b00100000000010000000;
        10'b1111001000: data <= 20'b00100000000010000000;
        10'b1111001001: data <= 20'b00000000000010000000;
        10'b1111001010: data <= 20'b00100000000000000000;
        10'b1111001011: data <= 20'b00000000000010000000;
        10'b1111001100: data <= 20'b00000000000010000000;
        10'b1111001101: data <= 20'b00000000000010000000;
        10'b1111001110: data <= 20'b00100000000010000000;
        10'b1111001111: data <= 20'b00000000000000000000;
        10'b1111010000: data <= 20'b00000000000010000000;
        10'b1111010001: data <= 20'b00000000000010000000;
        10'b1111010010: data <= 20'b00100000000000000000;
        10'b1111010011: data <= 20'b00100000000000000000;
        10'b1111010100: data <= 20'b00100000000010000000;
        10'b1111010101: data <= 20'b00000000000000000000;
        10'b1111010110: data <= 20'b00100000000000000000;
        10'b1111010111: data <= 20'b00100000000010000000;
        10'b1111011000: data <= 20'b00100000100000000000;
        10'b1111011001: data <= 20'b00000000000010000000;
        10'b1111011010: data <= 20'b00000000000010000000;
        10'b1111011011: data <= 20'b00000000000000000000;
        10'b1111011100: data <= 20'b00000000000010000000;
        10'b1111011101: data <= 20'b00000000000010000000;
        10'b1111011110: data <= 20'b00100000000000000000;
        10'b1111011111: data <= 20'b00000000000000000000;
        10'b1111100000: data <= 20'b00100000000010000000;
        10'b1111100001: data <= 20'b00000000000000000000;
        10'b1111100010: data <= 20'b00100000000000000000;
        10'b1111100011: data <= 20'b00000000000000000000;
        10'b1111100100: data <= 20'b00100000000000000000;
        10'b1111100101: data <= 20'b00000000000010000000;
        10'b1111100110: data <= 20'b00100000000000000000;
        10'b1111100111: data <= 20'b00000000000000000000;
        10'b1111101000: data <= 20'b00100000010010000000;
        10'b1111101001: data <= 20'b00000000000010000000;
        10'b1111101010: data <= 20'b00000000000000000000;
        10'b1111101011: data <= 20'b00000000000000000000;
        10'b1111101100: data <= 20'b00100000000000000000;
        10'b1111101101: data <= 20'b00100000000010000000;
        10'b1111101110: data <= 20'b00000000000010000000;
        10'b1111101111: data <= 20'b00000000000010000000;
        10'b1111110000: data <= 20'b00000000000000000000;
        10'b1111110001: data <= 20'b00100000000010000000;
        10'b1111110010: data <= 20'b00100000000010000000;
        10'b1111110011: data <= 20'b00000000000010000000;
        10'b1111110100: data <= 20'b00000000000010000000;
        10'b1111110101: data <= 20'b00100000000010000000;
        10'b1111110110: data <= 20'b00000000000000000000;
        10'b1111110111: data <= 20'b00000000000000000000;
        10'b1111111000: data <= 20'b00100000000010000000;
        10'b1111111001: data <= 20'b00100000000000000000;
        10'b1111111010: data <= 20'b00100000000010000000;
        10'b1111111011: data <= 20'b00100000000000000000;
        10'b1111111100: data <= 20'b00100000000010000000;
    
    endcase
    end
    end

    assign Q = data;

    endmodule

        