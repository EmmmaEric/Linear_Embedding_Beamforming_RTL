
module memory_rom_22(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3e57a8bf;
    11'b00000000001: data <= 32'h3adeac12;
    11'b00000000010: data <= 32'hbbc3a7a1;
    11'b00000000011: data <= 32'hbeb0bac9;
    11'b00000000100: data <= 32'hb01abee9;
    11'b00000000101: data <= 32'h3f12be46;
    11'b00000000110: data <= 32'h3e7aba83;
    11'b00000000111: data <= 32'hb1b1b841;
    11'b00000001000: data <= 32'hbd18b76d;
    11'b00000001001: data <= 32'hbade35f3;
    11'b00000001010: data <= 32'hb7363df6;
    11'b00000001011: data <= 32'hbc813ccc;
    11'b00000001100: data <= 32'hbf52b8f6;
    11'b00000001101: data <= 32'hbd0dbef2;
    11'b00000001110: data <= 32'h2778b86f;
    11'b00000001111: data <= 32'h39a43e00;
    11'b00000010000: data <= 32'h39e63fe5;
    11'b00000010001: data <= 32'h3bcb3ab5;
    11'b00000010010: data <= 32'h3cd33266;
    11'b00000010011: data <= 32'h36f13b2f;
    11'b00000010100: data <= 32'hbb993d6b;
    11'b00000010101: data <= 32'hbc513404;
    11'b00000010110: data <= 32'h3903bd8d;
    11'b00000010111: data <= 32'h405fbf5b;
    11'b00000011000: data <= 32'h3ec2bc9a;
    11'b00000011001: data <= 32'h29b1b893;
    11'b00000011010: data <= 32'hb764b5da;
    11'b00000011011: data <= 32'h35dd3105;
    11'b00000011100: data <= 32'h37f53a0f;
    11'b00000011101: data <= 32'hbc06342d;
    11'b00000011110: data <= 32'hc0e4bcf8;
    11'b00000011111: data <= 32'hc00cbf8b;
    11'b00000100000: data <= 32'hb677b8fc;
    11'b00000100001: data <= 32'h38573c0f;
    11'b00000100010: data <= 32'h36b73c56;
    11'b00000100011: data <= 32'h33a130b3;
    11'b00000100100: data <= 32'h346f351c;
    11'b00000100101: data <= 32'hb20d3f51;
    11'b00000100110: data <= 32'hbc1a40fb;
    11'b00000100111: data <= 32'hbb2b3beb;
    11'b00000101000: data <= 32'h3879bc68;
    11'b00000101001: data <= 32'h3eeabe57;
    11'b00000101010: data <= 32'h3d35b8a4;
    11'b00000101011: data <= 32'h359731af;
    11'b00000101100: data <= 32'h39382ddc;
    11'b00000101101: data <= 32'h3eed2844;
    11'b00000101110: data <= 32'h3da13458;
    11'b00000101111: data <= 32'hb9f9ad35;
    11'b00000110000: data <= 32'hc0ddbcc9;
    11'b00000110001: data <= 32'hbf2bbf12;
    11'b00000110010: data <= 32'h28d7bc0d;
    11'b00000110011: data <= 32'h3a08ae34;
    11'b00000110100: data <= 32'h2b8bb4bd;
    11'b00000110101: data <= 32'hb844ba1e;
    11'b00000110110: data <= 32'hb64b328f;
    11'b00000110111: data <= 32'hb6e94057;
    11'b00000111000: data <= 32'hbc32416e;
    11'b00000111001: data <= 32'hbcf03b72;
    11'b00000111010: data <= 32'hb5f4bc4c;
    11'b00000111011: data <= 32'h3854bc3d;
    11'b00000111100: data <= 32'h387435f1;
    11'b00000111101: data <= 32'h375d3c2d;
    11'b00000111110: data <= 32'h3d77375e;
    11'b00000111111: data <= 32'h40d826aa;
    11'b00001000000: data <= 32'h3eec3672;
    11'b00001000001: data <= 32'hb85e3841;
    11'b00001000010: data <= 32'hbf92b55c;
    11'b00001000011: data <= 32'hbacbbd2d;
    11'b00001000100: data <= 32'h3b6dbd80;
    11'b00001000101: data <= 32'h3c64bc79;
    11'b00001000110: data <= 32'hb00dbd63;
    11'b00001000111: data <= 32'hb9edbd7d;
    11'b00001001000: data <= 32'hb1f6abce;
    11'b00001001001: data <= 32'h2c303f23;
    11'b00001001010: data <= 32'hbac83ff9;
    11'b00001001011: data <= 32'hbf313294;
    11'b00001001100: data <= 32'hbe50bd1b;
    11'b00001001101: data <= 32'hb98cb90f;
    11'b00001001110: data <= 32'hb1273bb7;
    11'b00001001111: data <= 32'h344f3d0e;
    11'b00001010000: data <= 32'h3d13349a;
    11'b00001010001: data <= 32'h402b9ed3;
    11'b00001010010: data <= 32'h3d4a3c1c;
    11'b00001010011: data <= 32'hb8483f0c;
    11'b00001010100: data <= 32'hbd003b31;
    11'b00001010101: data <= 32'h2b85b938;
    11'b00001010110: data <= 32'h3e03bd9d;
    11'b00001010111: data <= 32'h3ca2bd97;
    11'b00001011000: data <= 32'hb072bdd3;
    11'b00001011001: data <= 32'hb3eabd5b;
    11'b00001011010: data <= 32'h3b08b4aa;
    11'b00001011011: data <= 32'h3c933c0f;
    11'b00001011100: data <= 32'hb67e3b7a;
    11'b00001011101: data <= 32'hc045b87a;
    11'b00001011110: data <= 32'hc088bdc0;
    11'b00001011111: data <= 32'hbce5b806;
    11'b00001100000: data <= 32'hb7143a34;
    11'b00001100001: data <= 32'hae62384b;
    11'b00001100010: data <= 32'h3807b830;
    11'b00001100011: data <= 32'h3c45b2e2;
    11'b00001100100: data <= 32'h389b3ea2;
    11'b00001100101: data <= 32'hb91d41a0;
    11'b00001100110: data <= 32'hbb3d3f0a;
    11'b00001100111: data <= 32'h343ab235;
    11'b00001101000: data <= 32'h3cdabc37;
    11'b00001101001: data <= 32'h395cba62;
    11'b00001101010: data <= 32'hb0fbb93d;
    11'b00001101011: data <= 32'h386eba4c;
    11'b00001101100: data <= 32'h404cb610;
    11'b00001101101: data <= 32'h4064366b;
    11'b00001101110: data <= 32'h2ce0357e;
    11'b00001101111: data <= 32'hbfecb980;
    11'b00001110000: data <= 32'hc000bcf9;
    11'b00001110001: data <= 32'hba20b8b2;
    11'b00001110010: data <= 32'hb19ea4d9;
    11'b00001110011: data <= 32'hb6e2b9ee;
    11'b00001110100: data <= 32'hb5e3be5f;
    11'b00001110101: data <= 32'h3195b8be;
    11'b00001110110: data <= 32'h30ee3f47;
    11'b00001110111: data <= 32'hb8f141ff;
    11'b00001111000: data <= 32'hbbb33ee2;
    11'b00001111001: data <= 32'hb59db18e;
    11'b00001111010: data <= 32'h3064b853;
    11'b00001111011: data <= 32'hb3b3337a;
    11'b00001111100: data <= 32'hb574367a;
    11'b00001111101: data <= 32'h3c37b3b4;
    11'b00001111110: data <= 32'h4199b670;
    11'b00001111111: data <= 32'h41283489;
    11'b00010000000: data <= 32'h3529392b;
    11'b00010000001: data <= 32'hbdb42a25;
    11'b00010000010: data <= 32'hbbecb8e2;
    11'b00010000011: data <= 32'h3497b90f;
    11'b00010000100: data <= 32'h355dba62;
    11'b00010000101: data <= 32'hb8dfbf00;
    11'b00010000110: data <= 32'hba55c099;
    11'b00010000111: data <= 32'h2d36bbae;
    11'b00010001000: data <= 32'h38123d8a;
    11'b00010001001: data <= 32'hb45d4070;
    11'b00010001010: data <= 32'hbcce3aef;
    11'b00010001011: data <= 32'hbd2cb830;
    11'b00010001100: data <= 32'hbc35b043;
    11'b00010001101: data <= 32'hbc5e3c0d;
    11'b00010001110: data <= 32'hb9823b4b;
    11'b00010001111: data <= 32'h3afcb411;
    11'b00010010000: data <= 32'h40d3b86c;
    11'b00010010001: data <= 32'h402938b8;
    11'b00010010010: data <= 32'h32e33e62;
    11'b00010010011: data <= 32'hba733ceb;
    11'b00010010100: data <= 32'h2d193232;
    11'b00010010101: data <= 32'h3c8ab73d;
    11'b00010010110: data <= 32'h388ebbab;
    11'b00010010111: data <= 32'hb9adbf4a;
    11'b00010011000: data <= 32'hb8cfc070;
    11'b00010011001: data <= 32'h3adcbc73;
    11'b00010011010: data <= 32'h3e18390f;
    11'b00010011011: data <= 32'h358b3c12;
    11'b00010011100: data <= 32'hbd27b0fc;
    11'b00010011101: data <= 32'hbf51baf3;
    11'b00010011110: data <= 32'hbe3a2b25;
    11'b00010011111: data <= 32'hbd833c6f;
    11'b00010100000: data <= 32'hbc1f37ac;
    11'b00010100001: data <= 32'h2f15bbe4;
    11'b00010100010: data <= 32'h3d19bb87;
    11'b00010100011: data <= 32'h3c643b87;
    11'b00010100100: data <= 32'hacf340ef;
    11'b00010100101: data <= 32'hb6d34024;
    11'b00010100110: data <= 32'h386539a8;
    11'b00010100111: data <= 32'h3c94acb4;
    11'b00010101000: data <= 32'h31c0b572;
    11'b00010101001: data <= 32'hbb2fbb5c;
    11'b00010101010: data <= 32'hae25bdda;
    11'b00010101011: data <= 32'h3fb3bc12;
    11'b00010101100: data <= 32'h41201cbc;
    11'b00010101101: data <= 32'h3b6d31d0;
    11'b00010101110: data <= 32'hbc30b8b5;
    11'b00010101111: data <= 32'hbe12ba60;
    11'b00010110000: data <= 32'hbc123012;
    11'b00010110001: data <= 32'hbb9438f1;
    11'b00010110010: data <= 32'hbccbb89e;
    11'b00010110011: data <= 32'hba19c016;
    11'b00010110100: data <= 32'h310abdd2;
    11'b00010110101: data <= 32'h35e53bb4;
    11'b00010110110: data <= 32'hb28e4128;
    11'b00010110111: data <= 32'hb5a23fe5;
    11'b00010111000: data <= 32'h33b038e3;
    11'b00010111001: data <= 32'h34ee34fc;
    11'b00010111010: data <= 32'hb9b73984;
    11'b00010111011: data <= 32'hbcfd357e;
    11'b00010111100: data <= 32'h3315b8e9;
    11'b00010111101: data <= 32'h40f5baf3;
    11'b00010111110: data <= 32'h41cfb2fa;
    11'b00010111111: data <= 32'h3c7131d1;
    11'b00011000000: data <= 32'hb89faf28;
    11'b00011000001: data <= 32'hb805b231;
    11'b00011000010: data <= 32'h32f63434;
    11'b00011000011: data <= 32'hb0b92b70;
    11'b00011000100: data <= 32'hbcc3bde1;
    11'b00011000101: data <= 32'hbd0ec177;
    11'b00011000110: data <= 32'hb35fbf3f;
    11'b00011000111: data <= 32'h371a3886;
    11'b00011001000: data <= 32'h2d9b3f22;
    11'b00011001001: data <= 32'hb6803baa;
    11'b00011001010: data <= 32'hb7419c89;
    11'b00011001011: data <= 32'hb9f7383e;
    11'b00011001100: data <= 32'hbe463e1b;
    11'b00011001101: data <= 32'hbe8d3c8a;
    11'b00011001110: data <= 32'h26ffb546;
    11'b00011001111: data <= 32'h4021bb7f;
    11'b00011010000: data <= 32'h408bada1;
    11'b00011010001: data <= 32'h3a293ae6;
    11'b00011010010: data <= 32'hb05c3b4c;
    11'b00011010011: data <= 32'h38e53900;
    11'b00011010100: data <= 32'h3d5c3847;
    11'b00011010101: data <= 32'h365fa92c;
    11'b00011010110: data <= 32'hbcb7be03;
    11'b00011010111: data <= 32'hbcefc119;
    11'b00011011000: data <= 32'h3435bf19;
    11'b00011011001: data <= 32'h3d1ba762;
    11'b00011011010: data <= 32'h39c8385d;
    11'b00011011011: data <= 32'hb5cab53f;
    11'b00011011100: data <= 32'hbb0db95c;
    11'b00011011101: data <= 32'hbccb38a5;
    11'b00011011110: data <= 32'hbf243f0d;
    11'b00011011111: data <= 32'hbf5d3bf4;
    11'b00011100000: data <= 32'hb8dabad4;
    11'b00011100001: data <= 32'h3b24bd53;
    11'b00011100010: data <= 32'h3c292ed3;
    11'b00011100011: data <= 32'h30f83e55;
    11'b00011100100: data <= 32'h2d5a3ec1;
    11'b00011100101: data <= 32'h3cd23c69;
    11'b00011100110: data <= 32'h3e983aaa;
    11'b00011100111: data <= 32'h33cd37cc;
    11'b00011101000: data <= 32'hbd6cb88d;
    11'b00011101001: data <= 32'hbb2ebe43;
    11'b00011101010: data <= 32'h3c98bd78;
    11'b00011101011: data <= 32'h4078b7be;
    11'b00011101100: data <= 32'h3d31b662;
    11'b00011101101: data <= 32'hb09dbc44;
    11'b00011101110: data <= 32'hb8f0bae7;
    11'b00011101111: data <= 32'hb90738ec;
    11'b00011110000: data <= 32'hbca33dc8;
    11'b00011110001: data <= 32'hbee230b0;
    11'b00011110010: data <= 32'hbd37bf41;
    11'b00011110011: data <= 32'hb51ebf71;
    11'b00011110100: data <= 32'h03f52e6b;
    11'b00011110101: data <= 32'hb43f3ecd;
    11'b00011110110: data <= 32'h2df43e3c;
    11'b00011110111: data <= 32'h3c453acb;
    11'b00011111000: data <= 32'h3c2f3bbd;
    11'b00011111001: data <= 32'hb8423d67;
    11'b00011111010: data <= 32'hbeec3a3a;
    11'b00011111011: data <= 32'hb936b680;
    11'b00011111100: data <= 32'h3eabbb33;
    11'b00011111101: data <= 32'h4117b8e3;
    11'b00011111110: data <= 32'h3d72b885;
    11'b00011111111: data <= 32'h2fd1baca;
    11'b00100000000: data <= 32'h3409b679;
    11'b00100000001: data <= 32'h39743a3c;
    11'b00100000010: data <= 32'hab773bed;
    11'b00100000011: data <= 32'hbd86b968;
    11'b00100000100: data <= 32'hbebcc0f0;
    11'b00100000101: data <= 32'hbaedc047;
    11'b00100000110: data <= 32'hb2a3b0ac;
    11'b00100000111: data <= 32'hb0e83c18;
    11'b00100001000: data <= 32'h2b75379d;
    11'b00100001001: data <= 32'h380baa55;
    11'b00100001010: data <= 32'h2e1b3ad7;
    11'b00100001011: data <= 32'hbd674018;
    11'b00100001100: data <= 32'hc02a3ee0;
    11'b00100001101: data <= 32'hb9f931d7;
    11'b00100001110: data <= 32'h3d5eb9ff;
    11'b00100001111: data <= 32'h3f68b7b1;
    11'b00100010000: data <= 32'h3a1ca85e;
    11'b00100010001: data <= 32'h33df28dd;
    11'b00100010010: data <= 32'h3ce035ec;
    11'b00100010011: data <= 32'h3fc83c2f;
    11'b00100010100: data <= 32'h3a793ac3;
    11'b00100010101: data <= 32'hbc74ba28;
    11'b00100010110: data <= 32'hbe81c07a;
    11'b00100010111: data <= 32'hb842bf83;
    11'b00100011000: data <= 32'h3743b728;
    11'b00100011001: data <= 32'h36b7ac5c;
    11'b00100011010: data <= 32'h2fb3bb91;
    11'b00100011011: data <= 32'h2d02bc31;
    11'b00100011100: data <= 32'hb63938ef;
    11'b00100011101: data <= 32'hbe244076;
    11'b00100011110: data <= 32'hc0363ef9;
    11'b00100011111: data <= 32'hbc7db059;
    11'b00100100000: data <= 32'h34f1bc37;
    11'b00100100001: data <= 32'h37e0b507;
    11'b00100100010: data <= 32'hb2023929;
    11'b00100100011: data <= 32'h30f13a88;
    11'b00100100100: data <= 32'h3ef23aa0;
    11'b00100100101: data <= 32'h40d93cd8;
    11'b00100100110: data <= 32'h3b273ca1;
    11'b00100100111: data <= 32'hbcaa28bc;
    11'b00100101000: data <= 32'hbd44bc8d;
    11'b00100101001: data <= 32'h3476bc8f;
    11'b00100101010: data <= 32'h3d87b89e;
    11'b00100101011: data <= 32'h3bdcbb5d;
    11'b00100101100: data <= 32'h3406bf72;
    11'b00100101101: data <= 32'h319ebe0e;
    11'b00100101110: data <= 32'h2c5b37d7;
    11'b00100101111: data <= 32'hba7a3fb7;
    11'b00100110000: data <= 32'hbeb13bf5;
    11'b00100110001: data <= 32'hbdf9bc23;
    11'b00100110010: data <= 32'hba64be47;
    11'b00100110011: data <= 32'hb9d6b45e;
    11'b00100110100: data <= 32'hbb533b0d;
    11'b00100110101: data <= 32'ha8e73a3f;
    11'b00100110110: data <= 32'h3e6737f2;
    11'b00100110111: data <= 32'h3fc53c44;
    11'b00100111000: data <= 32'h32d53ed4;
    11'b00100111001: data <= 32'hbe133d16;
    11'b00100111010: data <= 32'hbc353283;
    11'b00100111011: data <= 32'h3afbb568;
    11'b00100111100: data <= 32'h3f13b76a;
    11'b00100111101: data <= 32'h3bedbc49;
    11'b00100111110: data <= 32'h347bbf25;
    11'b00100111111: data <= 32'h3a0bbcc3;
    11'b00101000000: data <= 32'h3d0e38e7;
    11'b00101000001: data <= 32'h377e3de8;
    11'b00101000010: data <= 32'hbbda3050;
    11'b00101000011: data <= 32'hbe64befd;
    11'b00101000100: data <= 32'hbd41bf41;
    11'b00101000101: data <= 32'hbc68b538;
    11'b00101000110: data <= 32'hbbdc3760;
    11'b00101000111: data <= 32'hb08db218;
    11'b00101001000: data <= 32'h3c35b889;
    11'b00101001001: data <= 32'h3beb38cb;
    11'b00101001010: data <= 32'hb9254036;
    11'b00101001011: data <= 32'hbf6b4054;
    11'b00101001100: data <= 32'hbbfd3bce;
    11'b00101001101: data <= 32'h3a272906;
    11'b00101001110: data <= 32'h3cbbb33f;
    11'b00101001111: data <= 32'h33d7b876;
    11'b00101010000: data <= 32'h2b9ebb72;
    11'b00101010001: data <= 32'h3da9b673;
    11'b00101010010: data <= 32'h40f03b03;
    11'b00101010011: data <= 32'h3e233ce5;
    11'b00101010100: data <= 32'hb715b0a5;
    11'b00101010101: data <= 32'hbd91be7c;
    11'b00101010110: data <= 32'hbbf0bdb6;
    11'b00101010111: data <= 32'hb80cb4e0;
    11'b00101011000: data <= 32'hb6e3b537;
    11'b00101011001: data <= 32'had26be30;
    11'b00101011010: data <= 32'h386fbf1a;
    11'b00101011011: data <= 32'h35ab2ac2;
    11'b00101011100: data <= 32'hbb704033;
    11'b00101011101: data <= 32'hbf204063;
    11'b00101011110: data <= 32'hbc543a0c;
    11'b00101011111: data <= 32'h27edb277;
    11'b00101100000: data <= 32'haedfaa47;
    11'b00101100001: data <= 32'hbb5f313d;
    11'b00101100010: data <= 32'hb5e4a8c2;
    11'b00101100011: data <= 32'h3ed830ea;
    11'b00101100100: data <= 32'h41e43bd3;
    11'b00101100101: data <= 32'h3f003d21;
    11'b00101100110: data <= 32'hb624361f;
    11'b00101100111: data <= 32'hbc31b8c6;
    11'b00101101000: data <= 32'hb112b7a5;
    11'b00101101001: data <= 32'h3803ad34;
    11'b00101101010: data <= 32'h3307bb71;
    11'b00101101011: data <= 32'h2403c0e9;
    11'b00101101100: data <= 32'h370bc0cf;
    11'b00101101101: data <= 32'h386bb38a;
    11'b00101101110: data <= 32'hb4a03ef1;
    11'b00101101111: data <= 32'hbc9b3dbd;
    11'b00101110000: data <= 32'hbc61b1f8;
    11'b00101110001: data <= 32'hba7dba49;
    11'b00101110010: data <= 32'hbd471f25;
    11'b00101110011: data <= 32'hbf5f388d;
    11'b00101110100: data <= 32'hba2e312f;
    11'b00101110101: data <= 32'h3de9ad4f;
    11'b00101110110: data <= 32'h40eb3949;
    11'b00101110111: data <= 32'h3c3f3def;
    11'b00101111000: data <= 32'hba3a3d5d;
    11'b00101111001: data <= 32'hba3b39d9;
    11'b00101111010: data <= 32'h388d385b;
    11'b00101111011: data <= 32'h3c6334ae;
    11'b00101111100: data <= 32'h3551bb9b;
    11'b00101111101: data <= 32'hae29c0c4;
    11'b00101111110: data <= 32'h398dc039;
    11'b00101111111: data <= 32'h3de1aed3;
    11'b00110000000: data <= 32'h3bbc3d1a;
    11'b00110000001: data <= 32'hb3273783;
    11'b00110000010: data <= 32'hbb30bc54;
    11'b00110000011: data <= 32'hbca5bc90;
    11'b00110000100: data <= 32'hbecf2bce;
    11'b00110000101: data <= 32'hbff23721;
    11'b00110000110: data <= 32'hbb52b846;
    11'b00110000111: data <= 32'h3b4cbc75;
    11'b00110001000: data <= 32'h3db4aa06;
    11'b00110001001: data <= 32'h2a293e35;
    11'b00110001010: data <= 32'hbce74015;
    11'b00110001011: data <= 32'hb9303e16;
    11'b00110001100: data <= 32'h39d63c2e;
    11'b00110001101: data <= 32'h3a3a38f5;
    11'b00110001110: data <= 32'hb5e0b66d;
    11'b00110001111: data <= 32'hb863bde1;
    11'b00110010000: data <= 32'h3c09bccc;
    11'b00110010001: data <= 32'h40ec343a;
    11'b00110010010: data <= 32'h401c3bc7;
    11'b00110010011: data <= 32'h37b8a98e;
    11'b00110010100: data <= 32'hb85fbcdc;
    11'b00110010101: data <= 32'hba40ba8a;
    11'b00110010110: data <= 32'hbc4734bd;
    11'b00110010111: data <= 32'hbd641b4a;
    11'b00110011000: data <= 32'hba18bea6;
    11'b00110011001: data <= 32'h3622c0b1;
    11'b00110011010: data <= 32'h38b4ba5f;
    11'b00110011011: data <= 32'hb7d03d63;
    11'b00110011100: data <= 32'hbcf13fef;
    11'b00110011101: data <= 32'hb8593d22;
    11'b00110011110: data <= 32'h35433a1a;
    11'b00110011111: data <= 32'hb46539e1;
    11'b00110100000: data <= 32'hbe3a3571;
    11'b00110100001: data <= 32'hbcd3b670;
    11'b00110100010: data <= 32'h3c3fb678;
    11'b00110100011: data <= 32'h41a5377c;
    11'b00110100100: data <= 32'h408b3afd;
    11'b00110100101: data <= 32'h38693123;
    11'b00110100110: data <= 32'hb32eb6f9;
    11'b00110100111: data <= 32'h2cbc30c7;
    11'b00110101000: data <= 32'h2d623a21;
    11'b00110101001: data <= 32'hb7a4b529;
    11'b00110101010: data <= 32'hb863c0de;
    11'b00110101011: data <= 32'h30a7c1fd;
    11'b00110101100: data <= 32'h37b1bc96;
    11'b00110101101: data <= 32'hae7e3ba4;
    11'b00110101110: data <= 32'hb8d53cc5;
    11'b00110101111: data <= 32'hb4e13316;
    11'b00110110000: data <= 32'hb2b5a396;
    11'b00110110001: data <= 32'hbd55395a;
    11'b00110110010: data <= 32'hc1083ab7;
    11'b00110110011: data <= 32'hbee62d26;
    11'b00110110100: data <= 32'h3a02b611;
    11'b00110110101: data <= 32'h40953183;
    11'b00110110110: data <= 32'h3df53aa6;
    11'b00110110111: data <= 32'h99883a65;
    11'b00110111000: data <= 32'hac6539c8;
    11'b00110111001: data <= 32'h3afc3ce5;
    11'b00110111010: data <= 32'h3b853d35;
    11'b00110111011: data <= 32'hae51b2ec;
    11'b00110111100: data <= 32'hb8e3c09b;
    11'b00110111101: data <= 32'h319ac146;
    11'b00110111110: data <= 32'h3c49bb34;
    11'b00110111111: data <= 32'h3bc038ba;
    11'b00111000000: data <= 32'h3622316a;
    11'b00111000001: data <= 32'h2e08bb4e;
    11'b00111000010: data <= 32'hb62fb915;
    11'b00111000011: data <= 32'hbe94392e;
    11'b00111000100: data <= 32'hc1403b4f;
    11'b00111000101: data <= 32'hbf32b4a7;
    11'b00111000110: data <= 32'h3407bcd4;
    11'b00111000111: data <= 32'h3cd3b8ba;
    11'b00111001000: data <= 32'h34243959;
    11'b00111001001: data <= 32'hb9b03d24;
    11'b00111001010: data <= 32'ha8713db6;
    11'b00111001011: data <= 32'h3cd13ee5;
    11'b00111001100: data <= 32'h3b853e79;
    11'b00111001101: data <= 32'hb8a034dc;
    11'b00111001110: data <= 32'hbc6bbd5d;
    11'b00111001111: data <= 32'h33d7be20;
    11'b00111010000: data <= 32'h3f42b482;
    11'b00111010001: data <= 32'h3fd5365b;
    11'b00111010010: data <= 32'h3c7cb7da;
    11'b00111010011: data <= 32'h37ebbd6e;
    11'b00111010100: data <= 32'h2069b866;
    11'b00111010101: data <= 32'hbbb43b3a;
    11'b00111010110: data <= 32'hbf4d39c0;
    11'b00111010111: data <= 32'hbdafbc98;
    11'b00111011000: data <= 32'hb131c0a7;
    11'b00111011001: data <= 32'h33b7bd95;
    11'b00111011010: data <= 32'hb8a935bf;
    11'b00111011011: data <= 32'hbbcd3ca9;
    11'b00111011100: data <= 32'h2c2f3c8f;
    11'b00111011101: data <= 32'h3c2c3d46;
    11'b00111011110: data <= 32'h318f3e2f;
    11'b00111011111: data <= 32'hbe8f3b7f;
    11'b00111100000: data <= 32'hbf56b144;
    11'b00111100001: data <= 32'h30a9b70d;
    11'b00111100010: data <= 32'h4024322f;
    11'b00111100011: data <= 32'h403d354e;
    11'b00111100100: data <= 32'h3c6db81d;
    11'b00111100101: data <= 32'h396ebb05;
    11'b00111100110: data <= 32'h3a313456;
    11'b00111100111: data <= 32'h34933dce;
    11'b00111101000: data <= 32'hb96638a3;
    11'b00111101001: data <= 32'hbb6abf1c;
    11'b00111101010: data <= 32'hb56ec1d5;
    11'b00111101011: data <= 32'hacf9bed1;
    11'b00111101100: data <= 32'hb80e2a62;
    11'b00111101101: data <= 32'hb81a36f8;
    11'b00111101110: data <= 32'h360d9f8f;
    11'b00111101111: data <= 32'h39bf3487;
    11'b00111110000: data <= 32'hb9ae3ccd;
    11'b00111110001: data <= 32'hc1143d6a;
    11'b00111110010: data <= 32'hc0b33818;
    11'b00111110011: data <= 32'hb072ae05;
    11'b00111110100: data <= 32'h3e452e12;
    11'b00111110101: data <= 32'h3d0b3357;
    11'b00111110110: data <= 32'h3530aeb8;
    11'b00111110111: data <= 32'h38902cf9;
    11'b00111111000: data <= 32'h3dea3d21;
    11'b00111111001: data <= 32'h3d45400b;
    11'b00111111010: data <= 32'h281739ba;
    11'b00111111011: data <= 32'hba19be8e;
    11'b00111111100: data <= 32'hb587c0fb;
    11'b00111111101: data <= 32'h346bbd10;
    11'b00111111110: data <= 32'h3553ad06;
    11'b00111111111: data <= 32'h366fb7e3;
    11'b01000000000: data <= 32'h3abcbd37;
    11'b01000000001: data <= 32'h38fbb956;
    11'b01000000010: data <= 32'hbbda3b68;
    11'b01000000011: data <= 32'hc12f3dbd;
    11'b01000000100: data <= 32'hc08c3606;
    11'b01000000101: data <= 32'hb70bb955;
    11'b01000000110: data <= 32'h388ab89e;
    11'b01000000111: data <= 32'hafb1a3b5;
    11'b01000001000: data <= 32'hb9ac3411;
    11'b01000001001: data <= 32'h354e39b0;
    11'b01000001010: data <= 32'h3f293ef4;
    11'b01000001011: data <= 32'h3e324079;
    11'b01000001100: data <= 32'hb1643c56;
    11'b01000001101: data <= 32'hbc8eb9fa;
    11'b01000001110: data <= 32'hb5c8bcfd;
    11'b01000001111: data <= 32'h3adbb553;
    11'b01000010000: data <= 32'h3ce0211e;
    11'b01000010001: data <= 32'h3c6bbc73;
    11'b01000010010: data <= 32'h3cc4bfe5;
    11'b01000010011: data <= 32'h3b59bb0e;
    11'b01000010100: data <= 32'hb5a23c22;
    11'b01000010101: data <= 32'hbead3d45;
    11'b01000010110: data <= 32'hbe6ab4b4;
    11'b01000010111: data <= 32'hb896be9c;
    11'b01000011000: data <= 32'hb57fbd68;
    11'b01000011001: data <= 32'hbcbab51f;
    11'b01000011010: data <= 32'hbd2e31bb;
    11'b01000011011: data <= 32'h34023742;
    11'b01000011100: data <= 32'h3ec53cec;
    11'b01000011101: data <= 32'h3be43f9e;
    11'b01000011110: data <= 32'hbc453dcd;
    11'b01000011111: data <= 32'hbf5535df;
    11'b01000100000: data <= 32'hb7e22b96;
    11'b01000100001: data <= 32'h3c6d37ba;
    11'b01000100010: data <= 32'h3d8e3110;
    11'b01000100011: data <= 32'h3c0bbcb9;
    11'b01000100100: data <= 32'h3ca3bed7;
    11'b01000100101: data <= 32'h3dc6b40a;
    11'b01000100110: data <= 32'h3aa83e23;
    11'b01000100111: data <= 32'hb4fc3cf2;
    11'b01000101000: data <= 32'hba0ebaf7;
    11'b01000101001: data <= 32'hb80ec074;
    11'b01000101010: data <= 32'hb980be69;
    11'b01000101011: data <= 32'hbd58b76e;
    11'b01000101100: data <= 32'hbc3ab597;
    11'b01000101101: data <= 32'h37f6b910;
    11'b01000101110: data <= 32'h3dc2190c;
    11'b01000101111: data <= 32'h32213cd4;
    11'b01000110000: data <= 32'hbfb83e67;
    11'b01000110001: data <= 32'hc09f3c33;
    11'b01000110010: data <= 32'hb94f392a;
    11'b01000110011: data <= 32'h3a143928;
    11'b01000110100: data <= 32'h38a530d1;
    11'b01000110101: data <= 32'h2afebace;
    11'b01000110110: data <= 32'h39b5bb03;
    11'b01000110111: data <= 32'h3f7e3996;
    11'b01000111000: data <= 32'h3f6b402a;
    11'b01000111001: data <= 32'h39243d3a;
    11'b01000111010: data <= 32'hb4bcbac3;
    11'b01000111011: data <= 32'hb61fbf5f;
    11'b01000111100: data <= 32'hb68fbc0c;
    11'b01000111101: data <= 32'hb92db47f;
    11'b01000111110: data <= 32'hb358bc08;
    11'b01000111111: data <= 32'h3b96bfa4;
    11'b01001000000: data <= 32'h3d49bccb;
    11'b01001000001: data <= 32'hb0c938d6;
    11'b01001000010: data <= 32'hc0073e0e;
    11'b01001000011: data <= 32'hc0393bd9;
    11'b01001000100: data <= 32'hb9833408;
    11'b01001000101: data <= 32'h22ef2e06;
    11'b01001000110: data <= 32'hba36ad17;
    11'b01001000111: data <= 32'hbceab80a;
    11'b01001001000: data <= 32'h3001b2dc;
    11'b01001001001: data <= 32'h3ff03cb8;
    11'b01001001010: data <= 32'h40474069;
    11'b01001001011: data <= 32'h392a3dc5;
    11'b01001001100: data <= 32'hb816b1de;
    11'b01001001101: data <= 32'hb5eab8fe;
    11'b01001001110: data <= 32'h3031314a;
    11'b01001001111: data <= 32'h33503168;
    11'b01001010000: data <= 32'h37cfbd9b;
    11'b01001010001: data <= 32'h3cf4c13f;
    11'b01001010010: data <= 32'h3dbdbe8f;
    11'b01001010011: data <= 32'h34753810;
    11'b01001010100: data <= 32'hbc7b3d5f;
    11'b01001010101: data <= 32'hbcd735da;
    11'b01001010110: data <= 32'hb75db97d;
    11'b01001010111: data <= 32'hb93fb96d;
    11'b01001011000: data <= 32'hbf80b5a4;
    11'b01001011001: data <= 32'hc020b72b;
    11'b01001011010: data <= 32'hb27cb4da;
    11'b01001011011: data <= 32'h3f3439a3;
    11'b01001011100: data <= 32'h3e8e3eab;
    11'b01001011101: data <= 32'hb17c3dd6;
    11'b01001011110: data <= 32'hbcb83976;
    11'b01001011111: data <= 32'hb7c739b5;
    11'b01001100000: data <= 32'h37753cfe;
    11'b01001100001: data <= 32'h384038d6;
    11'b01001100010: data <= 32'h36ebbd69;
    11'b01001100011: data <= 32'h3c22c0d9;
    11'b01001100100: data <= 32'h3e8cbc81;
    11'b01001100101: data <= 32'h3cdd3ba1;
    11'b01001100110: data <= 32'h34333d02;
    11'b01001100111: data <= 32'had41b423;
    11'b01001101000: data <= 32'hac84bd70;
    11'b01001101001: data <= 32'hbad0bbc4;
    11'b01001101010: data <= 32'hc031b5c5;
    11'b01001101011: data <= 32'hbfe8b987;
    11'b01001101100: data <= 32'haa29bc9d;
    11'b01001101101: data <= 32'h3e23b853;
    11'b01001101110: data <= 32'h3a9d397c;
    11'b01001101111: data <= 32'hbc663d0b;
    11'b01001110000: data <= 32'hbecc3cc2;
    11'b01001110001: data <= 32'hb8753d7b;
    11'b01001110010: data <= 32'h35ca3e67;
    11'b01001110011: data <= 32'hab5939dd;
    11'b01001110100: data <= 32'hb83fbbf6;
    11'b01001110101: data <= 32'h34ffbe63;
    11'b01001110110: data <= 32'h3ed1b085;
    11'b01001110111: data <= 32'h40153e28;
    11'b01001111000: data <= 32'h3d283d05;
    11'b01001111001: data <= 32'h38dcb6eb;
    11'b01001111010: data <= 32'h33a6bcb1;
    11'b01001111011: data <= 32'hb835b628;
    11'b01001111100: data <= 32'hbdbc2ceb;
    11'b01001111101: data <= 32'hbc9abbec;
    11'b01001111110: data <= 32'h36d8c070;
    11'b01001111111: data <= 32'h3d7fbf41;
    11'b01010000000: data <= 32'h353ab1b5;
    11'b01010000001: data <= 32'hbd743b83;
    11'b01010000010: data <= 32'hbe123c2f;
    11'b01010000011: data <= 32'hb5b73c16;
    11'b01010000100: data <= 32'ha9303c5e;
    11'b01010000101: data <= 32'hbccc37ff;
    11'b01010000110: data <= 32'hbf8ab901;
    11'b01010000111: data <= 32'hb87dba81;
    11'b01010001000: data <= 32'h3e2537fb;
    11'b01010001001: data <= 32'h40723ec8;
    11'b01010001010: data <= 32'h3d683ccc;
    11'b01010001011: data <= 32'h37b1adcd;
    11'b01010001100: data <= 32'h3487b16a;
    11'b01010001101: data <= 32'h28193add;
    11'b01010001110: data <= 32'hb78c3a9b;
    11'b01010001111: data <= 32'hb4bdbc4a;
    11'b01010010000: data <= 32'h3a21c19c;
    11'b01010010001: data <= 32'h3d56c0a8;
    11'b01010010010: data <= 32'h3769b692;
    11'b01010010011: data <= 32'hb970398b;
    11'b01010010100: data <= 32'hb87c368d;
    11'b01010010101: data <= 32'h318b2745;
    11'b01010010110: data <= 32'hb60932c3;
    11'b01010010111: data <= 32'hc04e3172;
    11'b01010011000: data <= 32'hc19cb73f;
    11'b01010011001: data <= 32'hbc49b925;
    11'b01010011010: data <= 32'h3cec3370;
    11'b01010011011: data <= 32'h3ec13c79;
    11'b01010011100: data <= 32'h380e3b63;
    11'b01010011101: data <= 32'hb43236e9;
    11'b01010011110: data <= 32'h2f363c0b;
    11'b01010011111: data <= 32'h37324015;
    11'b01010100000: data <= 32'h2b243df3;
    11'b01010100001: data <= 32'hb0bbbad3;
    11'b01010100010: data <= 32'h385dc11d;
    11'b01010100011: data <= 32'h3d0fbf40;
    11'b01010100100: data <= 32'h3c3a2c6c;
    11'b01010100101: data <= 32'h38493921;
    11'b01010100110: data <= 32'h3968b465;
    11'b01010100111: data <= 32'h3a9ebab0;
    11'b01010101000: data <= 32'hb5b9b470;
    11'b01010101001: data <= 32'hc09e30dc;
    11'b01010101010: data <= 32'hc17db74d;
    11'b01010101011: data <= 32'hbb6dbca2;
    11'b01010101100: data <= 32'h3bd0bab0;
    11'b01010101101: data <= 32'h3aa126f3;
    11'b01010101110: data <= 32'hb8a536e9;
    11'b01010101111: data <= 32'hbbb93978;
    11'b01010110000: data <= 32'h20b33e5b;
    11'b01010110001: data <= 32'h386440e5;
    11'b01010110010: data <= 32'hb2e63eb7;
    11'b01010110011: data <= 32'hbb67b798;
    11'b01010110100: data <= 32'hb465bec0;
    11'b01010110101: data <= 32'h3c19b993;
    11'b01010110110: data <= 32'h3e613a92;
    11'b01010110111: data <= 32'h3de13989;
    11'b01010111000: data <= 32'h3dccb8f1;
    11'b01010111001: data <= 32'h3d06bb92;
    11'b01010111010: data <= 32'h27702f61;
    11'b01010111011: data <= 32'hbe6c395d;
    11'b01010111100: data <= 32'hbf45b72c;
    11'b01010111101: data <= 32'hb4f3bfac;
    11'b01010111110: data <= 32'h3afbc002;
    11'b01010111111: data <= 32'h3210bb91;
    11'b01011000000: data <= 32'hbc7bac1f;
    11'b01011000001: data <= 32'hbbe036f1;
    11'b01011000010: data <= 32'h34443cca;
    11'b01011000011: data <= 32'h37113f7f;
    11'b01011000100: data <= 32'hbc293d58;
    11'b01011000101: data <= 32'hc053b115;
    11'b01011000110: data <= 32'hbd18ba50;
    11'b01011000111: data <= 32'h39123258;
    11'b01011001000: data <= 32'h3e813cbd;
    11'b01011001001: data <= 32'h3df238d8;
    11'b01011001010: data <= 32'h3d30b868;
    11'b01011001011: data <= 32'h3cf1b42c;
    11'b01011001100: data <= 32'h385f3cec;
    11'b01011001101: data <= 32'hb8643e36;
    11'b01011001110: data <= 32'hb9d8b456;
    11'b01011001111: data <= 32'h33b0c09f;
    11'b01011010000: data <= 32'h3aa2c0ef;
    11'b01011010001: data <= 32'h2cd7bcc5;
    11'b01011010010: data <= 32'hba08b4cf;
    11'b01011010011: data <= 32'hb15ab1ff;
    11'b01011010100: data <= 32'h3b713004;
    11'b01011010101: data <= 32'h36393a4c;
    11'b01011010110: data <= 32'hbf153a63;
    11'b01011010111: data <= 32'hc20ea086;
    11'b01011011000: data <= 32'hbf5ab654;
    11'b01011011001: data <= 32'h347933e3;
    11'b01011011010: data <= 32'h3c493a1d;
    11'b01011011011: data <= 32'h3895329f;
    11'b01011011100: data <= 32'h361ab535;
    11'b01011011101: data <= 32'h3afb3961;
    11'b01011011110: data <= 32'h3b6540b5;
    11'b01011011111: data <= 32'h3196409c;
    11'b01011100000: data <= 32'hb45d2ae4;
    11'b01011100001: data <= 32'h3254c003;
    11'b01011100010: data <= 32'h3943bf90;
    11'b01011100011: data <= 32'h35e8b89f;
    11'b01011100100: data <= 32'h323cb1ff;
    11'b01011100101: data <= 32'h3c06ba9a;
    11'b01011100110: data <= 32'h3ed2bb48;
    11'b01011100111: data <= 32'h38869603;
    11'b01011101000: data <= 32'hbf5638a7;
    11'b01011101001: data <= 32'hc1d32bdb;
    11'b01011101010: data <= 32'hbe68b8f1;
    11'b01011101011: data <= 32'h30e1b84f;
    11'b01011101100: data <= 32'h3409b40e;
    11'b01011101101: data <= 32'hb954b6d6;
    11'b01011101110: data <= 32'hb8deb46d;
    11'b01011101111: data <= 32'h38723c80;
    11'b01011110000: data <= 32'h3c44416f;
    11'b01011110001: data <= 32'h31d440e6;
    11'b01011110010: data <= 32'hba0835a3;
    11'b01011110011: data <= 32'hb842bca6;
    11'b01011110100: data <= 32'h3441b91d;
    11'b01011110101: data <= 32'h39563717;
    11'b01011110110: data <= 32'h3bcb2d55;
    11'b01011110111: data <= 32'h3efdbcbd;
    11'b01011111000: data <= 32'h4046bd20;
    11'b01011111001: data <= 32'h3b682d6f;
    11'b01011111010: data <= 32'hbc8c3be4;
    11'b01011111011: data <= 32'hbf7832ef;
    11'b01011111100: data <= 32'hb9e7bc72;
    11'b01011111101: data <= 32'h343dbe18;
    11'b01011111110: data <= 32'hb626bcce;
    11'b01011111111: data <= 32'hbdccbbce;
    11'b01100000000: data <= 32'hbb88b873;
    11'b01100000001: data <= 32'h396339ba;
    11'b01100000010: data <= 32'h3c5d4017;
    11'b01100000011: data <= 32'hb5d53f95;
    11'b01100000100: data <= 32'hbf233772;
    11'b01100000101: data <= 32'hbe07b474;
    11'b01100000110: data <= 32'hb2fe37c3;
    11'b01100000111: data <= 32'h38e53c81;
    11'b01100001000: data <= 32'h3b933138;
    11'b01100001001: data <= 32'h3e11bcea;
    11'b01100001010: data <= 32'h3fccbb08;
    11'b01100001011: data <= 32'h3d113bc6;
    11'b01100001100: data <= 32'hae573f5b;
    11'b01100001101: data <= 32'hb8873825;
    11'b01100001110: data <= 32'h3051bd7a;
    11'b01100001111: data <= 32'h3698bfab;
    11'b01100010000: data <= 32'hb8afbd92;
    11'b01100010001: data <= 32'hbd78bc63;
    11'b01100010010: data <= 32'hb5fabc29;
    11'b01100010011: data <= 32'h3d2cb56f;
    11'b01100010100: data <= 32'h3cb93a18;
    11'b01100010101: data <= 32'hbb5a3c28;
    11'b01100010110: data <= 32'hc11c367c;
    11'b01100010111: data <= 32'hc01231be;
    11'b01100011000: data <= 32'hb81b3a87;
    11'b01100011001: data <= 32'h30b53bd4;
    11'b01100011010: data <= 32'h2944b182;
    11'b01100011011: data <= 32'h36d0bc9c;
    11'b01100011100: data <= 32'h3d22b0df;
    11'b01100011101: data <= 32'h3db33feb;
    11'b01100011110: data <= 32'h39574125;
    11'b01100011111: data <= 32'h31833ab1;
    11'b01100100000: data <= 32'h3639bc69;
    11'b01100100001: data <= 32'h354fbd56;
    11'b01100100010: data <= 32'hb70ab903;
    11'b01100100011: data <= 32'hb931b9b0;
    11'b01100100100: data <= 32'h394dbdd9;
    11'b01100100101: data <= 32'h4020bd9c;
    11'b01100100110: data <= 32'h3d98b4d5;
    11'b01100100111: data <= 32'hbbc53806;
    11'b01100101000: data <= 32'hc0d635a1;
    11'b01100101001: data <= 32'hbeb42e0e;
    11'b01100101010: data <= 32'hb6843482;
    11'b01100101011: data <= 32'hb7972fd5;
    11'b01100101100: data <= 32'hbcddba76;
    11'b01100101101: data <= 32'hbaa4bcbe;
    11'b01100101110: data <= 32'h390e33d1;
    11'b01100101111: data <= 32'h3da5409f;
    11'b01100110000: data <= 32'h3a5e413f;
    11'b01100110001: data <= 32'ha94e3b97;
    11'b01100110010: data <= 32'hb0c8b6db;
    11'b01100110011: data <= 32'hab1bac5a;
    11'b01100110100: data <= 32'hb413392f;
    11'b01100110101: data <= 32'h281fae61;
    11'b01100110110: data <= 32'h3d71be90;
    11'b01100110111: data <= 32'h40debf81;
    11'b01100111000: data <= 32'h3e80b7ee;
    11'b01100111001: data <= 32'hb68c3977;
    11'b01100111010: data <= 32'hbd6f37c1;
    11'b01100111011: data <= 32'hb899b445;
    11'b01100111100: data <= 32'h293fb88b;
    11'b01100111101: data <= 32'hbb50ba25;
    11'b01100111110: data <= 32'hc02cbd4f;
    11'b01100111111: data <= 32'hbdcfbd8d;
    11'b01101000000: data <= 32'h37ddac5a;
    11'b01101000001: data <= 32'h3d8b3e7d;
    11'b01101000010: data <= 32'h36393f6c;
    11'b01101000011: data <= 32'hbb3939f0;
    11'b01101000100: data <= 32'hbc323411;
    11'b01101000101: data <= 32'hb84a3c88;
    11'b01101000110: data <= 32'hb4953e85;
    11'b01101000111: data <= 32'h2be43451;
    11'b01101001000: data <= 32'h3c76be6b;
    11'b01101001001: data <= 32'h4022be73;
    11'b01101001010: data <= 32'h3eb33237;
    11'b01101001011: data <= 32'h36e73dbe;
    11'b01101001100: data <= 32'h22503a5d;
    11'b01101001101: data <= 32'h38d1b803;
    11'b01101001110: data <= 32'h380bbbd0;
    11'b01101001111: data <= 32'hbc06bb93;
    11'b01101010000: data <= 32'hc047bd3a;
    11'b01101010001: data <= 32'hbc6ebe7d;
    11'b01101010010: data <= 32'h3bddbb85;
    11'b01101010011: data <= 32'h3df2346f;
    11'b01101010100: data <= 32'haec33992;
    11'b01101010101: data <= 32'hbe9a357f;
    11'b01101010110: data <= 32'hbe40389c;
    11'b01101010111: data <= 32'hb9d73e61;
    11'b01101011000: data <= 32'hb8693eed;
    11'b01101011001: data <= 32'hb9752e3d;
    11'b01101011010: data <= 32'ha715be20;
    11'b01101011011: data <= 32'h3c6fbbc6;
    11'b01101011100: data <= 32'h3def3c94;
    11'b01101011101: data <= 32'h3c29404d;
    11'b01101011110: data <= 32'h3b063c34;
    11'b01101011111: data <= 32'h3c89b61b;
    11'b01101100000: data <= 32'h3905b838;
    11'b01101100001: data <= 32'hbac6b06b;
    11'b01101100010: data <= 32'hbe1bb935;
    11'b01101100011: data <= 32'hb12dbecd;
    11'b01101100100: data <= 32'h3ee7bf53;
    11'b01101100101: data <= 32'h3eb1bb45;
    11'b01101100110: data <= 32'hb412b08e;
    11'b01101100111: data <= 32'hbe7a29e1;
    11'b01101101000: data <= 32'hbcae3745;
    11'b01101101001: data <= 32'hb62d3cba;
    11'b01101101010: data <= 32'hbaca3bfe;
    11'b01101101011: data <= 32'hbf0eb7ee;
    11'b01101101100: data <= 32'hbd99be3a;
    11'b01101101101: data <= 32'h3058b831;
    11'b01101101110: data <= 32'h3cbf3e34;
    11'b01101101111: data <= 32'h3c6b405c;
    11'b01101110000: data <= 32'h3a5e3bb4;
    11'b01101110001: data <= 32'h3a0e02c6;
    11'b01101110010: data <= 32'h34e9388d;
    11'b01101110011: data <= 32'hb9593cfb;
    11'b01101110100: data <= 32'hbaac34a4;
    11'b01101110101: data <= 32'h38adbe41;
    11'b01101110110: data <= 32'h402dc06d;
    11'b01101110111: data <= 32'h3ef7bcf8;
    11'b01101111000: data <= 32'h2abdb141;
    11'b01101111001: data <= 32'hb9bc2ce5;
    11'b01101111010: data <= 32'h280e2e98;
    11'b01101111011: data <= 32'h363f35b2;
    11'b01101111100: data <= 32'hbba62da8;
    11'b01101111101: data <= 32'hc10bbc11;
    11'b01101111110: data <= 32'hc056be93;
    11'b01101111111: data <= 32'hb3dfb8fb;
    11'b01110000000: data <= 32'h3c113c09;
    11'b01110000001: data <= 32'h39983d4c;
    11'b01110000010: data <= 32'ha223370c;
    11'b01110000011: data <= 32'hb0263582;
    11'b01110000100: data <= 32'hb1b23e95;
    11'b01110000101: data <= 32'hb90240c2;
    11'b01110000110: data <= 32'hb9143b7e;
    11'b01110000111: data <= 32'h3796bd5b;
    11'b01110001000: data <= 32'h3e9abfbe;
    11'b01110001001: data <= 32'h3dffb90b;
    11'b01110001010: data <= 32'h387b384f;
    11'b01110001011: data <= 32'h382b3622;
    11'b01110001100: data <= 32'h3d76b18a;
    11'b01110001101: data <= 32'h3ca7b1b7;
    11'b01110001110: data <= 32'hba8bb2b6;
    11'b01110001111: data <= 32'hc116bb9b;
    11'b01110010000: data <= 32'hbfb1be7b;
    11'b01110010001: data <= 32'h30f7bcb5;
    11'b01110010010: data <= 32'h3c60b261;
    11'b01110010011: data <= 32'h31e41e5f;
    11'b01110010100: data <= 32'hbac2b4aa;
    11'b01110010101: data <= 32'hb9f73667;
    11'b01110010110: data <= 32'hb59b401e;
    11'b01110010111: data <= 32'hb9674134;
    11'b01110011000: data <= 32'hbc583b30;
    11'b01110011001: data <= 32'hb83fbcda;
    11'b01110011010: data <= 32'h3854bd24;
    11'b01110011011: data <= 32'h3bb035ee;
    11'b01110011100: data <= 32'h3afe3d56;
    11'b01110011101: data <= 32'h3d4c3916;
    11'b01110011110: data <= 32'h4015b331;
    11'b01110011111: data <= 32'h3dde2116;
    11'b01110100000: data <= 32'hb891375d;
    11'b01110100001: data <= 32'hbfb1b11a;
    11'b01110100010: data <= 32'hbbaabd6a;
    11'b01110100011: data <= 32'h3ba2bf05;
    11'b01110100100: data <= 32'h3d27bd3e;
    11'b01110100101: data <= 32'hae24bbfc;
    11'b01110100110: data <= 32'hbc29ba8f;
    11'b01110100111: data <= 32'hb7d930cd;
    11'b01110101000: data <= 32'h2ecc3e8c;
    11'b01110101001: data <= 32'hb9283f89;
    11'b01110101010: data <= 32'hbf653477;
    11'b01110101011: data <= 32'hbf46bd00;
    11'b01110101100: data <= 32'hb8e9b9ea;
    11'b01110101101: data <= 32'h36333bc4;
    11'b01110101110: data <= 32'h3a233dff;
    11'b01110101111: data <= 32'h3ceb3765;
    11'b01110110000: data <= 32'h3edab09b;
    11'b01110110001: data <= 32'h3ca33a57;
    11'b01110110010: data <= 32'hb6593f01;
    11'b01110110011: data <= 32'hbca43bc4;
    11'b01110110100: data <= 32'haa3ebb3d;
    11'b01110110101: data <= 32'h3dccbfb4;
    11'b01110110110: data <= 32'h3d32be7f;
    11'b01110110111: data <= 32'hab3bbc6b;
    11'b01110111000: data <= 32'hb706bacd;
    11'b01110111001: data <= 32'h38e6b2e8;
    11'b01110111010: data <= 32'h3c493a17;
    11'b01110111011: data <= 32'hb6ad3abb;
    11'b01110111100: data <= 32'hc0bab5e6;
    11'b01110111101: data <= 32'hc11ebd3a;
    11'b01110111110: data <= 32'hbc76b8da;
    11'b01110111111: data <= 32'h2e9239b6;
    11'b01111000000: data <= 32'h35163a00;
    11'b01111000001: data <= 32'h3630b3ab;
    11'b01111000010: data <= 32'h39d7b09d;
    11'b01111000011: data <= 32'h387d3e69;
    11'b01111000100: data <= 32'hb58e41b4;
    11'b01111000101: data <= 32'hba213f14;
    11'b01111000110: data <= 32'h2ef9b814;
    11'b01111000111: data <= 32'h3c84be45;
    11'b01111001000: data <= 32'h3b2bbbe4;
    11'b01111001001: data <= 32'h2ef4b57f;
    11'b01111001010: data <= 32'h382ab746;
    11'b01111001011: data <= 32'h3fa5b7c4;
    11'b01111001100: data <= 32'h400c2c49;
    11'b01111001101: data <= 32'hab8434b6;
    11'b01111001110: data <= 32'hc088b6f0;
    11'b01111001111: data <= 32'hc096bc99;
    11'b01111010000: data <= 32'hb992baa6;
    11'b01111010001: data <= 32'h336eb2ac;
    11'b01111010010: data <= 32'hb20fb839;
    11'b01111010011: data <= 32'hb89abcb2;
    11'b01111010100: data <= 32'haf34b5a2;
    11'b01111010101: data <= 32'h33e13f76;
    11'b01111010110: data <= 32'hb4bc421f;
    11'b01111010111: data <= 32'hbb483f06;
    11'b01111011000: data <= 32'hb8dab648;
    11'b01111011001: data <= 32'h2c73bb4f;
    11'b01111011010: data <= 32'h309f2fa8;
    11'b01111011011: data <= 32'h2fee3938;
    11'b01111011100: data <= 32'h3c93ab16;
    11'b01111011101: data <= 32'h4129b8d6;
    11'b01111011110: data <= 32'h40cca5fc;
    11'b01111011111: data <= 32'h33643968;
    11'b01111100000: data <= 32'hbe7f34ac;
    11'b01111100001: data <= 32'hbcf8b95d;
    11'b01111100010: data <= 32'h3465bc57;
    11'b01111100011: data <= 32'h388fbc75;
    11'b01111100100: data <= 32'hb816be22;
    11'b01111100101: data <= 32'hbc13bf46;
    11'b01111100110: data <= 32'hb084b997;
    11'b01111100111: data <= 32'h38f03d96;
    11'b01111101000: data <= 32'hac54408c;
    11'b01111101001: data <= 32'hbd5b3bfe;
    11'b01111101010: data <= 32'hbeacb878;
    11'b01111101011: data <= 32'hbc5cb582;
    11'b01111101100: data <= 32'hb8b53b87;
    11'b01111101101: data <= 32'hb0543c61;
    11'b01111101110: data <= 32'h3bd0afde;
    11'b01111101111: data <= 32'h4068b994;
    11'b01111110000: data <= 32'h3ff936d8;
    11'b01111110001: data <= 32'h34cc3ee6;
    11'b01111110010: data <= 32'hbac63db3;
    11'b01111110011: data <= 32'hb059a773;
    11'b01111110100: data <= 32'h3c27bc37;
    11'b01111110101: data <= 32'h39a5bd51;
    11'b01111110110: data <= 32'hb8eebe73;
    11'b01111110111: data <= 32'hb9eabf35;
    11'b01111111000: data <= 32'h39aabbf6;
    11'b01111111001: data <= 32'h3e4f3813;
    11'b01111111010: data <= 32'h35f63c3b;
    11'b01111111011: data <= 32'hbe6f2df1;
    11'b01111111100: data <= 32'hc091ba0e;
    11'b01111111101: data <= 32'hbe56ae14;
    11'b01111111110: data <= 32'hbb0c3bef;
    11'b01111111111: data <= 32'hb87d38de;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    