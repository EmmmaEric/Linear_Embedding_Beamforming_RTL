
module memory_rom_42(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hb7e13e03;
    11'b00000000001: data <= 32'hb3373b0d;
    11'b00000000010: data <= 32'h3506bae4;
    11'b00000000011: data <= 32'h3d43bd55;
    11'b00000000100: data <= 32'h3ebd35dc;
    11'b00000000101: data <= 32'h3b8c404e;
    11'b00000000110: data <= 32'h34083f5d;
    11'b00000000111: data <= 32'h38562b88;
    11'b00000001000: data <= 32'h3adfbc2d;
    11'b00000001001: data <= 32'ha797bb8a;
    11'b00000001010: data <= 32'hbcfbbb2f;
    11'b00000001011: data <= 32'hba8bbdbf;
    11'b00000001100: data <= 32'h3c7abe2f;
    11'b00000001101: data <= 32'h4020b959;
    11'b00000001110: data <= 32'h38b63231;
    11'b00000001111: data <= 32'hbe64321d;
    11'b00000010000: data <= 32'hc03f2ab2;
    11'b00000010001: data <= 32'hbc923901;
    11'b00000010010: data <= 32'hb89f3c53;
    11'b00000010011: data <= 32'hbbcd316b;
    11'b00000010100: data <= 32'hbbf3bd3a;
    11'b00000010101: data <= 32'h2c7abc96;
    11'b00000010110: data <= 32'h3c603bbb;
    11'b00000010111: data <= 32'h3c31414a;
    11'b00000011000: data <= 32'h386a400b;
    11'b00000011001: data <= 32'h382c345a;
    11'b00000011010: data <= 32'h380eb53c;
    11'b00000011011: data <= 32'hb38e3471;
    11'b00000011100: data <= 32'hbb063402;
    11'b00000011101: data <= 32'h25fcbbf0;
    11'b00000011110: data <= 32'h3fabbfa0;
    11'b00000011111: data <= 32'h40edbd5e;
    11'b00000100000: data <= 32'h3a56b2a8;
    11'b00000100001: data <= 32'hbc6731f7;
    11'b00000100010: data <= 32'hbcc02a38;
    11'b00000100011: data <= 32'hb3963176;
    11'b00000100100: data <= 32'hb5c83185;
    11'b00000100101: data <= 32'hbe87b9d8;
    11'b00000100110: data <= 32'hc016bf0d;
    11'b00000100111: data <= 32'hb9a2bcdf;
    11'b00000101000: data <= 32'h3aaa3a8e;
    11'b00000101001: data <= 32'h3bac4048;
    11'b00000101010: data <= 32'h30dd3dda;
    11'b00000101011: data <= 32'hb47434ab;
    11'b00000101100: data <= 32'hb4b73871;
    11'b00000101101: data <= 32'hb8a23e6e;
    11'b00000101110: data <= 32'hb9c93d26;
    11'b00000101111: data <= 32'h344bb8ee;
    11'b00000110000: data <= 32'h3f83bfa0;
    11'b00000110001: data <= 32'h408bbcb0;
    11'b00000110010: data <= 32'h3bf9353e;
    11'b00000110011: data <= 32'hb07e3a08;
    11'b00000110100: data <= 32'h336f3183;
    11'b00000110101: data <= 32'h3b2ab407;
    11'b00000110110: data <= 32'ha189b6d8;
    11'b00000110111: data <= 32'hbf78bc54;
    11'b00000111000: data <= 32'hc084bf70;
    11'b00000111001: data <= 32'hb866be05;
    11'b00000111010: data <= 32'h3c73aa90;
    11'b00000111011: data <= 32'h3aea3acd;
    11'b00000111100: data <= 32'hb7e436df;
    11'b00000111101: data <= 32'hbc8b2d92;
    11'b00000111110: data <= 32'hbb1a3c63;
    11'b00000111111: data <= 32'hba6d408a;
    11'b00001000000: data <= 32'hbb8e3e42;
    11'b00001000001: data <= 32'hb5c8b8fc;
    11'b00001000010: data <= 32'h3b25bec2;
    11'b00001000011: data <= 32'h3e01b726;
    11'b00001000100: data <= 32'h3c163d27;
    11'b00001000101: data <= 32'h39923db3;
    11'b00001000110: data <= 32'h3d2b3598;
    11'b00001000111: data <= 32'h3e39b410;
    11'b00001001000: data <= 32'h31d7b110;
    11'b00001001001: data <= 32'hbeb0b7da;
    11'b00001001010: data <= 32'hbe9dbdae;
    11'b00001001011: data <= 32'h3518bf1a;
    11'b00001001100: data <= 32'h3ed8bc6f;
    11'b00001001101: data <= 32'h3b03b75d;
    11'b00001001110: data <= 32'hba8fb763;
    11'b00001001111: data <= 32'hbd2cb1c4;
    11'b00001010000: data <= 32'hb9993c40;
    11'b00001010001: data <= 32'hb9363fe4;
    11'b00001010010: data <= 32'hbd843bd7;
    11'b00001010011: data <= 32'hbe0bbc1a;
    11'b00001010100: data <= 32'hb7ccbe00;
    11'b00001010101: data <= 32'h389f3257;
    11'b00001010110: data <= 32'h3abc3f69;
    11'b00001010111: data <= 32'h3b7f3e56;
    11'b00001011000: data <= 32'h3da335e5;
    11'b00001011001: data <= 32'h3d7b31d5;
    11'b00001011010: data <= 32'h29db3b44;
    11'b00001011011: data <= 32'hbd3f3a46;
    11'b00001011100: data <= 32'hba6eb915;
    11'b00001011101: data <= 32'h3ca5bf4a;
    11'b00001011110: data <= 32'h4034becd;
    11'b00001011111: data <= 32'h3b6ebc0d;
    11'b00001100000: data <= 32'hb885b968;
    11'b00001100001: data <= 32'hb803b4a3;
    11'b00001100010: data <= 32'h351b38ee;
    11'b00001100011: data <= 32'hae733c59;
    11'b00001100100: data <= 32'hbed42bcb;
    11'b00001100101: data <= 32'hc0ecbdee;
    11'b00001100110: data <= 32'hbdb1bdd8;
    11'b00001100111: data <= 32'h2c11340c;
    11'b00001101000: data <= 32'h38d33dec;
    11'b00001101001: data <= 32'h384f3b6c;
    11'b00001101010: data <= 32'h39502c8a;
    11'b00001101011: data <= 32'h38a639df;
    11'b00001101100: data <= 32'hb4d34041;
    11'b00001101101: data <= 32'hbc573ff5;
    11'b00001101110: data <= 32'hb6582809;
    11'b00001101111: data <= 32'h3cfdbe82;
    11'b00001110000: data <= 32'h3f58be12;
    11'b00001110001: data <= 32'h3abfb87b;
    11'b00001110010: data <= 32'h2cc0b127;
    11'b00001110011: data <= 32'h3a6cb178;
    11'b00001110100: data <= 32'h3e8130e4;
    11'b00001110101: data <= 32'h389035d5;
    11'b00001110110: data <= 32'hbed5b678;
    11'b00001110111: data <= 32'hc14bbe20;
    11'b00001111000: data <= 32'hbd82bdfa;
    11'b00001111001: data <= 32'h33dcb504;
    11'b00001111010: data <= 32'h37b434ef;
    11'b00001111011: data <= 32'hb013b478;
    11'b00001111100: data <= 32'hb474b799;
    11'b00001111101: data <= 32'haf2b3c0a;
    11'b00001111110: data <= 32'hb8064180;
    11'b00001111111: data <= 32'hbc6140cd;
    11'b00010000000: data <= 32'hb9f7316f;
    11'b00010000001: data <= 32'h3622bd68;
    11'b00010000010: data <= 32'h3b34ba40;
    11'b00010000011: data <= 32'h38263735;
    11'b00010000100: data <= 32'h38fa38b9;
    11'b00010000101: data <= 32'h3f3f1c0e;
    11'b00010000110: data <= 32'h40e3a469;
    11'b00010000111: data <= 32'h3baa361d;
    11'b00010001000: data <= 32'hbdab2bb5;
    11'b00010001001: data <= 32'hc011bb92;
    11'b00010001010: data <= 32'hb7e2bdad;
    11'b00010001011: data <= 32'h3b2ebc45;
    11'b00010001100: data <= 32'h3803bb8e;
    11'b00010001101: data <= 32'hb8a9bd69;
    11'b00010001110: data <= 32'hb940bbe1;
    11'b00010001111: data <= 32'haaeb3ab9;
    11'b00010010000: data <= 32'hb37640e2;
    11'b00010010001: data <= 32'hbcd03f55;
    11'b00010010010: data <= 32'hbe59b40b;
    11'b00010010011: data <= 32'hbb73bcad;
    11'b00010010100: data <= 32'hb31fa8fb;
    11'b00010010101: data <= 32'h2a993cd1;
    11'b00010010110: data <= 32'h39833b0b;
    11'b00010010111: data <= 32'h3fadac24;
    11'b00010011000: data <= 32'h40a02fc6;
    11'b00010011001: data <= 32'h3abe3c95;
    11'b00010011010: data <= 32'hbc363d0a;
    11'b00010011011: data <= 32'hbc7129ca;
    11'b00010011100: data <= 32'h3816bc94;
    11'b00010011101: data <= 32'h3dacbdcd;
    11'b00010011110: data <= 32'h37efbdf1;
    11'b00010011111: data <= 32'hb8b9bea6;
    11'b00010100000: data <= 32'hb0fabcaa;
    11'b00010100001: data <= 32'h3b0a35ee;
    11'b00010100010: data <= 32'h38273e03;
    11'b00010100011: data <= 32'hbcc23a45;
    11'b00010100100: data <= 32'hc099baa9;
    11'b00010100101: data <= 32'hbf6abc65;
    11'b00010100110: data <= 32'hbafa33cd;
    11'b00010100111: data <= 32'hb5063c6f;
    11'b00010101000: data <= 32'h33a5351e;
    11'b00010101001: data <= 32'h3c8ab865;
    11'b00010101010: data <= 32'h3db7353e;
    11'b00010101011: data <= 32'h36314037;
    11'b00010101100: data <= 32'hba8540e6;
    11'b00010101101: data <= 32'hb8123b0f;
    11'b00010101110: data <= 32'h3adeba24;
    11'b00010101111: data <= 32'h3d0bbcba;
    11'b00010110000: data <= 32'h33dcbc06;
    11'b00010110001: data <= 32'hb4a5bc5e;
    11'b00010110010: data <= 32'h3b0bbbb7;
    11'b00010110011: data <= 32'h4055adf5;
    11'b00010110100: data <= 32'h3d8d38ed;
    11'b00010110101: data <= 32'hbbab2c9e;
    11'b00010110110: data <= 32'hc0bbbc06;
    11'b00010110111: data <= 32'hbf2abbf7;
    11'b00010111000: data <= 32'hb9701675;
    11'b00010111001: data <= 32'hb64532ba;
    11'b00010111010: data <= 32'hb6d8bae6;
    11'b00010111011: data <= 32'h2b5dbd3e;
    11'b00010111100: data <= 32'h3811354b;
    11'b00010111101: data <= 32'h2a094128;
    11'b00010111110: data <= 32'hb9c441b5;
    11'b00010111111: data <= 32'hb86f3c3b;
    11'b00011000000: data <= 32'h345cb7cf;
    11'b00011000001: data <= 32'h35c9b6ec;
    11'b00011000010: data <= 32'hb4db2f51;
    11'b00011000011: data <= 32'ha9b6b073;
    11'b00011000100: data <= 32'h3edbb929;
    11'b00011000101: data <= 32'h41fab55c;
    11'b00011000110: data <= 32'h3f7235af;
    11'b00011000111: data <= 32'hb8e23419;
    11'b00011001000: data <= 32'hbee1b797;
    11'b00011001001: data <= 32'hba8ab99a;
    11'b00011001010: data <= 32'h3089b6e4;
    11'b00011001011: data <= 32'hb378bac5;
    11'b00011001100: data <= 32'hbb6fbfcd;
    11'b00011001101: data <= 32'hb892bfd0;
    11'b00011001110: data <= 32'h34922a81;
    11'b00011001111: data <= 32'h33ab406e;
    11'b00011010000: data <= 32'hb901406f;
    11'b00011010001: data <= 32'hbc433807;
    11'b00011010010: data <= 32'hba9fb6d1;
    11'b00011010011: data <= 32'hba433572;
    11'b00011010100: data <= 32'hbb8e3c5f;
    11'b00011010101: data <= 32'hb07836d9;
    11'b00011010110: data <= 32'h3efab8e6;
    11'b00011010111: data <= 32'h41a0b5f9;
    11'b00011011000: data <= 32'h3ea23a52;
    11'b00011011001: data <= 32'hb56c3ce7;
    11'b00011011010: data <= 32'hba2b384a;
    11'b00011011011: data <= 32'h3637b30e;
    11'b00011011100: data <= 32'h3b73b8d5;
    11'b00011011101: data <= 32'haf79bd29;
    11'b00011011110: data <= 32'hbc56c07a;
    11'b00011011111: data <= 32'hb63dc032;
    11'b00011100000: data <= 32'h3bcdb5d2;
    11'b00011100001: data <= 32'h3c003d01;
    11'b00011100010: data <= 32'hb6373be7;
    11'b00011100011: data <= 32'hbe1fb554;
    11'b00011100100: data <= 32'hbe87b7e1;
    11'b00011100101: data <= 32'hbdbf39f1;
    11'b00011100110: data <= 32'hbd533d37;
    11'b00011100111: data <= 32'hb8a53000;
    11'b00011101000: data <= 32'h3b71bc58;
    11'b00011101001: data <= 32'h3f17b652;
    11'b00011101010: data <= 32'h3bba3de8;
    11'b00011101011: data <= 32'hb3d1408e;
    11'b00011101100: data <= 32'hacaa3d98;
    11'b00011101101: data <= 32'h3c1e3387;
    11'b00011101110: data <= 32'h3c2eb4b3;
    11'b00011101111: data <= 32'hb556ba2d;
    11'b00011110000: data <= 32'hbc05be2c;
    11'b00011110001: data <= 32'h35a8bec5;
    11'b00011110010: data <= 32'h4036b980;
    11'b00011110011: data <= 32'h3fa23497;
    11'b00011110100: data <= 32'ha78a9d9b;
    11'b00011110101: data <= 32'hbe02ba51;
    11'b00011110110: data <= 32'hbe13b730;
    11'b00011110111: data <= 32'hbc9c39a9;
    11'b00011111000: data <= 32'hbcfe39ac;
    11'b00011111001: data <= 32'hbc7fbb14;
    11'b00011111010: data <= 32'hb2c1bf94;
    11'b00011111011: data <= 32'h38b0b878;
    11'b00011111100: data <= 32'h35563f3c;
    11'b00011111101: data <= 32'hb3a0413c;
    11'b00011111110: data <= 32'h2c7a3e12;
    11'b00011111111: data <= 32'h3a093684;
    11'b00100000000: data <= 32'h356435c9;
    11'b00100000001: data <= 32'hbb6a3678;
    11'b00100000010: data <= 32'hbba4b584;
    11'b00100000011: data <= 32'h3c0abc52;
    11'b00100000100: data <= 32'h41b6ba88;
    11'b00100000101: data <= 32'h40b7b080;
    11'b00100000110: data <= 32'h344bb066;
    11'b00100000111: data <= 32'hbb4db794;
    11'b00100001000: data <= 32'hb7e1afcc;
    11'b00100001001: data <= 32'haf1137d3;
    11'b00100001010: data <= 32'hba77b079;
    11'b00100001011: data <= 32'hbdfcbf8f;
    11'b00100001100: data <= 32'hbbe2c117;
    11'b00100001101: data <= 32'h29c1bac3;
    11'b00100001110: data <= 32'h34893dd8;
    11'b00100001111: data <= 32'hb0413fb8;
    11'b00100010000: data <= 32'hb30c3a2d;
    11'b00100010001: data <= 32'haf1232c9;
    11'b00100010010: data <= 32'hb9b43c01;
    11'b00100010011: data <= 32'hbe6b3e0b;
    11'b00100010100: data <= 32'hbc713850;
    11'b00100010101: data <= 32'h3c0fba3b;
    11'b00100010110: data <= 32'h4141baaf;
    11'b00100010111: data <= 32'h40002cdb;
    11'b00100011000: data <= 32'h35153894;
    11'b00100011001: data <= 32'hadaa36cd;
    11'b00100011010: data <= 32'h3aa036a4;
    11'b00100011011: data <= 32'h3bec36ca;
    11'b00100011100: data <= 32'hb677b827;
    11'b00100011101: data <= 32'hbe69c043;
    11'b00100011110: data <= 32'hbc0dc127;
    11'b00100011111: data <= 32'h3746bc54;
    11'b00100100000: data <= 32'h3b4338d3;
    11'b00100100001: data <= 32'h315b38c2;
    11'b00100100010: data <= 32'hb84bb5dd;
    11'b00100100011: data <= 32'hba81b0ea;
    11'b00100100100: data <= 32'hbd4a3d52;
    11'b00100100101: data <= 32'hbfb23fac;
    11'b00100100110: data <= 32'hbdb43844;
    11'b00100100111: data <= 32'h348fbc5a;
    11'b00100101000: data <= 32'h3df8bb50;
    11'b00100101001: data <= 32'h3c1638b0;
    11'b00100101010: data <= 32'h2f1f3df4;
    11'b00100101011: data <= 32'h38243cf9;
    11'b00100101100: data <= 32'h3ea03ac6;
    11'b00100101101: data <= 32'h3dab3954;
    11'b00100101110: data <= 32'hb6c9ab51;
    11'b00100101111: data <= 32'hbe41bd69;
    11'b00100110000: data <= 32'hb764bfa6;
    11'b00100110001: data <= 32'h3dadbc75;
    11'b00100110010: data <= 32'h3f10b41f;
    11'b00100110011: data <= 32'h3851b89e;
    11'b00100110100: data <= 32'hb829bc9b;
    11'b00100110101: data <= 32'hb9cdb56d;
    11'b00100110110: data <= 32'hbbc43d42;
    11'b00100110111: data <= 32'hbe7b3e1a;
    11'b00100111000: data <= 32'hbeceb480;
    11'b00100111001: data <= 32'hb9ffbf55;
    11'b00100111010: data <= 32'h3056bc79;
    11'b00100111011: data <= 32'h2a693b09;
    11'b00100111100: data <= 32'hb08e3f4b;
    11'b00100111101: data <= 32'h39403d3b;
    11'b00100111110: data <= 32'h3e5c3abf;
    11'b00100111111: data <= 32'h3b773c5c;
    11'b00101000000: data <= 32'hbb7e3c11;
    11'b00101000001: data <= 32'hbe471c83;
    11'b00101000010: data <= 32'h2f5ebba8;
    11'b00101000011: data <= 32'h4044bbaa;
    11'b00101000100: data <= 32'h4059b942;
    11'b00101000101: data <= 32'h39b0bb62;
    11'b00101000110: data <= 32'haf67bc5c;
    11'b00101000111: data <= 32'h32c9afa2;
    11'b00101001000: data <= 32'h32e83ca1;
    11'b00101001001: data <= 32'hbac53a52;
    11'b00101001010: data <= 32'hbf19bce5;
    11'b00101001011: data <= 32'hbde6c0e9;
    11'b00101001100: data <= 32'hb8f9bd4d;
    11'b00101001101: data <= 32'hb49a3958;
    11'b00101001110: data <= 32'hb1bb3cd3;
    11'b00101001111: data <= 32'h36ca36f7;
    11'b00101010000: data <= 32'h3aee3561;
    11'b00101010001: data <= 32'ha6e43dba;
    11'b00101010010: data <= 32'hbe5e401e;
    11'b00101010011: data <= 32'hbec23c6b;
    11'b00101010100: data <= 32'h32a5b569;
    11'b00101010101: data <= 32'h3fd6ba5f;
    11'b00101010110: data <= 32'h3ed6b7ca;
    11'b00101010111: data <= 32'h37adb60f;
    11'b00101011000: data <= 32'h36c4b503;
    11'b00101011001: data <= 32'h3dd9364e;
    11'b00101011010: data <= 32'h3e1f3c61;
    11'b00101011011: data <= 32'hae7835e6;
    11'b00101011100: data <= 32'hbea6be04;
    11'b00101011101: data <= 32'hbe1ec0ce;
    11'b00101011110: data <= 32'hb65ebd49;
    11'b00101011111: data <= 32'h31b22c94;
    11'b00101100000: data <= 32'h2d6dab72;
    11'b00101100001: data <= 32'h3065bb4c;
    11'b00101100010: data <= 32'h3146b626;
    11'b00101100011: data <= 32'hb9453e0b;
    11'b00101100100: data <= 32'hbf6a40f4;
    11'b00101100101: data <= 32'hbf3e3d34;
    11'b00101100110: data <= 32'hb4adb72d;
    11'b00101100111: data <= 32'h3b23ba82;
    11'b00101101000: data <= 32'h383fa5ab;
    11'b00101101001: data <= 32'had7d37f2;
    11'b00101101010: data <= 32'h3a13380f;
    11'b00101101011: data <= 32'h40923a58;
    11'b00101101100: data <= 32'h405a3cc5;
    11'b00101101101: data <= 32'h2f8d3918;
    11'b00101101110: data <= 32'hbe1eba55;
    11'b00101101111: data <= 32'hbc1ebe37;
    11'b00101110000: data <= 32'h37ddbc02;
    11'b00101110001: data <= 32'h3c0db813;
    11'b00101110010: data <= 32'h370fbcdd;
    11'b00101110011: data <= 32'h2b99bfb8;
    11'b00101110100: data <= 32'h2e57baca;
    11'b00101110101: data <= 32'hb5ef3d76;
    11'b00101110110: data <= 32'hbd924043;
    11'b00101110111: data <= 32'hbf0638bd;
    11'b00101111000: data <= 32'hbc2fbc91;
    11'b00101111001: data <= 32'hb718bc08;
    11'b00101111010: data <= 32'hb97e352f;
    11'b00101111011: data <= 32'hb93c3b8e;
    11'b00101111100: data <= 32'h39dd3910;
    11'b00101111101: data <= 32'h40863951;
    11'b00101111110: data <= 32'h3f4e3d49;
    11'b00101111111: data <= 32'hb4ea3dc3;
    11'b00110000000: data <= 32'hbe15384d;
    11'b00110000001: data <= 32'hb6e7b591;
    11'b00110000010: data <= 32'h3d1eb801;
    11'b00110000011: data <= 32'h3de8b9b0;
    11'b00110000100: data <= 32'h382abe67;
    11'b00110000101: data <= 32'h32c2c012;
    11'b00110000110: data <= 32'h3a47ba0e;
    11'b00110000111: data <= 32'h3a3f3cb8;
    11'b00110001000: data <= 32'hb5f73d98;
    11'b00110001001: data <= 32'hbdddb640;
    11'b00110001010: data <= 32'hbe2ebf3c;
    11'b00110001011: data <= 32'hbcf0bc9d;
    11'b00110001100: data <= 32'hbce6351c;
    11'b00110001101: data <= 32'hbaee386d;
    11'b00110001110: data <= 32'h3733b260;
    11'b00110001111: data <= 32'h3e3bacb1;
    11'b00110010000: data <= 32'h3ae23d2f;
    11'b00110010001: data <= 32'hbbf74079;
    11'b00110010010: data <= 32'hbe6a3eaa;
    11'b00110010011: data <= 32'hb19f3802;
    11'b00110010100: data <= 32'h3d38af46;
    11'b00110010101: data <= 32'h3c3bb758;
    11'b00110010110: data <= 32'h2d4abc5a;
    11'b00110010111: data <= 32'h3656bd29;
    11'b00110011000: data <= 32'h3f20b367;
    11'b00110011001: data <= 32'h403d3c65;
    11'b00110011010: data <= 32'h39023ad5;
    11'b00110011011: data <= 32'hbc53babf;
    11'b00110011100: data <= 32'hbdf1bf3f;
    11'b00110011101: data <= 32'hbc35bbc8;
    11'b00110011110: data <= 32'hbaa52aec;
    11'b00110011111: data <= 32'hb8fab75a;
    11'b00110100000: data <= 32'h30e0be43;
    11'b00110100001: data <= 32'h3a28bc40;
    11'b00110100010: data <= 32'h2d3c3c43;
    11'b00110100011: data <= 32'hbd494104;
    11'b00110100100: data <= 32'hbe553fa3;
    11'b00110100101: data <= 32'hb5fe380a;
    11'b00110100110: data <= 32'h37baac73;
    11'b00110100111: data <= 32'hb03e253a;
    11'b00110101000: data <= 32'hba0fb108;
    11'b00110101001: data <= 32'h3655b5a2;
    11'b00110101010: data <= 32'h40dd33a2;
    11'b00110101011: data <= 32'h41a23c5e;
    11'b00110101100: data <= 32'h3c023ad9;
    11'b00110101101: data <= 32'hbab5b5e2;
    11'b00110101110: data <= 32'hbba2bbb1;
    11'b00110101111: data <= 32'hb039b622;
    11'b00110110000: data <= 32'h2dabb19c;
    11'b00110110001: data <= 32'hb24dbdb4;
    11'b00110110010: data <= 32'h1a30c149;
    11'b00110110011: data <= 32'h379cbee6;
    11'b00110110100: data <= 32'h30953a13;
    11'b00110110101: data <= 32'hbb014038;
    11'b00110110110: data <= 32'hbd193cc4;
    11'b00110110111: data <= 32'hba2fb37c;
    11'b00110111000: data <= 32'hb92eb517;
    11'b00110111001: data <= 32'hbda9369c;
    11'b00110111010: data <= 32'hbe3f37b2;
    11'b00110111011: data <= 32'h311fa2c0;
    11'b00110111100: data <= 32'h40aa30ab;
    11'b00110111101: data <= 32'h40f43bf4;
    11'b00110111110: data <= 32'h38953d40;
    11'b00110111111: data <= 32'hbae039fb;
    11'b00111000000: data <= 32'hb52d34f8;
    11'b00111000001: data <= 32'h3a803627;
    11'b00111000010: data <= 32'h39ffafe1;
    11'b00111000011: data <= 32'habffbed9;
    11'b00111000100: data <= 32'ha892c18e;
    11'b00111000101: data <= 32'h3aa8beb3;
    11'b00111000110: data <= 32'h3c4c388f;
    11'b00111000111: data <= 32'h32883d64;
    11'b00111001000: data <= 32'hb9972d35;
    11'b00111001001: data <= 32'hbbd9bc50;
    11'b00111001010: data <= 32'hbd48b844;
    11'b00111001011: data <= 32'hc0023880;
    11'b00111001100: data <= 32'hbf783650;
    11'b00111001101: data <= 32'hb164b8f8;
    11'b00111001110: data <= 32'h3e62b91a;
    11'b00111001111: data <= 32'h3da5396f;
    11'b00111010000: data <= 32'hb4513f2b;
    11'b00111010001: data <= 32'hbc143ef5;
    11'b00111010010: data <= 32'h2af23ced;
    11'b00111010011: data <= 32'h3c763b5a;
    11'b00111010100: data <= 32'h3872331c;
    11'b00111010101: data <= 32'hb836bca3;
    11'b00111010110: data <= 32'hb033bfd9;
    11'b00111010111: data <= 32'h3dfebc1a;
    11'b00111011000: data <= 32'h40853883;
    11'b00111011001: data <= 32'h3d2939a9;
    11'b00111011010: data <= 32'haf7cb8fd;
    11'b00111011011: data <= 32'hba38bd3b;
    11'b00111011100: data <= 32'hbc58b599;
    11'b00111011101: data <= 32'hbe4a3877;
    11'b00111011110: data <= 32'hbe28b48e;
    11'b00111011111: data <= 32'hb66fbf4b;
    11'b00111100000: data <= 32'h39ddbee4;
    11'b00111100001: data <= 32'h367932c0;
    11'b00111100010: data <= 32'hba933f7b;
    11'b00111100011: data <= 32'hbc153fac;
    11'b00111100100: data <= 32'h2dd43cec;
    11'b00111100101: data <= 32'h38fb3b71;
    11'b00111100110: data <= 32'hb75b394c;
    11'b00111100111: data <= 32'hbddab163;
    11'b00111101000: data <= 32'hb65cba94;
    11'b00111101001: data <= 32'h3facb555;
    11'b00111101010: data <= 32'h41c238d6;
    11'b00111101011: data <= 32'h3ec63805;
    11'b00111101100: data <= 32'h30c7b784;
    11'b00111101101: data <= 32'hb3fdb929;
    11'b00111101110: data <= 32'haf453542;
    11'b00111101111: data <= 32'hb7b338e3;
    11'b00111110000: data <= 32'hbb3dbbed;
    11'b00111110001: data <= 32'hb7c2c19f;
    11'b00111110010: data <= 32'h3431c0e2;
    11'b00111110011: data <= 32'h30edb1a2;
    11'b00111110100: data <= 32'hb8a13dbc;
    11'b00111110101: data <= 32'hb91f3c97;
    11'b00111110110: data <= 32'ha51935a6;
    11'b00111110111: data <= 32'hb33f37f1;
    11'b00111111000: data <= 32'hbe953bd6;
    11'b00111111001: data <= 32'hc0b538f3;
    11'b00111111010: data <= 32'hba25b1e5;
    11'b00111111011: data <= 32'h3ef2b29d;
    11'b00111111100: data <= 32'h40f9375c;
    11'b00111111101: data <= 32'h3ca5396a;
    11'b00111111110: data <= 32'ha55f3590;
    11'b00111111111: data <= 32'h34f5382a;
    11'b01000000000: data <= 32'h3ba83cd1;
    11'b01000000001: data <= 32'h37663ac7;
    11'b01000000010: data <= 32'hb84dbc9e;
    11'b01000000011: data <= 32'hb851c1ca;
    11'b01000000100: data <= 32'h35a3c0a8;
    11'b01000000101: data <= 32'h3a36b42c;
    11'b01000000110: data <= 32'h361039d0;
    11'b01000000111: data <= 32'h2b20aca5;
    11'b01000001000: data <= 32'h9acdba0c;
    11'b01000001001: data <= 32'hb9eb2969;
    11'b01000001010: data <= 32'hc05e3c77;
    11'b01000001011: data <= 32'hc1463a37;
    11'b01000001100: data <= 32'hbc2db7a1;
    11'b01000001101: data <= 32'h3c20baca;
    11'b01000001110: data <= 32'h3d4a26c1;
    11'b01000001111: data <= 32'h2ce83b38;
    11'b01000010000: data <= 32'hb6b03c96;
    11'b01000010001: data <= 32'h39383d92;
    11'b01000010010: data <= 32'h3dee3f0d;
    11'b01000010011: data <= 32'h38b23cc9;
    11'b01000010100: data <= 32'hbab1b8d7;
    11'b01000010101: data <= 32'hb9eebff7;
    11'b01000010110: data <= 32'h39fcbddd;
    11'b01000010111: data <= 32'h3ef7a93f;
    11'b01000011000: data <= 32'h3da73059;
    11'b01000011001: data <= 32'h399fbbd9;
    11'b01000011010: data <= 32'h343abd37;
    11'b01000011011: data <= 32'hb79d28b3;
    11'b01000011100: data <= 32'hbeb63cc9;
    11'b01000011101: data <= 32'hc04435f3;
    11'b01000011110: data <= 32'hbc4dbdbd;
    11'b01000011111: data <= 32'h3323bf7f;
    11'b01000100000: data <= 32'h3026b850;
    11'b01000100001: data <= 32'hba5c3ae6;
    11'b01000100010: data <= 32'hb90d3d0b;
    11'b01000100011: data <= 32'h39fd3d53;
    11'b01000100100: data <= 32'h3d0b3e93;
    11'b01000100101: data <= 32'hb14f3de2;
    11'b01000100110: data <= 32'hbece3557;
    11'b01000100111: data <= 32'hbc7fb973;
    11'b01000101000: data <= 32'h3c03b756;
    11'b01000101001: data <= 32'h40863364;
    11'b01000101010: data <= 32'h3f15ae8a;
    11'b01000101011: data <= 32'h3b1dbc5f;
    11'b01000101100: data <= 32'h3962bb60;
    11'b01000101101: data <= 32'h374d3901;
    11'b01000101110: data <= 32'hb6f53d80;
    11'b01000101111: data <= 32'hbcc9b053;
    11'b01000110000: data <= 32'hbb4ec098;
    11'b01000110001: data <= 32'hb41bc11e;
    11'b01000110010: data <= 32'hb612bb2d;
    11'b01000110011: data <= 32'hbad037d8;
    11'b01000110100: data <= 32'hb5d53819;
    11'b01000110101: data <= 32'h3a193520;
    11'b01000110110: data <= 32'h39183b74;
    11'b01000110111: data <= 32'hbcce3e2c;
    11'b01000111000: data <= 32'hc1213c70;
    11'b01000111001: data <= 32'hbe0d3298;
    11'b01000111010: data <= 32'h3aa7a280;
    11'b01000111011: data <= 32'h3f7a3368;
    11'b01000111100: data <= 32'h3c7fa95f;
    11'b01000111101: data <= 32'h379bb826;
    11'b01000111110: data <= 32'h3c022c66;
    11'b01000111111: data <= 32'h3e043dea;
    11'b01001000000: data <= 32'h39fa3eae;
    11'b01001000001: data <= 32'hb7ecb41e;
    11'b01001000010: data <= 32'hba53c0b7;
    11'b01001000011: data <= 32'hb42fc0b4;
    11'b01001000100: data <= 32'ha31cba40;
    11'b01001000101: data <= 32'hae1fa2d8;
    11'b01001000110: data <= 32'h34dfb974;
    11'b01001000111: data <= 32'h3af9bc0e;
    11'b01001001000: data <= 32'h32be305f;
    11'b01001001001: data <= 32'hbeca3de4;
    11'b01001001010: data <= 32'hc1903d5c;
    11'b01001001011: data <= 32'hbe8d31b8;
    11'b01001001100: data <= 32'h34b5b6c3;
    11'b01001001101: data <= 32'h39d2b11f;
    11'b01001001110: data <= 32'hb1862c6b;
    11'b01001001111: data <= 32'hb42930dc;
    11'b01001010000: data <= 32'h3c793b09;
    11'b01001010001: data <= 32'h40293ffc;
    11'b01001010010: data <= 32'h3c913fb0;
    11'b01001010011: data <= 32'hb8403152;
    11'b01001010100: data <= 32'hbb64bde1;
    11'b01001010101: data <= 32'h2193bd2e;
    11'b01001010110: data <= 32'h3a4cb38a;
    11'b01001010111: data <= 32'h3ad8b5e9;
    11'b01001011000: data <= 32'h3b76be80;
    11'b01001011001: data <= 32'h3c61bf58;
    11'b01001011010: data <= 32'h3651b123;
    11'b01001011011: data <= 32'hbccd3dd0;
    11'b01001011100: data <= 32'hc0373c39;
    11'b01001011101: data <= 32'hbd77b8b3;
    11'b01001011110: data <= 32'hb480bd5c;
    11'b01001011111: data <= 32'hb7d9b9c2;
    11'b01001100000: data <= 32'hbd4725ce;
    11'b01001100001: data <= 32'hba5534c9;
    11'b01001100010: data <= 32'h3c553a90;
    11'b01001100011: data <= 32'h3fe23ef4;
    11'b01001100100: data <= 32'h38d33fb8;
    11'b01001100101: data <= 32'hbd0a3b14;
    11'b01001100110: data <= 32'hbd37b08c;
    11'b01001100111: data <= 32'h330ca234;
    11'b01001101000: data <= 32'h3d303607;
    11'b01001101001: data <= 32'h3cd2b722;
    11'b01001101010: data <= 32'h3c10bf5a;
    11'b01001101011: data <= 32'h3d24bec1;
    11'b01001101100: data <= 32'h3c843428;
    11'b01001101101: data <= 32'h2b113e7b;
    11'b01001101110: data <= 32'hbb3738fc;
    11'b01001101111: data <= 32'hbacdbd97;
    11'b01001110000: data <= 32'hb895c003;
    11'b01001110001: data <= 32'hbc5dbc09;
    11'b01001110010: data <= 32'hbe89b1e4;
    11'b01001110011: data <= 32'hb9d5b489;
    11'b01001110100: data <= 32'h3c45b25e;
    11'b01001110101: data <= 32'h3dc13a33;
    11'b01001110110: data <= 32'hb5873e96;
    11'b01001110111: data <= 32'hc02f3dd0;
    11'b01001111000: data <= 32'hbe9d3a9d;
    11'b01001111001: data <= 32'h312239b1;
    11'b01001111010: data <= 32'h3c2238f8;
    11'b01001111011: data <= 32'h386fb551;
    11'b01001111100: data <= 32'h3607bd79;
    11'b01001111101: data <= 32'h3d19ba89;
    11'b01001111110: data <= 32'h3fd83c44;
    11'b01001111111: data <= 32'h3d3c3f9a;
    11'b01010000000: data <= 32'h2e0536fe;
    11'b01010000001: data <= 32'hb718be36;
    11'b01010000010: data <= 32'hb7e8bf32;
    11'b01010000011: data <= 32'hbab1b99a;
    11'b01010000100: data <= 32'hbc1fb606;
    11'b01010000101: data <= 32'hb025bd10;
    11'b01010000110: data <= 32'h3cb4be64;
    11'b01010000111: data <= 32'h3bf0b531;
    11'b01010001000: data <= 32'hbb383d09;
    11'b01010001001: data <= 32'hc0a03e46;
    11'b01010001010: data <= 32'hbe7c3b4d;
    11'b01010001011: data <= 32'hae9d37d5;
    11'b01010001100: data <= 32'h2dbd3550;
    11'b01010001101: data <= 32'hba66b32b;
    11'b01010001110: data <= 32'hb950b9b6;
    11'b01010001111: data <= 32'h3c32256f;
    11'b01010010000: data <= 32'h40ca3e5d;
    11'b01010010001: data <= 32'h3f444012;
    11'b01010010010: data <= 32'h347c390b;
    11'b01010010011: data <= 32'hb6efbac2;
    11'b01010010100: data <= 32'hb2e9b986;
    11'b01010010101: data <= 32'had323095;
    11'b01010010110: data <= 32'had6fb615;
    11'b01010010111: data <= 32'h380dc017;
    11'b01010011000: data <= 32'h3d4ac110;
    11'b01010011001: data <= 32'h3befbb04;
    11'b01010011010: data <= 32'hb8883c34;
    11'b01010011011: data <= 32'hbe643d09;
    11'b01010011100: data <= 32'hbc4732da;
    11'b01010011101: data <= 32'hb53fb629;
    11'b01010011110: data <= 32'hbba1b347;
    11'b01010011111: data <= 32'hc01fb345;
    11'b01010100000: data <= 32'hbdecb6e0;
    11'b01010100001: data <= 32'h3a402e93;
    11'b01010100010: data <= 32'h40783d3d;
    11'b01010100011: data <= 32'h3d723f2b;
    11'b01010100100: data <= 32'hb5de3c0b;
    11'b01010100101: data <= 32'hba5a34db;
    11'b01010100110: data <= 32'h22e039a5;
    11'b01010100111: data <= 32'h382c3c42;
    11'b01010101000: data <= 32'h361eb1e8;
    11'b01010101001: data <= 32'h38adc05f;
    11'b01010101010: data <= 32'h3d33c0f7;
    11'b01010101011: data <= 32'h3da6b89e;
    11'b01010101100: data <= 32'h38133caf;
    11'b01010101101: data <= 32'hb4893a89;
    11'b01010101110: data <= 32'hb34fb935;
    11'b01010101111: data <= 32'hb508bc93;
    11'b01010110000: data <= 32'hbdd8b836;
    11'b01010110001: data <= 32'hc0f9b43c;
    11'b01010110010: data <= 32'hbe53b9dc;
    11'b01010110011: data <= 32'h3977b9ec;
    11'b01010110100: data <= 32'h3ec833f0;
    11'b01010110101: data <= 32'h363e3cb8;
    11'b01010110110: data <= 32'hbd0f3d00;
    11'b01010110111: data <= 32'hbca63ca5;
    11'b01010111000: data <= 32'h2d363e3b;
    11'b01010111001: data <= 32'h37fb3e13;
    11'b01010111010: data <= 32'hae682adb;
    11'b01010111011: data <= 32'hb058becf;
    11'b01010111100: data <= 32'h3bc4be77;
    11'b01010111101: data <= 32'h3f9e343b;
    11'b01010111110: data <= 32'h3e8c3de3;
    11'b01010111111: data <= 32'h3ad4384f;
    11'b01011000000: data <= 32'h36ecbc08;
    11'b01011000001: data <= 32'hac30bc62;
    11'b01011000010: data <= 32'hbcb9b10f;
    11'b01011000011: data <= 32'hbfabb131;
    11'b01011000100: data <= 32'hbbdcbd82;
    11'b01011000101: data <= 32'h3a72c001;
    11'b01011000110: data <= 32'h3cbcbc00;
    11'b01011000111: data <= 32'hb55737fb;
    11'b01011001000: data <= 32'hbe8a3c99;
    11'b01011001001: data <= 32'hbc603cd5;
    11'b01011001010: data <= 32'h2d253d99;
    11'b01011001011: data <= 32'hafb63d18;
    11'b01011001100: data <= 32'hbd3f3146;
    11'b01011001101: data <= 32'hbd4dbc04;
    11'b01011001110: data <= 32'h36d1b926;
    11'b01011001111: data <= 32'h402a3b6e;
    11'b01011010000: data <= 32'h402e3e60;
    11'b01011010001: data <= 32'h3c88380b;
    11'b01011010010: data <= 32'h384eb8d7;
    11'b01011010011: data <= 32'h33d8b043;
    11'b01011010100: data <= 32'hb6553aa1;
    11'b01011010101: data <= 32'hbaf93157;
    11'b01011010110: data <= 32'hb310bf7e;
    11'b01011010111: data <= 32'h3bb2c1bc;
    11'b01011011000: data <= 32'h3bf6beb0;
    11'b01011011001: data <= 32'hb47b308b;
    11'b01011011010: data <= 32'hbc483a27;
    11'b01011011011: data <= 32'hb69e37bf;
    11'b01011011100: data <= 32'h32143759;
    11'b01011011101: data <= 32'hbae638e4;
    11'b01011011110: data <= 32'hc0fe3069;
    11'b01011011111: data <= 32'hc092b88d;
    11'b01011100000: data <= 32'ha971b4dd;
    11'b01011100001: data <= 32'h3f3c3a6f;
    11'b01011100010: data <= 32'h3e703cf8;
    11'b01011100011: data <= 32'h374b387e;
    11'b01011100100: data <= 32'h2ee73373;
    11'b01011100101: data <= 32'h372a3cb8;
    11'b01011100110: data <= 32'h35333fa8;
    11'b01011100111: data <= 32'hb18638e0;
    11'b01011101000: data <= 32'h2568bf6e;
    11'b01011101001: data <= 32'h3ae3c194;
    11'b01011101010: data <= 32'h3c73bd84;
    11'b01011101011: data <= 32'h37b9349f;
    11'b01011101100: data <= 32'h30e4357e;
    11'b01011101101: data <= 32'h38d7b794;
    11'b01011101110: data <= 32'h37d2b806;
    11'b01011101111: data <= 32'hbcb530aa;
    11'b01011110000: data <= 32'hc1c830b3;
    11'b01011110001: data <= 32'hc0ddb8c8;
    11'b01011110010: data <= 32'hb130bab3;
    11'b01011110011: data <= 32'h3d0eb0ef;
    11'b01011110100: data <= 32'h38803736;
    11'b01011110101: data <= 32'hb8ee37cd;
    11'b01011110110: data <= 32'hb6c23af0;
    11'b01011110111: data <= 32'h38464000;
    11'b01011111000: data <= 32'h385840e8;
    11'b01011111001: data <= 32'hb5ab3b62;
    11'b01011111010: data <= 32'hb8a5bd5d;
    11'b01011111011: data <= 32'h35cabf72;
    11'b01011111100: data <= 32'h3d1ab64d;
    11'b01011111101: data <= 32'h3d7239e7;
    11'b01011111110: data <= 32'h3d082c3a;
    11'b01011111111: data <= 32'h3d91bc28;
    11'b01100000000: data <= 32'h3af4b9f3;
    11'b01100000001: data <= 32'hbaab3613;
    11'b01100000010: data <= 32'hc08a365d;
    11'b01100000011: data <= 32'hbee6bb4d;
    11'b01100000100: data <= 32'h2d87bf55;
    11'b01100000101: data <= 32'h3a1dbd77;
    11'b01100000110: data <= 32'hb57cb63b;
    11'b01100000111: data <= 32'hbd0c3264;
    11'b01100001000: data <= 32'hb8083a86;
    11'b01100001001: data <= 32'h393c3f37;
    11'b01100001010: data <= 32'h33c44049;
    11'b01100001011: data <= 32'hbd263b86;
    11'b01100001100: data <= 32'hbee9b93f;
    11'b01100001101: data <= 32'hb5d7b9da;
    11'b01100001110: data <= 32'h3cdf3841;
    11'b01100001111: data <= 32'h3ebb3c19;
    11'b01100010000: data <= 32'h3e0bab94;
    11'b01100010001: data <= 32'h3dedbb81;
    11'b01100010010: data <= 32'h3c86ac3e;
    11'b01100010011: data <= 32'haaca3d3e;
    11'b01100010100: data <= 32'hbc5c3b5b;
    11'b01100010101: data <= 32'hb9c2bc8d;
    11'b01100010110: data <= 32'h36a9c112;
    11'b01100010111: data <= 32'h3818c00b;
    11'b01100011000: data <= 32'hb893ba41;
    11'b01100011001: data <= 32'hbbe8b1ee;
    11'b01100011010: data <= 32'h2ebb2d27;
    11'b01100011011: data <= 32'h3ba63a01;
    11'b01100011100: data <= 32'hb2943d0d;
    11'b01100011101: data <= 32'hc09139e8;
    11'b01100011110: data <= 32'hc15cb1d6;
    11'b01100011111: data <= 32'hbb56b020;
    11'b01100100000: data <= 32'h3b1239a1;
    11'b01100100001: data <= 32'h3cab3a21;
    11'b01100100010: data <= 32'h39f1b1e6;
    11'b01100100011: data <= 32'h3af5b683;
    11'b01100100100: data <= 32'h3cae3c2a;
    11'b01100100101: data <= 32'h397f40ca;
    11'b01100100110: data <= 32'hb0c53df4;
    11'b01100100111: data <= 32'hb1acbc07;
    11'b01100101000: data <= 32'h36f4c0cb;
    11'b01100101001: data <= 32'h3779bea3;
    11'b01100101010: data <= 32'hafbeb7f4;
    11'b01100101011: data <= 32'h2229b792;
    11'b01100101100: data <= 32'h3c7ebb18;
    11'b01100101101: data <= 32'h3daab6e6;
    11'b01100101110: data <= 32'hb5b437f8;
    11'b01100101111: data <= 32'hc13138d1;
    11'b01100110000: data <= 32'hc18eacd0;
    11'b01100110001: data <= 32'hbb97b59e;
    11'b01100110010: data <= 32'h3707a295;
    11'b01100110011: data <= 32'h2f04a4ca;
    11'b01100110100: data <= 32'hb838b71b;
    11'b01100110101: data <= 32'h2a3125bd;
    11'b01100110110: data <= 32'h3c5e3f09;
    11'b01100110111: data <= 32'h3c0d41d1;
    11'b01100111000: data <= 32'ha67e3f11;
    11'b01100111001: data <= 32'hb823b860;
    11'b01100111010: data <= 32'ha920bdcd;
    11'b01100111011: data <= 32'h36eab7f4;
    11'b01100111100: data <= 32'h38273336;
    11'b01100111101: data <= 32'h3bf7b89c;
    11'b01100111110: data <= 32'h3fa3be24;
    11'b01100111111: data <= 32'h3f45bbbe;
    11'b01101000000: data <= 32'ha5643739;
    11'b01101000001: data <= 32'hbfcb3a6c;
    11'b01101000010: data <= 32'hbfabb235;
    11'b01101000011: data <= 32'hb741bc54;
    11'b01101000100: data <= 32'h2f21bc55;
    11'b01101000101: data <= 32'hbae3bb02;
    11'b01101000110: data <= 32'hbdd6ba73;
    11'b01101000111: data <= 32'hb547ac83;
    11'b01101001000: data <= 32'h3c873e19;
    11'b01101001001: data <= 32'h3b2b40f4;
    11'b01101001010: data <= 32'hb96c3e4c;
    11'b01101001011: data <= 32'hbdffa53c;
    11'b01101001100: data <= 32'hba58b444;
    11'b01101001101: data <= 32'h341539a3;
    11'b01101001110: data <= 32'h3a003a90;
    11'b01101001111: data <= 32'h3ccdb8c0;
    11'b01101010000: data <= 32'h3fa5be67;
    11'b01101010001: data <= 32'h3faab8a8;
    11'b01101010010: data <= 32'h38fd3cc8;
    11'b01101010011: data <= 32'hb9c33d65;
    11'b01101010100: data <= 32'hb931b442;
    11'b01101010101: data <= 32'h3225be9b;
    11'b01101010110: data <= 32'ha063beb8;
    11'b01101010111: data <= 32'hbcf4bcde;
    11'b01101011000: data <= 32'hbdf1bc56;
    11'b01101011001: data <= 32'h2c49b99f;
    11'b01101011010: data <= 32'h3dc936dc;
    11'b01101011011: data <= 32'h38f93d69;
    11'b01101011100: data <= 32'hbe043c3c;
    11'b01101011101: data <= 32'hc0c234d5;
    11'b01101011110: data <= 32'hbd4e377e;
    11'b01101011111: data <= 32'ha80a3cbc;
    11'b01101100000: data <= 32'h34be3a6b;
    11'b01101100001: data <= 32'h3647b9b1;
    11'b01101100010: data <= 32'h3c54bd04;
    11'b01101100011: data <= 32'h3ea23538;
    11'b01101100100: data <= 32'h3ccf4063;
    11'b01101100101: data <= 32'h35653fb4;
    11'b01101100110: data <= 32'h32a8b015;
    11'b01101100111: data <= 32'h37afbe21;
    11'b01101101000: data <= 32'ha535bd1b;
    11'b01101101001: data <= 32'hbbccba01;
    11'b01101101010: data <= 32'hb9adbc6c;
    11'b01101101011: data <= 32'h3bdfbe0c;
    11'b01101101100: data <= 32'h3fbcbada;
    11'b01101101101: data <= 32'h38363454;
    11'b01101101110: data <= 32'hbf2f3901;
    11'b01101101111: data <= 32'hc0e0358a;
    11'b01101110000: data <= 32'hbcdc36e1;
    11'b01101110001: data <= 32'hb40839bd;
    11'b01101110010: data <= 32'hb8ed3088;
    11'b01101110011: data <= 32'hbbc4bc0a;
    11'b01101110100: data <= 32'haa62bb5d;
    11'b01101110101: data <= 32'h3d0d3be5;
    11'b01101110110: data <= 32'h3dbe4157;
    11'b01101110111: data <= 32'h391a4034;
    11'b01101111000: data <= 32'h308d310c;
    11'b01101111001: data <= 32'h311eb9a8;
    11'b01101111010: data <= 32'hadeca7ce;
    11'b01101111011: data <= 32'hb7673453;
    11'b01101111100: data <= 32'h31dfbb13;
    11'b01101111101: data <= 32'h3eefc017;
    11'b01101111110: data <= 32'h408dbe3e;
    11'b01101111111: data <= 32'h39eaacad;
    11'b01110000000: data <= 32'hbcf83915;
    11'b01110000001: data <= 32'hbe033405;
    11'b01110000010: data <= 32'hb715b0c3;
    11'b01110000011: data <= 32'hb42db354;
    11'b01110000100: data <= 32'hbdd5b96b;
    11'b01110000101: data <= 32'hc01fbd68;
    11'b01110000110: data <= 32'hb9f4bb8d;
    11'b01110000111: data <= 32'h3c4c3a90;
    11'b01110001000: data <= 32'h3d484059;
    11'b01110001001: data <= 32'h30dc3ea7;
    11'b01110001010: data <= 32'hb9753620;
    11'b01110001011: data <= 32'hb8583583;
    11'b01110001100: data <= 32'hb47e3d4c;
    11'b01110001101: data <= 32'hb2dd3cc9;
    11'b01110001110: data <= 32'h36d9b91e;
    11'b01110001111: data <= 32'h3ebfc02c;
    11'b01110010000: data <= 32'h4055bd66;
    11'b01110010001: data <= 32'h3c7237ae;
    11'b01110010010: data <= 32'hb09a3c71;
    11'b01110010011: data <= 32'had9132b4;
    11'b01110010100: data <= 32'h3858b986;
    11'b01110010101: data <= 32'hadccbab0;
    11'b01110010110: data <= 32'hbf27bbe1;
    11'b01110010111: data <= 32'hc089bde1;
    11'b01110011000: data <= 32'hb891bd5f;
    11'b01110011001: data <= 32'h3d28b0f0;
    11'b01110011010: data <= 32'h3c553b4c;
    11'b01110011011: data <= 32'hb8e13a75;
    11'b01110011100: data <= 32'hbe2c3652;
    11'b01110011101: data <= 32'hbc393c0c;
    11'b01110011110: data <= 32'hb7493ff6;
    11'b01110011111: data <= 32'hb7b03dbe;
    11'b01110100000: data <= 32'hb459b8fe;
    11'b01110100001: data <= 32'h39e3bf16;
    11'b01110100010: data <= 32'h3e52b848;
    11'b01110100011: data <= 32'h3d7c3db6;
    11'b01110100100: data <= 32'h3aa73eaf;
    11'b01110100101: data <= 32'h3bb4347c;
    11'b01110100110: data <= 32'h3c7eb9ad;
    11'b01110100111: data <= 32'h2c74b834;
    11'b01110101000: data <= 32'hbe30b6ab;
    11'b01110101001: data <= 32'hbe71bcc1;
    11'b01110101010: data <= 32'h343dbf59;
    11'b01110101011: data <= 32'h3f09bd63;
    11'b01110101100: data <= 32'h3ba6b5db;
    11'b01110101101: data <= 32'hbbf22a44;
    11'b01110101110: data <= 32'hbeb53345;
    11'b01110101111: data <= 32'hbaec3bdd;
    11'b01110110000: data <= 32'hb6933ea9;
    11'b01110110001: data <= 32'hbc633b21;
    11'b01110110010: data <= 32'hbe26bb26;
    11'b01110110011: data <= 32'hb8b9bdbc;
    11'b01110110100: data <= 32'h3ab331ab;
    11'b01110110101: data <= 32'h3d6b3fdc;
    11'b01110110110: data <= 32'h3c7f3f2c;
    11'b01110110111: data <= 32'h3c3f3581;
    11'b01110111000: data <= 32'h3bb0b0dd;
    11'b01110111001: data <= 32'h29f638fc;
    11'b01110111010: data <= 32'hbc323a51;
    11'b01110111011: data <= 32'hb9a0b8e0;
    11'b01110111100: data <= 32'h3c3ac02f;
    11'b01110111101: data <= 32'h4022c00d;
    11'b01110111110: data <= 32'h3bf0bb28;
    11'b01110111111: data <= 32'hb965b0a3;
    11'b01111000000: data <= 32'hbaaf2aa0;
    11'b01111000001: data <= 32'h2d1f36d7;
    11'b01111000010: data <= 32'hac2a39ed;
    11'b01111000011: data <= 32'hbe942a99;
    11'b01111000100: data <= 32'hc12ebce2;
    11'b01111000101: data <= 32'hbdf3bd4d;
    11'b01111000110: data <= 32'h366632b5;
    11'b01111000111: data <= 32'h3c7b3e3c;
    11'b01111001000: data <= 32'h394d3ccd;
    11'b01111001001: data <= 32'h34b03355;
    11'b01111001010: data <= 32'h344038d1;
    11'b01111001011: data <= 32'hb06a3fbc;
    11'b01111001100: data <= 32'hb9b03fbb;
    11'b01111001101: data <= 32'hb4b8acba;
    11'b01111001110: data <= 32'h3c66bfe5;
    11'b01111001111: data <= 32'h3f55bf56;
    11'b01111010000: data <= 32'h3c33b6e5;
    11'b01111010001: data <= 32'h30393490;
    11'b01111010010: data <= 32'h383e1c6c;
    11'b01111010011: data <= 32'h3d2bb163;
    11'b01111010100: data <= 32'h36de1e2e;
    11'b01111010101: data <= 32'hbf1eb587;
    11'b01111010110: data <= 32'hc19ebcfc;
    11'b01111010111: data <= 32'hbdbebdc8;
    11'b01111011000: data <= 32'h3835b7c1;
    11'b01111011001: data <= 32'h3ae535a5;
    11'b01111011010: data <= 32'hb0182f61;
    11'b01111011011: data <= 32'hb945aed8;
    11'b01111011100: data <= 32'hb5483c2d;
    11'b01111011101: data <= 32'hb40a4137;
    11'b01111011110: data <= 32'hb9eb40a7;
    11'b01111011111: data <= 32'hb9dc2cfc;
    11'b01111100000: data <= 32'h32d7be75;
    11'b01111100001: data <= 32'h3c1abc07;
    11'b01111100010: data <= 32'h3b973897;
    11'b01111100011: data <= 32'h3ae03b55;
    11'b01111100100: data <= 32'h3e59294b;
    11'b01111100101: data <= 32'h401fb619;
    11'b01111100110: data <= 32'h3a342ce8;
    11'b01111100111: data <= 32'hbddb30c0;
    11'b01111101000: data <= 32'hc04dba1d;
    11'b01111101001: data <= 32'hb8a0be52;
    11'b01111101010: data <= 32'h3c2ebda8;
    11'b01111101011: data <= 32'h39bfbb6e;
    11'b01111101100: data <= 32'hb952bae4;
    11'b01111101101: data <= 32'hbc07b816;
    11'b01111101110: data <= 32'hb32a3b44;
    11'b01111101111: data <= 32'ha8a14095;
    11'b01111110000: data <= 32'hbc0d3f32;
    11'b01111110001: data <= 32'hbee9b2cd;
    11'b01111110010: data <= 32'hbc71bd11;
    11'b01111110011: data <= 32'h294db196;
    11'b01111110100: data <= 32'h39343d32;
    11'b01111110101: data <= 32'h3c0d3c85;
    11'b01111110110: data <= 32'h3ed0a84a;
    11'b01111110111: data <= 32'h3fd5b07c;
    11'b01111111000: data <= 32'h3a283baa;
    11'b01111111001: data <= 32'hbba13d61;
    11'b01111111010: data <= 32'hbc9a2c4a;
    11'b01111111011: data <= 32'h360bbe12;
    11'b01111111100: data <= 32'h3dcfbfb2;
    11'b01111111101: data <= 32'h3931bdef;
    11'b01111111110: data <= 32'hb90dbca5;
    11'b01111111111: data <= 32'hb6d5ba03;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    