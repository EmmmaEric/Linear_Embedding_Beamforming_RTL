
module memory_rom_62(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbcfdbbb4;
    11'b00000000001: data <= 32'hba6cb82b;
    11'b00000000010: data <= 32'h39693845;
    11'b00000000011: data <= 32'h3aee3e9f;
    11'b00000000100: data <= 32'hba9d3e06;
    11'b00000000101: data <= 32'hc0a5338a;
    11'b00000000110: data <= 32'hbf78b5d5;
    11'b00000000111: data <= 32'hb4723755;
    11'b00000001000: data <= 32'h39923c9c;
    11'b00000001001: data <= 32'h3b2c3525;
    11'b00000001010: data <= 32'h3cf2baf8;
    11'b00000001011: data <= 32'h3e7eb5bc;
    11'b00000001100: data <= 32'h3c883e06;
    11'b00000001101: data <= 32'h9c144060;
    11'b00000001110: data <= 32'hb623388c;
    11'b00000001111: data <= 32'h34f9be1c;
    11'b00000010000: data <= 32'h392ec013;
    11'b00000010001: data <= 32'hb202bd3b;
    11'b00000010010: data <= 32'hbab9bb2d;
    11'b00000010011: data <= 32'h2eadbbd4;
    11'b00000010100: data <= 32'h3e22b85b;
    11'b00000010101: data <= 32'h3c773695;
    11'b00000010110: data <= 32'hbcc339d9;
    11'b00000010111: data <= 32'hc1a83104;
    11'b00000011000: data <= 32'hc049b06e;
    11'b00000011001: data <= 32'hb77f362c;
    11'b00000011010: data <= 32'h30c138c9;
    11'b00000011011: data <= 32'hb1b3b472;
    11'b00000011100: data <= 32'h2647bb59;
    11'b00000011101: data <= 32'h3b403470;
    11'b00000011110: data <= 32'h3cc640c2;
    11'b00000011111: data <= 32'h38004197;
    11'b00000100000: data <= 32'hab233b27;
    11'b00000100001: data <= 32'h3159bc45;
    11'b00000100010: data <= 32'h3580bca7;
    11'b00000100011: data <= 32'hac83b4c5;
    11'b00000100100: data <= 32'hac53b5fc;
    11'b00000100101: data <= 32'h3cadbd23;
    11'b00000100110: data <= 32'h40a3bd8a;
    11'b00000100111: data <= 32'h3dc7b4fb;
    11'b00000101000: data <= 32'hbbc6381f;
    11'b00000101001: data <= 32'hc0a93389;
    11'b00000101010: data <= 32'hbdedb51e;
    11'b00000101011: data <= 32'hb29ab5c6;
    11'b00000101100: data <= 32'hb66bb722;
    11'b00000101101: data <= 32'hbd44bc32;
    11'b00000101110: data <= 32'hbc15bc7e;
    11'b00000101111: data <= 32'h3738362c;
    11'b00000110000: data <= 32'h3ccc40b4;
    11'b00000110001: data <= 32'h369a411f;
    11'b00000110010: data <= 32'hb8e93b2d;
    11'b00000110011: data <= 32'hb970b5dc;
    11'b00000110100: data <= 32'hb3f6302b;
    11'b00000110101: data <= 32'hab3e3b66;
    11'b00000110110: data <= 32'h361731a6;
    11'b00000110111: data <= 32'h3e57bd85;
    11'b00000111000: data <= 32'h40f9be40;
    11'b00000111001: data <= 32'h3ea0ad93;
    11'b00000111010: data <= 32'hb4203c3c;
    11'b00000111011: data <= 32'hbc5c38a0;
    11'b00000111100: data <= 32'hb480b89c;
    11'b00000111101: data <= 32'h34afbc64;
    11'b00000111110: data <= 32'hb99fbcc2;
    11'b00000111111: data <= 32'hbf80bdf0;
    11'b00001000000: data <= 32'hbce9bdae;
    11'b00001000001: data <= 32'h393db234;
    11'b00001000010: data <= 32'h3d4d3d6e;
    11'b00001000011: data <= 32'h9cdd3e57;
    11'b00001000100: data <= 32'hbe1738a8;
    11'b00001000101: data <= 32'hbe6031f0;
    11'b00001000110: data <= 32'hba2f3c4d;
    11'b00001000111: data <= 32'hb4583e44;
    11'b00001001000: data <= 32'h2c9c348f;
    11'b00001001001: data <= 32'h3bc3bd93;
    11'b00001001010: data <= 32'h3f77bc9b;
    11'b00001001011: data <= 32'h3e6c3a80;
    11'b00001001100: data <= 32'h38333fe8;
    11'b00001001101: data <= 32'h30983c20;
    11'b00001001110: data <= 32'h397cb8b4;
    11'b00001001111: data <= 32'h38ecbcaa;
    11'b00001010000: data <= 32'hb9d7bc08;
    11'b00001010001: data <= 32'hbea1bcf5;
    11'b00001010010: data <= 32'hb85abe7c;
    11'b00001010011: data <= 32'h3da9bc85;
    11'b00001010100: data <= 32'h3e749f01;
    11'b00001010101: data <= 32'hb4d637be;
    11'b00001010110: data <= 32'hc0003293;
    11'b00001010111: data <= 32'hbf5435a8;
    11'b00001011000: data <= 32'hbaa03cc3;
    11'b00001011001: data <= 32'hb8dc3d0d;
    11'b00001011010: data <= 32'hbafeb22e;
    11'b00001011011: data <= 32'hb59dbdf0;
    11'b00001011100: data <= 32'h3aa0b8f1;
    11'b00001011101: data <= 32'h3d673e80;
    11'b00001011110: data <= 32'h3b90411a;
    11'b00001011111: data <= 32'h39413d10;
    11'b00001100000: data <= 32'h3a8fb49a;
    11'b00001100001: data <= 32'h376fb65c;
    11'b00001100010: data <= 32'hb9392e4f;
    11'b00001100011: data <= 32'hbc10b697;
    11'b00001100100: data <= 32'h36e0be6b;
    11'b00001100101: data <= 32'h4057bf77;
    11'b00001100110: data <= 32'h3f91bb48;
    11'b00001100111: data <= 32'hb220a89d;
    11'b00001101000: data <= 32'hbe572df9;
    11'b00001101001: data <= 32'hbc57325e;
    11'b00001101010: data <= 32'hb49b38c7;
    11'b00001101011: data <= 32'hbac43574;
    11'b00001101100: data <= 32'hbf98bb71;
    11'b00001101101: data <= 32'hbe48beb6;
    11'b00001101110: data <= 32'h29e8b73a;
    11'b00001101111: data <= 32'h3c813e9e;
    11'b00001110000: data <= 32'h3ae8407e;
    11'b00001110001: data <= 32'h344b3c1a;
    11'b00001110010: data <= 32'h30242ff1;
    11'b00001110011: data <= 32'had4e3a3e;
    11'b00001110100: data <= 32'hb9403df6;
    11'b00001110101: data <= 32'hb87337b0;
    11'b00001110110: data <= 32'h3b07bdbf;
    11'b00001110111: data <= 32'h4092c00d;
    11'b00001111000: data <= 32'h3f9cbaf0;
    11'b00001111001: data <= 32'h343b3508;
    11'b00001111010: data <= 32'hb74435e3;
    11'b00001111011: data <= 32'h346fa5b7;
    11'b00001111100: data <= 32'h3879aef0;
    11'b00001111101: data <= 32'hbadcb694;
    11'b00001111110: data <= 32'hc0d5bd57;
    11'b00001111111: data <= 32'hbfdfbf48;
    11'b00010000000: data <= 32'h24f3ba7f;
    11'b00010000001: data <= 32'h3c9b3a1c;
    11'b00010000010: data <= 32'h37c53c7a;
    11'b00010000011: data <= 32'hb89535db;
    11'b00010000100: data <= 32'hba2035f0;
    11'b00010000101: data <= 32'hb8b83ead;
    11'b00010000110: data <= 32'hba2240a9;
    11'b00010000111: data <= 32'hb9843ad9;
    11'b00010001000: data <= 32'h35b9bd3f;
    11'b00010001001: data <= 32'h3e20be97;
    11'b00010001010: data <= 32'h3e18ac23;
    11'b00010001011: data <= 32'h39e83cba;
    11'b00010001100: data <= 32'h39b33a7b;
    11'b00010001101: data <= 32'h3dceae0a;
    11'b00010001110: data <= 32'h3cbcb4e3;
    11'b00010001111: data <= 32'hb9abb503;
    11'b00010010000: data <= 32'hc071bbda;
    11'b00010010001: data <= 32'hbda0bee3;
    11'b00010010010: data <= 32'h3992bdc9;
    11'b00010010011: data <= 32'h3db1b837;
    11'b00010010100: data <= 32'h3130b23b;
    11'b00010010101: data <= 32'hbc8bb57f;
    11'b00010010110: data <= 32'hbc4c3537;
    11'b00010010111: data <= 32'hb8853f30;
    11'b00010011000: data <= 32'hbabf4059;
    11'b00010011001: data <= 32'hbd6937fa;
    11'b00010011010: data <= 32'hbb12bd7e;
    11'b00010011011: data <= 32'h3487bc73;
    11'b00010011100: data <= 32'h3b4d3a5d;
    11'b00010011101: data <= 32'h3b4d3f3f;
    11'b00010011110: data <= 32'h3ce83bed;
    11'b00010011111: data <= 32'h3f09a006;
    11'b00010100000: data <= 32'h3cca32ac;
    11'b00010100001: data <= 32'hb8a039b2;
    11'b00010100010: data <= 32'hbe5f29ec;
    11'b00010100011: data <= 32'hb6babd5e;
    11'b00010100100: data <= 32'h3df6bfa4;
    11'b00010100101: data <= 32'h3eafbdad;
    11'b00010100110: data <= 32'h2ebdbb4e;
    11'b00010100111: data <= 32'hbb8ab958;
    11'b00010101000: data <= 32'hb68d2d8b;
    11'b00010101001: data <= 32'h31023ce6;
    11'b00010101010: data <= 32'hb9cd3d19;
    11'b00010101011: data <= 32'hc02fb41e;
    11'b00010101100: data <= 32'hc02abe35;
    11'b00010101101: data <= 32'hb9bfba91;
    11'b00010101110: data <= 32'h36d93c0d;
    11'b00010101111: data <= 32'h39aa3e5c;
    11'b00010110000: data <= 32'h3ae838c1;
    11'b00010110001: data <= 32'h3c812c55;
    11'b00010110010: data <= 32'h39483c66;
    11'b00010110011: data <= 32'hb89c4027;
    11'b00010110100: data <= 32'hbc2f3cb0;
    11'b00010110101: data <= 32'h31f1bafb;
    11'b00010110110: data <= 32'h3ec3bfa2;
    11'b00010110111: data <= 32'h3e38bd9a;
    11'b00010111000: data <= 32'h3410b944;
    11'b00010111001: data <= 32'hadbfb715;
    11'b00010111010: data <= 32'h3b5db095;
    11'b00010111011: data <= 32'h3cfb376d;
    11'b00010111100: data <= 32'hb6793659;
    11'b00010111101: data <= 32'hc0d4b9fb;
    11'b00010111110: data <= 32'hc101be68;
    11'b00010111111: data <= 32'hbb06bb46;
    11'b00011000000: data <= 32'h35b83634;
    11'b00011000001: data <= 32'h34e43805;
    11'b00011000010: data <= 32'ha02cb4e6;
    11'b00011000011: data <= 32'h3077a8c0;
    11'b00011000100: data <= 32'h2c863f13;
    11'b00011000101: data <= 32'hb90341e0;
    11'b00011000110: data <= 32'hbb953ede;
    11'b00011000111: data <= 32'had6fb8cd;
    11'b00011001000: data <= 32'h3be4bded;
    11'b00011001001: data <= 32'h3b92b8af;
    11'b00011001010: data <= 32'h35e6343b;
    11'b00011001011: data <= 32'h3ab72c64;
    11'b00011001100: data <= 32'h403bb3fa;
    11'b00011001101: data <= 32'h40252cde;
    11'b00011001110: data <= 32'hab5a3434;
    11'b00011001111: data <= 32'hc048b753;
    11'b00011010000: data <= 32'hbfc3bd2f;
    11'b00011010001: data <= 32'hb1e4bcc1;
    11'b00011010010: data <= 32'h3964b93b;
    11'b00011010011: data <= 32'ha8a3baaa;
    11'b00011010100: data <= 32'hb9ccbcff;
    11'b00011010101: data <= 32'hb614b540;
    11'b00011010110: data <= 32'h24553f25;
    11'b00011010111: data <= 32'hb83a4195;
    11'b00011011000: data <= 32'hbd183d89;
    11'b00011011001: data <= 32'hbc4ab963;
    11'b00011011010: data <= 32'hb478bb73;
    11'b00011011011: data <= 32'h2d213655;
    11'b00011011100: data <= 32'h34143c54;
    11'b00011011101: data <= 32'h3cdc356f;
    11'b00011011110: data <= 32'h40e5b4d3;
    11'b00011011111: data <= 32'h40503476;
    11'b00011100000: data <= 32'h2e7e3c21;
    11'b00011100001: data <= 32'hbdf7389b;
    11'b00011100010: data <= 32'hbadfb937;
    11'b00011100011: data <= 32'h3a2dbd55;
    11'b00011100100: data <= 32'h3c13bd89;
    11'b00011100101: data <= 32'hb257be5b;
    11'b00011100110: data <= 32'hba7cbec6;
    11'b00011100111: data <= 32'h2842b927;
    11'b00011101000: data <= 32'h39d63cbb;
    11'b00011101001: data <= 32'hb0d23f49;
    11'b00011101010: data <= 32'hbeb137e9;
    11'b00011101011: data <= 32'hc02cbb95;
    11'b00011101100: data <= 32'hbd51b880;
    11'b00011101101: data <= 32'hb8953ae7;
    11'b00011101110: data <= 32'had163c6d;
    11'b00011101111: data <= 32'h3a6ca76b;
    11'b00011110000: data <= 32'h3f13b780;
    11'b00011110001: data <= 32'h3e163a9c;
    11'b00011110010: data <= 32'h24cf4065;
    11'b00011110011: data <= 32'hbb1e3f07;
    11'b00011110100: data <= 32'ha80a2724;
    11'b00011110101: data <= 32'h3cdabc98;
    11'b00011110110: data <= 32'h3b9cbd2d;
    11'b00011110111: data <= 32'hb449bd42;
    11'b00011111000: data <= 32'hb4c2bda9;
    11'b00011111001: data <= 32'h3c9cba7e;
    11'b00011111010: data <= 32'h3f7f3618;
    11'b00011111011: data <= 32'h369539fe;
    11'b00011111100: data <= 32'hbf11b359;
    11'b00011111101: data <= 32'hc0d3bc46;
    11'b00011111110: data <= 32'hbdfab764;
    11'b00011111111: data <= 32'hb9253887;
    11'b00100000000: data <= 32'hb7473398;
    11'b00100000001: data <= 32'hae9cbbd8;
    11'b00100000010: data <= 32'h38efbaad;
    11'b00100000011: data <= 32'h39af3ceb;
    11'b00100000100: data <= 32'hafcb41e4;
    11'b00100000101: data <= 32'hb91140a9;
    11'b00100000110: data <= 32'h222635af;
    11'b00100000111: data <= 32'h39e6b9a0;
    11'b00100001000: data <= 32'h34dbb710;
    11'b00100001001: data <= 32'hb6c1b417;
    11'b00100001010: data <= 32'h3574b9a3;
    11'b00100001011: data <= 32'h4071ba88;
    11'b00100001100: data <= 32'h4182b04a;
    11'b00100001101: data <= 32'h3af13516;
    11'b00100001110: data <= 32'hbdb4b1c2;
    11'b00100001111: data <= 32'hbf39b9f6;
    11'b00100010000: data <= 32'hb98eb79c;
    11'b00100010001: data <= 32'hb11db157;
    11'b00100010010: data <= 32'hb993bbab;
    11'b00100010011: data <= 32'hbb5ebffb;
    11'b00100010100: data <= 32'hb1c4bd23;
    11'b00100010101: data <= 32'h36813c88;
    11'b00100010110: data <= 32'ha860417d;
    11'b00100010111: data <= 32'hb9a93fb2;
    11'b00100011000: data <= 32'hb93f3104;
    11'b00100011001: data <= 32'hb5fdb39e;
    11'b00100011010: data <= 32'hb92d38fc;
    11'b00100011011: data <= 32'hb9e93a8b;
    11'b00100011100: data <= 32'h387ab1b5;
    11'b00100011101: data <= 32'h40fbbaa1;
    11'b00100011110: data <= 32'h4198b117;
    11'b00100011111: data <= 32'h3b9a3a1e;
    11'b00100100000: data <= 32'hbab33976;
    11'b00100100001: data <= 32'hb935a391;
    11'b00100100010: data <= 32'h37efb623;
    11'b00100100011: data <= 32'h3701b999;
    11'b00100100100: data <= 32'hba5bbe95;
    11'b00100100101: data <= 32'hbcd5c0e0;
    11'b00100100110: data <= 32'hadb2be51;
    11'b00100100111: data <= 32'h3b6c3875;
    11'b00100101000: data <= 32'h36b73ed4;
    11'b00100101001: data <= 32'hbacf3a98;
    11'b00100101010: data <= 32'hbdc3b5c5;
    11'b00100101011: data <= 32'hbd642a56;
    11'b00100101100: data <= 32'hbd583d12;
    11'b00100101101: data <= 32'hbc723ca4;
    11'b00100101110: data <= 32'h3061b55e;
    11'b00100101111: data <= 32'h3f00bc35;
    11'b00100110000: data <= 32'h3fef3003;
    11'b00100110001: data <= 32'h39273eb1;
    11'b00100110010: data <= 32'hb52e3f1b;
    11'b00100110011: data <= 32'h355839dc;
    11'b00100110100: data <= 32'h3cffae96;
    11'b00100110101: data <= 32'h38d0b879;
    11'b00100110110: data <= 32'hbb29bd42;
    11'b00100110111: data <= 32'hbba1c009;
    11'b00100111000: data <= 32'h3a0cbe39;
    11'b00100111001: data <= 32'h3fe3b109;
    11'b00100111010: data <= 32'h3c4837eb;
    11'b00100111011: data <= 32'hba63b29d;
    11'b00100111100: data <= 32'hbeb2b9d8;
    11'b00100111101: data <= 32'hbdd830f0;
    11'b00100111110: data <= 32'hbd3e3ce1;
    11'b00100111111: data <= 32'hbd5c38a4;
    11'b00101000000: data <= 32'hb98ebcae;
    11'b00101000001: data <= 32'h3790be11;
    11'b00101000010: data <= 32'h3b03357b;
    11'b00101000011: data <= 32'h33b14096;
    11'b00101000100: data <= 32'hadc4409a;
    11'b00101000101: data <= 32'h38ea3c0b;
    11'b00101000110: data <= 32'h3c4f3401;
    11'b00101000111: data <= 32'h2de833b0;
    11'b00101001000: data <= 32'hbc98b0a7;
    11'b00101001001: data <= 32'hb83dbc21;
    11'b00101001010: data <= 32'h3ea9bd2c;
    11'b00101001011: data <= 32'h419cb902;
    11'b00101001100: data <= 32'h3e16b11c;
    11'b00101001101: data <= 32'hb7dfb797;
    11'b00101001110: data <= 32'hbc5db895;
    11'b00101001111: data <= 32'hb883335b;
    11'b00101010000: data <= 32'hb8a539c3;
    11'b00101010001: data <= 32'hbd4db6e1;
    11'b00101010010: data <= 32'hbdcdc047;
    11'b00101010011: data <= 32'hb843c001;
    11'b00101010100: data <= 32'h33c93338;
    11'b00101010101: data <= 32'h3034402c;
    11'b00101010110: data <= 32'hae093f3f;
    11'b00101010111: data <= 32'h322538d3;
    11'b00101011000: data <= 32'h31aa37b8;
    11'b00101011001: data <= 32'hba763cf4;
    11'b00101011010: data <= 32'hbe233c7d;
    11'b00101011011: data <= 32'hb621b176;
    11'b00101011100: data <= 32'h3f98bc51;
    11'b00101011101: data <= 32'h4190b992;
    11'b00101011110: data <= 32'h3dc228ab;
    11'b00101011111: data <= 32'hae6d30c9;
    11'b00101100000: data <= 32'h14952e05;
    11'b00101100001: data <= 32'h3a7536a3;
    11'b00101100010: data <= 32'h359e34de;
    11'b00101100011: data <= 32'hbcb1bc39;
    11'b00101100100: data <= 32'hbf06c110;
    11'b00101100101: data <= 32'hb989c05d;
    11'b00101100110: data <= 32'h37fbb248;
    11'b00101100111: data <= 32'h37fa3c65;
    11'b00101101000: data <= 32'hb049385a;
    11'b00101101001: data <= 32'hb700b3a4;
    11'b00101101010: data <= 32'hb9ab3811;
    11'b00101101011: data <= 32'hbddb3f85;
    11'b00101101100: data <= 32'hbf5f3ed9;
    11'b00101101101: data <= 32'hb999a89f;
    11'b00101101110: data <= 32'h3cc8bcbe;
    11'b00101101111: data <= 32'h3f44b81b;
    11'b00101110000: data <= 32'h3a9f3a14;
    11'b00101110001: data <= 32'h30cd3c83;
    11'b00101110010: data <= 32'h3bc03a8f;
    11'b00101110011: data <= 32'h3f393975;
    11'b00101110100: data <= 32'h3aa43640;
    11'b00101110101: data <= 32'hbc7eb9f9;
    11'b00101110110: data <= 32'hbe5dbff1;
    11'b00101110111: data <= 32'haadbbf87;
    11'b00101111000: data <= 32'h3d98b943;
    11'b00101111001: data <= 32'h3c85ad9b;
    11'b00101111010: data <= 32'haa99b9d7;
    11'b00101111011: data <= 32'hb965bb8f;
    11'b00101111100: data <= 32'hba9f36e1;
    11'b00101111101: data <= 32'hbd5b3f9f;
    11'b00101111110: data <= 32'hbf5b3d6b;
    11'b00101111111: data <= 32'hbd32b992;
    11'b00110000000: data <= 32'haa8dbe7d;
    11'b00110000001: data <= 32'h378fb5b3;
    11'b00110000010: data <= 32'h2ca43d5a;
    11'b00110000011: data <= 32'h317a3e90;
    11'b00110000100: data <= 32'h3d3b3c1c;
    11'b00110000101: data <= 32'h3f7c3ad4;
    11'b00110000110: data <= 32'h38383bee;
    11'b00110000111: data <= 32'hbd553643;
    11'b00110001000: data <= 32'hbcfdba30;
    11'b00110001001: data <= 32'h3a32bd0d;
    11'b00110001010: data <= 32'h4066bb20;
    11'b00110001011: data <= 32'h3e25ba49;
    11'b00110001100: data <= 32'h300cbd00;
    11'b00110001101: data <= 32'hb400bc1e;
    11'b00110001110: data <= 32'h29323700;
    11'b00110001111: data <= 32'hb6773dfc;
    11'b00110010000: data <= 32'hbde83755;
    11'b00110010001: data <= 32'hbf39be75;
    11'b00110010010: data <= 32'hbc58c02b;
    11'b00110010011: data <= 32'hb6d6b655;
    11'b00110010100: data <= 32'hb5143cfc;
    11'b00110010101: data <= 32'h2c533cb2;
    11'b00110010110: data <= 32'h3bd3370f;
    11'b00110010111: data <= 32'h3c763a19;
    11'b00110011000: data <= 32'hb4ca3ef5;
    11'b00110011001: data <= 32'hbed53eb6;
    11'b00110011010: data <= 32'hbc4535cf;
    11'b00110011011: data <= 32'h3c55b9dc;
    11'b00110011100: data <= 32'h4064ba9b;
    11'b00110011101: data <= 32'h3d39b96f;
    11'b00110011110: data <= 32'h335bba6a;
    11'b00110011111: data <= 32'h38d7b775;
    11'b00110100000: data <= 32'h3db238ee;
    11'b00110100001: data <= 32'h3a6f3c57;
    11'b00110100010: data <= 32'hbbdab28e;
    11'b00110100011: data <= 32'hbfc6c00c;
    11'b00110100100: data <= 32'hbd50c04c;
    11'b00110100101: data <= 32'hb608b893;
    11'b00110100110: data <= 32'hadde379b;
    11'b00110100111: data <= 32'h2384ae74;
    11'b00110101000: data <= 32'h3628b961;
    11'b00110101001: data <= 32'h335536e1;
    11'b00110101010: data <= 32'hbbbe405f;
    11'b00110101011: data <= 32'hbfc140af;
    11'b00110101100: data <= 32'hbcbe39d8;
    11'b00110101101: data <= 32'h3893b93b;
    11'b00110101110: data <= 32'h3ce9b8e1;
    11'b00110101111: data <= 32'h36f4a338;
    11'b00110110000: data <= 32'h2fa93083;
    11'b00110110001: data <= 32'h3d713434;
    11'b00110110010: data <= 32'h40fc3ab5;
    11'b00110110011: data <= 32'h3e2b3c17;
    11'b00110110100: data <= 32'hb99dabbb;
    11'b00110110101: data <= 32'hbedfbded;
    11'b00110110110: data <= 32'hba17be73;
    11'b00110110111: data <= 32'h3733b975;
    11'b00110111000: data <= 32'h3831b7de;
    11'b00110111001: data <= 32'h2cdcbdc4;
    11'b00110111010: data <= 32'h29e6bea3;
    11'b00110111011: data <= 32'ha6732d25;
    11'b00110111100: data <= 32'hbadd403e;
    11'b00110111101: data <= 32'hbeeb4021;
    11'b00110111110: data <= 32'hbdd231c2;
    11'b00110111111: data <= 32'hb748bc31;
    11'b00111000000: data <= 32'hb1c1b71c;
    11'b00111000001: data <= 32'hb8f338fc;
    11'b00111000010: data <= 32'hb1583a11;
    11'b00111000011: data <= 32'h3e5337ec;
    11'b00111000100: data <= 32'h41493ac3;
    11'b00111000101: data <= 32'h3d8b3d4e;
    11'b00111000110: data <= 32'hbaab3ae9;
    11'b00111000111: data <= 32'hbd75b2d6;
    11'b00111001000: data <= 32'h2df5b97f;
    11'b00111001001: data <= 32'h3d4db8a1;
    11'b00111001010: data <= 32'h3bb1bc30;
    11'b00111001011: data <= 32'h302bc01c;
    11'b00111001100: data <= 32'h32debfba;
    11'b00111001101: data <= 32'h391fa7ee;
    11'b00111001110: data <= 32'h2fc43ec7;
    11'b00111001111: data <= 32'hbc443cac;
    11'b00111010000: data <= 32'hbe6fba3e;
    11'b00111010001: data <= 32'hbd4fbe29;
    11'b00111010010: data <= 32'hbcb9b657;
    11'b00111010011: data <= 32'hbcf339f5;
    11'b00111010100: data <= 32'hb6f837a9;
    11'b00111010101: data <= 32'h3ce0afae;
    11'b00111010110: data <= 32'h3fa6378e;
    11'b00111010111: data <= 32'h38683ee0;
    11'b00111011000: data <= 32'hbced3fe4;
    11'b00111011001: data <= 32'hbc823c1d;
    11'b00111011010: data <= 32'h38982f0b;
    11'b00111011011: data <= 32'h3df7b4ce;
    11'b00111011100: data <= 32'h39c0bb1c;
    11'b00111011101: data <= 32'ha4fabe9d;
    11'b00111011110: data <= 32'h39cfbd98;
    11'b00111011111: data <= 32'h3f5b30f7;
    11'b00111100000: data <= 32'h3dbe3cfd;
    11'b00111100001: data <= 32'hb46735e7;
    11'b00111100010: data <= 32'hbdf3bd5f;
    11'b00111100011: data <= 32'hbdfbbe72;
    11'b00111100100: data <= 32'hbcccb5aa;
    11'b00111100101: data <= 32'hbc5a34be;
    11'b00111100110: data <= 32'hb813b8e1;
    11'b00111100111: data <= 32'h38d1bd57;
    11'b00111101000: data <= 32'h3b63b190;
    11'b00111101001: data <= 32'hb4133f7c;
    11'b00111101010: data <= 32'hbdf34115;
    11'b00111101011: data <= 32'hbc423df1;
    11'b00111101100: data <= 32'h35c13510;
    11'b00111101101: data <= 32'h39aba659;
    11'b00111101110: data <= 32'hb3ceb278;
    11'b00111101111: data <= 32'hb72db923;
    11'b00111110000: data <= 32'h3ca8b872;
    11'b00111110001: data <= 32'h419736a9;
    11'b00111110010: data <= 32'h408f3c2a;
    11'b00111110011: data <= 32'h31d533da;
    11'b00111110100: data <= 32'hbca0bbe6;
    11'b00111110101: data <= 32'hbb35bbff;
    11'b00111110110: data <= 32'hb55eb0dc;
    11'b00111110111: data <= 32'hb63cb573;
    11'b00111111000: data <= 32'hb679bf4e;
    11'b00111111001: data <= 32'h30fdc0e4;
    11'b00111111010: data <= 32'h36e6b9fc;
    11'b00111111011: data <= 32'hb54c3e9e;
    11'b00111111100: data <= 32'hbce84073;
    11'b00111111101: data <= 32'hbc283b6e;
    11'b00111111110: data <= 32'hb55aafc6;
    11'b00111111111: data <= 32'hb8882eca;
    11'b01000000000: data <= 32'hbdbc381e;
    11'b01000000001: data <= 32'hbc0031ca;
    11'b01000000010: data <= 32'h3cc1b06f;
    11'b01000000011: data <= 32'h41cb3662;
    11'b01000000100: data <= 32'h404c3c50;
    11'b01000000101: data <= 32'h2ac93aba;
    11'b01000000110: data <= 32'hba893070;
    11'b01000000111: data <= 32'h23d22c4c;
    11'b01000001000: data <= 32'h39b733f2;
    11'b01000001001: data <= 32'h3336b94d;
    11'b01000001010: data <= 32'hb58dc0c4;
    11'b01000001011: data <= 32'h2de7c18d;
    11'b01000001100: data <= 32'h3a3dbb4e;
    11'b01000001101: data <= 32'h37eb3cd7;
    11'b01000001110: data <= 32'hb6d73d1c;
    11'b01000001111: data <= 32'hbb01b1a1;
    11'b01000010000: data <= 32'hbb8aba37;
    11'b01000010001: data <= 32'hbe02302b;
    11'b01000010010: data <= 32'hc0493aa9;
    11'b01000010011: data <= 32'hbd823272;
    11'b01000010100: data <= 32'h3a32b8b5;
    11'b01000010101: data <= 32'h403cadf8;
    11'b01000010110: data <= 32'h3cce3c98;
    11'b01000010111: data <= 32'hb7d13ea6;
    11'b01000011000: data <= 32'hb8ea3d3b;
    11'b01000011001: data <= 32'h394b3be8;
    11'b01000011010: data <= 32'h3ca53988;
    11'b01000011011: data <= 32'h3118b69a;
    11'b01000011100: data <= 32'hb8babfc1;
    11'b01000011101: data <= 32'h34a5c055;
    11'b01000011110: data <= 32'h3eb5b8e9;
    11'b01000011111: data <= 32'h3ee83a67;
    11'b01000100000: data <= 32'h3816356b;
    11'b01000100001: data <= 32'hb84dbc02;
    11'b01000100010: data <= 32'hbbd2bc23;
    11'b01000100011: data <= 32'hbded33a4;
    11'b01000100100: data <= 32'hbfd7396f;
    11'b01000100101: data <= 32'hbd84b8a6;
    11'b01000100110: data <= 32'h31f8bed7;
    11'b01000100111: data <= 32'h3c0cbb31;
    11'b01000101000: data <= 32'h30e13c2c;
    11'b01000101001: data <= 32'hbb7f401f;
    11'b01000101010: data <= 32'hb81c3eea;
    11'b01000101011: data <= 32'h39c13cd2;
    11'b01000101100: data <= 32'h397d3b92;
    11'b01000101101: data <= 32'hb9933432;
    11'b01000101110: data <= 32'hbcbabaa0;
    11'b01000101111: data <= 32'h3714bc69;
    11'b01000110000: data <= 32'h40dcb10c;
    11'b01000110001: data <= 32'h411238aa;
    11'b01000110010: data <= 32'h3c18a847;
    11'b01000110011: data <= 32'hb16bbb9f;
    11'b01000110100: data <= 32'hb5e0b85e;
    11'b01000110101: data <= 32'hb84938c2;
    11'b01000110110: data <= 32'hbc4b3580;
    11'b01000110111: data <= 32'hbc59be48;
    11'b01000111000: data <= 32'hb400c192;
    11'b01000111001: data <= 32'h34babe47;
    11'b01000111010: data <= 32'hb36039d8;
    11'b01000111011: data <= 32'hba913ec8;
    11'b01000111100: data <= 32'hb5a23c69;
    11'b01000111101: data <= 32'h355238f1;
    11'b01000111110: data <= 32'hb57f3b4f;
    11'b01000111111: data <= 32'hbf673baa;
    11'b01001000000: data <= 32'hbf74323d;
    11'b01001000001: data <= 32'h351ab620;
    11'b01001000010: data <= 32'h40e79edc;
    11'b01001000011: data <= 32'h40b33812;
    11'b01001000100: data <= 32'h3a52341b;
    11'b01001000101: data <= 32'h2956adaa;
    11'b01001000110: data <= 32'h383737aa;
    11'b01001000111: data <= 32'h39883c9b;
    11'b01001001000: data <= 32'hb14332ea;
    11'b01001001001: data <= 32'hbabbc009;
    11'b01001001010: data <= 32'hb651c226;
    11'b01001001011: data <= 32'h3590beb6;
    11'b01001001100: data <= 32'h351435ee;
    11'b01001001101: data <= 32'hacf33a13;
    11'b01001001110: data <= 32'ha449b119;
    11'b01001001111: data <= 32'ha986b50b;
    11'b01001010000: data <= 32'hbc9339e6;
    11'b01001010001: data <= 32'hc1123d50;
    11'b01001010010: data <= 32'hc07937f8;
    11'b01001010011: data <= 32'habefb851;
    11'b01001010100: data <= 32'h3eacb6bc;
    11'b01001010101: data <= 32'h3d0d3680;
    11'b01001010110: data <= 32'h9ded3a8a;
    11'b01001010111: data <= 32'h29993b5f;
    11'b01001011000: data <= 32'h3cd13d8f;
    11'b01001011001: data <= 32'h3da03e91;
    11'b01001011010: data <= 32'h2cc037c7;
    11'b01001011011: data <= 32'hbbd7be34;
    11'b01001011100: data <= 32'hb5bdc0b1;
    11'b01001011101: data <= 32'h3bbabca0;
    11'b01001011110: data <= 32'h3d7730cd;
    11'b01001011111: data <= 32'h3adeb24c;
    11'b01001100000: data <= 32'h36a5bcf4;
    11'b01001100001: data <= 32'h9ca5bb18;
    11'b01001100010: data <= 32'hbc5539b3;
    11'b01001100011: data <= 32'hc0853d45;
    11'b01001100100: data <= 32'hc01d1c29;
    11'b01001100101: data <= 32'hb7b7bdd2;
    11'b01001100110: data <= 32'h3869bce4;
    11'b01001100111: data <= 32'ha6bd316a;
    11'b01001101000: data <= 32'hba303c5e;
    11'b01001101001: data <= 32'ha38d3d20;
    11'b01001101010: data <= 32'h3d883e2d;
    11'b01001101011: data <= 32'h3ce43f12;
    11'b01001101100: data <= 32'hb86d3c1b;
    11'b01001101101: data <= 32'hbe39b6e6;
    11'b01001101110: data <= 32'hb5c7bc3e;
    11'b01001101111: data <= 32'h3e36b619;
    11'b01001110000: data <= 32'h40302f36;
    11'b01001110001: data <= 32'h3d58b959;
    11'b01001110010: data <= 32'h39b2bdef;
    11'b01001110011: data <= 32'h381bb934;
    11'b01001110100: data <= 32'hb0033c24;
    11'b01001110101: data <= 32'hbcb03c97;
    11'b01001110110: data <= 32'hbdd5ba4d;
    11'b01001110111: data <= 32'hb9cdc0dd;
    11'b01001111000: data <= 32'hb3dabf86;
    11'b01001111001: data <= 32'hb9a4b017;
    11'b01001111010: data <= 32'hbb7c3a2a;
    11'b01001111011: data <= 32'h2dbf391b;
    11'b01001111100: data <= 32'h3ca73a42;
    11'b01001111101: data <= 32'h36ab3dcf;
    11'b01001111110: data <= 32'hbe5b3e1b;
    11'b01001111111: data <= 32'hc07d393f;
    11'b01010000000: data <= 32'hb829a9be;
    11'b01010000001: data <= 32'h3e472cb0;
    11'b01010000010: data <= 32'h3f883005;
    11'b01010000011: data <= 32'h3baeb853;
    11'b01010000100: data <= 32'h396fbaec;
    11'b01010000101: data <= 32'h3ce63387;
    11'b01010000110: data <= 32'h3c9e3e6f;
    11'b01010000111: data <= 32'h26de3c65;
    11'b01010001000: data <= 32'hbb1abcbf;
    11'b01010001001: data <= 32'hba02c15f;
    11'b01010001010: data <= 32'hb582bf87;
    11'b01010001011: data <= 32'hb6c7b4a9;
    11'b01010001100: data <= 32'hb5bc9ef8;
    11'b01010001101: data <= 32'h3710b95c;
    11'b01010001110: data <= 32'h3b34b6e0;
    11'b01010001111: data <= 32'hb4c23b88;
    11'b01010010000: data <= 32'hc0783f00;
    11'b01010010001: data <= 32'hc1173c62;
    11'b01010010010: data <= 32'hba0e2d4a;
    11'b01010010011: data <= 32'h3b52b085;
    11'b01010010100: data <= 32'h3a0524ae;
    11'b01010010101: data <= 32'hae3aaf85;
    11'b01010010110: data <= 32'h359125c7;
    11'b01010010111: data <= 32'h3ef23c65;
    11'b01010011000: data <= 32'h3ff74020;
    11'b01010011001: data <= 32'h38853d1d;
    11'b01010011010: data <= 32'hba53ba82;
    11'b01010011011: data <= 32'hb994bfad;
    11'b01010011100: data <= 32'h2fd0bc7d;
    11'b01010011101: data <= 32'h3780b229;
    11'b01010011110: data <= 32'h3824ba51;
    11'b01010011111: data <= 32'h3af4bf72;
    11'b01010100000: data <= 32'h3b39bd3f;
    11'b01010100001: data <= 32'hb4b9392b;
    11'b01010100010: data <= 32'hbfb43ec6;
    11'b01010100011: data <= 32'hc0523a11;
    11'b01010100100: data <= 32'hbb10b929;
    11'b01010100101: data <= 32'ha805bae7;
    11'b01010100110: data <= 32'hb921b384;
    11'b01010100111: data <= 32'hbcbd3096;
    11'b01010101000: data <= 32'ha15c367c;
    11'b01010101001: data <= 32'h3f5c3ce9;
    11'b01010101010: data <= 32'h3fdb400c;
    11'b01010101011: data <= 32'h30f23e3f;
    11'b01010101100: data <= 32'hbd0930a1;
    11'b01010101101: data <= 32'hb9c9b848;
    11'b01010101110: data <= 32'h393da696;
    11'b01010101111: data <= 32'h3cbd2df1;
    11'b01010110000: data <= 32'h3bd0bca5;
    11'b01010110001: data <= 32'h3c2fc086;
    11'b01010110010: data <= 32'h3cd7bd49;
    11'b01010110011: data <= 32'h38233aa1;
    11'b01010110100: data <= 32'hb9fe3e2c;
    11'b01010110101: data <= 32'hbcfd2a9f;
    11'b01010110110: data <= 32'hba52be4c;
    11'b01010110111: data <= 32'hb9a9be04;
    11'b01010111000: data <= 32'hbde7b74a;
    11'b01010111001: data <= 32'hbe7da4cd;
    11'b01010111010: data <= 32'had61af51;
    11'b01010111011: data <= 32'h3e823647;
    11'b01010111100: data <= 32'h3d103da8;
    11'b01010111101: data <= 32'hba6a3ee7;
    11'b01010111110: data <= 32'hbfb33c63;
    11'b01010111111: data <= 32'hbabe3916;
    11'b01011000000: data <= 32'h3a3c39df;
    11'b01011000001: data <= 32'h3c493531;
    11'b01011000010: data <= 32'h3856bc17;
    11'b01011000011: data <= 32'h3a00bf14;
    11'b01011000100: data <= 32'h3e66b862;
    11'b01011000101: data <= 32'h3e9e3d7a;
    11'b01011000110: data <= 32'h38d13ded;
    11'b01011000111: data <= 32'hb58eb68c;
    11'b01011001000: data <= 32'hb875bf9c;
    11'b01011001001: data <= 32'hba30bdda;
    11'b01011001010: data <= 32'hbd58b656;
    11'b01011001011: data <= 32'hbcc7b804;
    11'b01011001100: data <= 32'h32e7bd1f;
    11'b01011001101: data <= 32'h3d7cbbb9;
    11'b01011001110: data <= 32'h383d387c;
    11'b01011001111: data <= 32'hbdfe3ea0;
    11'b01011010000: data <= 32'hc0663dec;
    11'b01011010001: data <= 32'hbb323b5d;
    11'b01011010010: data <= 32'h361f39ae;
    11'b01011010011: data <= 32'h2cd634c8;
    11'b01011010100: data <= 32'hb935b8ec;
    11'b01011010101: data <= 32'h2cc9bb2a;
    11'b01011010110: data <= 32'h3f303578;
    11'b01011010111: data <= 32'h40d53f41;
    11'b01011011000: data <= 32'h3d3c3e1a;
    11'b01011011001: data <= 32'ha41eb415;
    11'b01011011010: data <= 32'hb61ebd0b;
    11'b01011011011: data <= 32'hb529b8a7;
    11'b01011011100: data <= 32'hb7db28ad;
    11'b01011011101: data <= 32'hb51cbbb2;
    11'b01011011110: data <= 32'h3924c0c3;
    11'b01011011111: data <= 32'h3d20c00d;
    11'b01011100000: data <= 32'h35a8a091;
    11'b01011100001: data <= 32'hbd393dbd;
    11'b01011100010: data <= 32'hbedb3c98;
    11'b01011100011: data <= 32'hb9b5344f;
    11'b01011100100: data <= 32'hb3ca265f;
    11'b01011100101: data <= 32'hbce22a08;
    11'b01011100110: data <= 32'hbfb2b4c7;
    11'b01011100111: data <= 32'hb8bdb5fe;
    11'b01011101000: data <= 32'h3ec638a2;
    11'b01011101001: data <= 32'h40c23ecb;
    11'b01011101010: data <= 32'h3c023e1d;
    11'b01011101011: data <= 32'hb6823652;
    11'b01011101100: data <= 32'hb64b25b9;
    11'b01011101101: data <= 32'h33a339a4;
    11'b01011101110: data <= 32'h352d3942;
    11'b01011101111: data <= 32'h3394bc5e;
    11'b01011110000: data <= 32'h3a2cc186;
    11'b01011110001: data <= 32'h3d64c054;
    11'b01011110010: data <= 32'h3b052a83;
    11'b01011110011: data <= 32'hb37d3cfa;
    11'b01011110100: data <= 32'hb8ea36e2;
    11'b01011110101: data <= 32'hb44cb9c5;
    11'b01011110110: data <= 32'hb933b994;
    11'b01011110111: data <= 32'hc00cb0d5;
    11'b01011111000: data <= 32'hc109b43f;
    11'b01011111001: data <= 32'hbab1b90f;
    11'b01011111010: data <= 32'h3da3b0b2;
    11'b01011111011: data <= 32'h3eb53b54;
    11'b01011111100: data <= 32'h24a63d59;
    11'b01011111101: data <= 32'hbc883c3b;
    11'b01011111110: data <= 32'hb80f3c9e;
    11'b01011111111: data <= 32'h38203e96;
    11'b01100000000: data <= 32'h370d3c6f;
    11'b01100000001: data <= 32'had61bac1;
    11'b01100000010: data <= 32'h353ec089;
    11'b01100000011: data <= 32'h3d93bd97;
    11'b01100000100: data <= 32'h3edd38fc;
    11'b01100000101: data <= 32'h3c483cbe;
    11'b01100000110: data <= 32'h37d4b0b0;
    11'b01100000111: data <= 32'h336abcff;
    11'b01100001000: data <= 32'hb88dba2f;
    11'b01100001001: data <= 32'hbf8a2704;
    11'b01100001010: data <= 32'hc043b6e0;
    11'b01100001011: data <= 32'hb851be00;
    11'b01100001100: data <= 32'h3c9cbdcc;
    11'b01100001101: data <= 32'h3ad6b0f3;
    11'b01100001110: data <= 32'hbaca3baf;
    11'b01100001111: data <= 32'hbe1a3d08;
    11'b01100010000: data <= 32'hb79f3dc1;
    11'b01100010001: data <= 32'h367e3ed2;
    11'b01100010010: data <= 32'hb43d3c86;
    11'b01100010011: data <= 32'hbcdbb6cb;
    11'b01100010100: data <= 32'hb889bd52;
    11'b01100010101: data <= 32'h3d06b5da;
    11'b01100010110: data <= 32'h40853cbb;
    11'b01100010111: data <= 32'h3f1c3caf;
    11'b01100011000: data <= 32'h3b8eb3d2;
    11'b01100011001: data <= 32'h380fbb13;
    11'b01100011010: data <= 32'had50288c;
    11'b01100011011: data <= 32'hbbf8395d;
    11'b01100011100: data <= 32'hbc97b855;
    11'b01100011101: data <= 32'h9d91c0b9;
    11'b01100011110: data <= 32'h3c1ec104;
    11'b01100011111: data <= 32'h3760bb16;
    11'b01100100000: data <= 32'hbb5a38a8;
    11'b01100100001: data <= 32'hbc7f3ae1;
    11'b01100100010: data <= 32'hae323a15;
    11'b01100100011: data <= 32'h30153b97;
    11'b01100100100: data <= 32'hbd3b3a51;
    11'b01100100101: data <= 32'hc0f7ae07;
    11'b01100100110: data <= 32'hbdb6b903;
    11'b01100100111: data <= 32'h3b8c2fa9;
    11'b01100101000: data <= 32'h40403cad;
    11'b01100101001: data <= 32'h3dd13c05;
    11'b01100101010: data <= 32'h38342c52;
    11'b01100101011: data <= 32'h37023060;
    11'b01100101100: data <= 32'h37bd3d44;
    11'b01100101101: data <= 32'ha7b33e0a;
    11'b01100101110: data <= 32'hb5c5b6ac;
    11'b01100101111: data <= 32'h33b7c138;
    11'b01100110000: data <= 32'h3bb0c149;
    11'b01100110001: data <= 32'h3950bac2;
    11'b01100110010: data <= 32'haf563686;
    11'b01100110011: data <= 32'ha8c03036;
    11'b01100110100: data <= 32'h38a9b5a9;
    11'b01100110101: data <= 32'h21b52499;
    11'b01100110110: data <= 32'hbfd13769;
    11'b01100110111: data <= 32'hc22b293d;
    11'b01100111000: data <= 32'hbef4b8b3;
    11'b01100111001: data <= 32'h3902b55d;
    11'b01100111010: data <= 32'h3d98369e;
    11'b01100111011: data <= 32'h35ed389c;
    11'b01100111100: data <= 32'hb61836a1;
    11'b01100111101: data <= 32'h32353c5c;
    11'b01100111110: data <= 32'h3aa8408e;
    11'b01100111111: data <= 32'h35b44027;
    11'b01101000000: data <= 32'hb68cad69;
    11'b01101000001: data <= 32'hb0f7c025;
    11'b01101000010: data <= 32'h3a3abf2f;
    11'b01101000011: data <= 32'h3cafb000;
    11'b01101000100: data <= 32'h3bf2377f;
    11'b01101000101: data <= 32'h3c64b7e9;
    11'b01101000110: data <= 32'h3cfabc7f;
    11'b01101000111: data <= 32'h3356b53d;
    11'b01101001000: data <= 32'hbf02388f;
    11'b01101001001: data <= 32'hc1492d51;
    11'b01101001010: data <= 32'hbd57bc7c;
    11'b01101001011: data <= 32'h3781bdb2;
    11'b01101001100: data <= 32'h384fb989;
    11'b01101001101: data <= 32'hb9b69492;
    11'b01101001110: data <= 32'hbc2736d2;
    11'b01101001111: data <= 32'h302c3d2b;
    11'b01101010000: data <= 32'h3b34409d;
    11'b01101010001: data <= 32'ha57e4014;
    11'b01101010010: data <= 32'hbd3e3441;
    11'b01101010011: data <= 32'hbc51bc6b;
    11'b01101010100: data <= 32'h369db88f;
    11'b01101010101: data <= 32'h3df03988;
    11'b01101010110: data <= 32'h3e62388b;
    11'b01101010111: data <= 32'h3e33b9ef;
    11'b01101011000: data <= 32'h3e11bc4d;
    11'b01101011001: data <= 32'h397e33b1;
    11'b01101011010: data <= 32'hbaa53ceb;
    11'b01101011011: data <= 32'hbdf432bb;
    11'b01101011100: data <= 32'hb878bedf;
    11'b01101011101: data <= 32'h3790c0b8;
    11'b01101011110: data <= 32'h25b6bdc8;
    11'b01101011111: data <= 32'hbc5bb6f3;
    11'b01101100000: data <= 32'hbb1f20c1;
    11'b01101100001: data <= 32'h380e389b;
    11'b01101100010: data <= 32'h3ae33da4;
    11'b01101100011: data <= 32'hba383dee;
    11'b01101100100: data <= 32'hc0e23774;
    11'b01101100101: data <= 32'hbfedb4ce;
    11'b01101100110: data <= 32'ha01c32a8;
    11'b01101100111: data <= 32'h3d1d3b8d;
    11'b01101101000: data <= 32'h3ce836e1;
    11'b01101101001: data <= 32'h3c17b946;
    11'b01101101010: data <= 32'h3d13b5ae;
    11'b01101101011: data <= 32'h3c863d77;
    11'b01101101100: data <= 32'h32f1403f;
    11'b01101101101: data <= 32'hb6c737d5;
    11'b01101101110: data <= 32'ha83dbf64;
    11'b01101101111: data <= 32'h375bc0df;
    11'b01101110000: data <= 32'h222abd52;
    11'b01101110001: data <= 32'hb8c1b7a8;
    11'b01101110010: data <= 32'h267eb8f3;
    11'b01101110011: data <= 32'h3cfcb8db;
    11'b01101110100: data <= 32'h3b7b3307;
    11'b01101110101: data <= 32'hbd0f3af8;
    11'b01101110110: data <= 32'hc1f33822;
    11'b01101110111: data <= 32'hc082ac63;
    11'b01101111000: data <= 32'hb3ff2c76;
    11'b01101111001: data <= 32'h38f53618;
    11'b01101111010: data <= 32'h2d20aafc;
    11'b01101111011: data <= 32'hafadb83a;
    11'b01101111100: data <= 32'h39f5367b;
    11'b01101111101: data <= 32'h3d7e4082;
    11'b01101111110: data <= 32'h3a30415f;
    11'b01101111111: data <= 32'hb0de3a6d;
    11'b01110000000: data <= 32'hb2c4bd5c;
    11'b01110000001: data <= 32'h33a0be1f;
    11'b01110000010: data <= 32'h349fb66d;
    11'b01110000011: data <= 32'h34a3b0f1;
    11'b01110000100: data <= 32'h3c4fbc83;
    11'b01110000101: data <= 32'h3fc1be1c;
    11'b01110000110: data <= 32'h3cc3b721;
    11'b01110000111: data <= 32'hbc3539de;
    11'b01110001000: data <= 32'hc0f33894;
    11'b01110001001: data <= 32'hbeb2b5e6;
    11'b01110001010: data <= 32'hb17fba29;
    11'b01110001011: data <= 32'haff2b908;
    11'b01110001100: data <= 32'hbc8db983;
    11'b01110001101: data <= 32'hbc60b8dc;
    11'b01110001110: data <= 32'h36a13876;
    11'b01110001111: data <= 32'h3db44076;
    11'b01110010000: data <= 32'h38fb4107;
    11'b01110010001: data <= 32'hba433ba8;
    11'b01110010010: data <= 32'hbc14b7a0;
    11'b01110010011: data <= 32'hb25cb1d2;
    11'b01110010100: data <= 32'h377139cc;
    11'b01110010101: data <= 32'h3a73334c;
    11'b01110010110: data <= 32'h3defbd54;
    11'b01110010111: data <= 32'h403dbec8;
    11'b01110011000: data <= 32'h3e00b156;
    11'b01110011001: data <= 32'hb2fa3d03;
    11'b01110011010: data <= 32'hbcd73a2f;
    11'b01110011011: data <= 32'hb8ccba5a;
    11'b01110011100: data <= 32'h2fe5be56;
    11'b01110011101: data <= 32'hb899bd5b;
    11'b01110011110: data <= 32'hbee0bc4f;
    11'b01110011111: data <= 32'hbd01bb74;
    11'b01110100000: data <= 32'h38faae24;
    11'b01110100001: data <= 32'h3dcd3cf0;
    11'b01110100010: data <= 32'h2bcc3eb7;
    11'b01110100011: data <= 32'hbf093af0;
    11'b01110100100: data <= 32'hbf8333dd;
    11'b01110100101: data <= 32'hb8f33a58;
    11'b01110100110: data <= 32'h34b63d32;
    11'b01110100111: data <= 32'h378834a2;
    11'b01110101000: data <= 32'h3afabd30;
    11'b01110101001: data <= 32'h3e83bcba;
    11'b01110101010: data <= 32'h3eae3a39;
    11'b01110101011: data <= 32'h39e84031;
    11'b01110101100: data <= 32'h29733c56;
    11'b01110101101: data <= 32'h3431bb3e;
    11'b01110101110: data <= 32'h3579bea7;
    11'b01110101111: data <= 32'hb8e3bc9f;
    11'b01110110000: data <= 32'hbdc3bb5e;
    11'b01110110001: data <= 32'hb85bbd43;
    11'b01110110010: data <= 32'h3d31bcc0;
    11'b01110110011: data <= 32'h3e53b03e;
    11'b01110110100: data <= 32'hb5c839ca;
    11'b01110110101: data <= 32'hc0883941;
    11'b01110110110: data <= 32'hc03137ab;
    11'b01110110111: data <= 32'hb9a83b06;
    11'b01110111000: data <= 32'hb12e3bcd;
    11'b01110111001: data <= 32'hb8beaf1b;
    11'b01110111010: data <= 32'hb6f2bcf2;
    11'b01110111011: data <= 32'h3a19b833;
    11'b01110111100: data <= 32'h3e853e74;
    11'b01110111101: data <= 32'h3d18413e;
    11'b01110111110: data <= 32'h38543d2d;
    11'b01110111111: data <= 32'h35adb86d;
    11'b01111000000: data <= 32'h337eba9b;
    11'b01111000001: data <= 32'hb686ad0e;
    11'b01111000010: data <= 32'hb98ab454;
    11'b01111000011: data <= 32'h36dfbe24;
    11'b01111000100: data <= 32'h3fdbc022;
    11'b01111000101: data <= 32'h3f1fbc1a;
    11'b01111000110: data <= 32'hb41a3489;
    11'b01111000111: data <= 32'hbf483880;
    11'b01111001000: data <= 32'hbd8c33df;
    11'b01111001001: data <= 32'hb542326e;
    11'b01111001010: data <= 32'hb8fa2c99;
    11'b01111001011: data <= 32'hbf0ab9ce;
    11'b01111001100: data <= 32'hbe8abd35;
    11'b01111001101: data <= 32'h2e9db4ff;
    11'b01111001110: data <= 32'h3dfa3e82;
    11'b01111001111: data <= 32'h3cb340ae;
    11'b01111010000: data <= 32'h2e1e3cbb;
    11'b01111010001: data <= 32'hb50329ae;
    11'b01111010010: data <= 32'hb1b5377e;
    11'b01111010011: data <= 32'hb40f3d16;
    11'b01111010100: data <= 32'hb12b375c;
    11'b01111010101: data <= 32'h3adebe11;
    11'b01111010110: data <= 32'h4022c08a;
    11'b01111010111: data <= 32'h3f78bb9a;
    11'b01111011000: data <= 32'h35693900;
    11'b01111011001: data <= 32'hb8e039c7;
    11'b01111011010: data <= 32'hae0eb043;
    11'b01111011011: data <= 32'h3534b8ae;
    11'b01111011100: data <= 32'hba9ab928;
    11'b01111011101: data <= 32'hc0b8bc41;
    11'b01111011110: data <= 32'hc006bdd1;
    11'b01111011111: data <= 32'h2e09ba14;
    11'b01111100000: data <= 32'h3dce397a;
    11'b01111100001: data <= 32'h395d3d34;
    11'b01111100010: data <= 32'hba8739e0;
    11'b01111100011: data <= 32'hbca03805;
    11'b01111100100: data <= 32'hb8903dce;
    11'b01111100101: data <= 32'hb4e0402a;
    11'b01111100110: data <= 32'hb5463a39;
    11'b01111100111: data <= 32'h34ccbd86;
    11'b01111101000: data <= 32'h3d91bf44;
    11'b01111101001: data <= 32'h3ec5ae92;
    11'b01111101010: data <= 32'h3c183db6;
    11'b01111101011: data <= 32'h39253c14;
    11'b01111101100: data <= 32'h3c12b511;
    11'b01111101101: data <= 32'h3ab7ba54;
    11'b01111101110: data <= 32'hb9d0b817;
    11'b01111101111: data <= 32'hc048ba07;
    11'b01111110000: data <= 32'hbdbbbe16;
    11'b01111110001: data <= 32'h3999be56;
    11'b01111110010: data <= 32'h3e48b965;
    11'b01111110011: data <= 32'h32d82d66;
    11'b01111110100: data <= 32'hbda53232;
    11'b01111110101: data <= 32'hbdb03889;
    11'b01111110110: data <= 32'hb8513e5d;
    11'b01111110111: data <= 32'hb7be3fab;
    11'b01111111000: data <= 32'hbc9037bc;
    11'b01111111001: data <= 32'hbbeebd37;
    11'b01111111010: data <= 32'h343bbc9e;
    11'b01111111011: data <= 32'h3d313a47;
    11'b01111111100: data <= 32'h3d6e3ff9;
    11'b01111111101: data <= 32'h3cc53c92;
    11'b01111111110: data <= 32'h3d36b251;
    11'b01111111111: data <= 32'h3b0cb1dd;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    