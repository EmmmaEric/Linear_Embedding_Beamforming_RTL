
module memory_rom_19(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3d1e3b81;
    11'b00000000001: data <= 32'h39b13788;
    11'b00000000010: data <= 32'hba0ab8fb;
    11'b00000000011: data <= 32'hba67bec8;
    11'b00000000100: data <= 32'h3bb5bdc3;
    11'b00000000101: data <= 32'h40b8b0fa;
    11'b00000000110: data <= 32'h3f173581;
    11'b00000000111: data <= 32'h31aeb848;
    11'b00000001000: data <= 32'hb9d0bc95;
    11'b00000001001: data <= 32'hbb43b326;
    11'b00000001010: data <= 32'hbd143b41;
    11'b00000001011: data <= 32'hbe80340c;
    11'b00000001100: data <= 32'hbc42be78;
    11'b00000001101: data <= 32'h2c35c049;
    11'b00000001110: data <= 32'h35c3b68f;
    11'b00000001111: data <= 32'hb5cc3e80;
    11'b00000010000: data <= 32'hb8f74005;
    11'b00000010001: data <= 32'h34393d06;
    11'b00000010010: data <= 32'h3aa73b2a;
    11'b00000010011: data <= 32'hb2d13bce;
    11'b00000010100: data <= 32'hbe5537cd;
    11'b00000010101: data <= 32'hbbffb76f;
    11'b00000010110: data <= 32'h3d6cb9b6;
    11'b00000010111: data <= 32'h41b6af76;
    11'b00000011000: data <= 32'h40102fb5;
    11'b00000011001: data <= 32'h360eb6da;
    11'b00000011010: data <= 32'hb087b88e;
    11'b00000011011: data <= 32'h324035a7;
    11'b00000011100: data <= 32'haca83b37;
    11'b00000011101: data <= 32'hbbaeb6b2;
    11'b00000011110: data <= 32'hbcb2c0f8;
    11'b00000011111: data <= 32'hb725c173;
    11'b00000100000: data <= 32'h2bdbb9d4;
    11'b00000100001: data <= 32'hb2283c8f;
    11'b00000100010: data <= 32'hb5443c71;
    11'b00000100011: data <= 32'h2e763427;
    11'b00000100100: data <= 32'h255636d0;
    11'b00000100101: data <= 32'hbd193d57;
    11'b00000100110: data <= 32'hc0ab3d5e;
    11'b00000100111: data <= 32'hbd37335c;
    11'b00000101000: data <= 32'h3c81b840;
    11'b00000101001: data <= 32'h40acb23d;
    11'b00000101010: data <= 32'h3d833567;
    11'b00000101011: data <= 32'h314b35a9;
    11'b00000101100: data <= 32'h37703792;
    11'b00000101101: data <= 32'h3d693c59;
    11'b00000101110: data <= 32'h3b893c48;
    11'b00000101111: data <= 32'hb862b83f;
    11'b00000110000: data <= 32'hbcc5c0e0;
    11'b00000110001: data <= 32'hb554c0fa;
    11'b00000110010: data <= 32'h3936ba28;
    11'b00000110011: data <= 32'h393c362a;
    11'b00000110100: data <= 32'h333cb283;
    11'b00000110101: data <= 32'h29aabb74;
    11'b00000110110: data <= 32'hb70eac86;
    11'b00000110111: data <= 32'hbeb33dd6;
    11'b00000111000: data <= 32'hc0fb3e03;
    11'b00000111001: data <= 32'hbe26a682;
    11'b00000111010: data <= 32'h35eabc51;
    11'b00000111011: data <= 32'h3c4cb805;
    11'b00000111100: data <= 32'h32ac391b;
    11'b00000111101: data <= 32'hb45b3c6f;
    11'b00000111110: data <= 32'h3a763ccd;
    11'b00000111111: data <= 32'h3f9c3e02;
    11'b00001000000: data <= 32'h3c763d7e;
    11'b00001000001: data <= 32'hba1d2d12;
    11'b00001000010: data <= 32'hbd2abdb5;
    11'b00001000011: data <= 32'h3017be29;
    11'b00001000100: data <= 32'h3e50b822;
    11'b00001000101: data <= 32'h3e32b2ec;
    11'b00001000110: data <= 32'h39c1bc98;
    11'b00001000111: data <= 32'h3404be26;
    11'b00001001000: data <= 32'haf3db0e4;
    11'b00001001001: data <= 32'hbc2d3dd3;
    11'b00001001010: data <= 32'hbf903c35;
    11'b00001001011: data <= 32'hbe2dbb8f;
    11'b00001001100: data <= 32'hb770bfe6;
    11'b00001001101: data <= 32'hb140bb54;
    11'b00001001110: data <= 32'hb9c1395d;
    11'b00001001111: data <= 32'hb8703ca8;
    11'b00001010000: data <= 32'h3ab03c03;
    11'b00001010001: data <= 32'h3e9c3d15;
    11'b00001010010: data <= 32'h368d3e7d;
    11'b00001010011: data <= 32'hbe063c3f;
    11'b00001010100: data <= 32'hbe21ab3f;
    11'b00001010101: data <= 32'h374bb7af;
    11'b00001010110: data <= 32'h401ab21f;
    11'b00001010111: data <= 32'h3f11b66b;
    11'b00001011000: data <= 32'h3a37bcf7;
    11'b00001011001: data <= 32'h38febcd4;
    11'b00001011010: data <= 32'h3afd350a;
    11'b00001011011: data <= 32'h347c3e04;
    11'b00001011100: data <= 32'hbb2d37b6;
    11'b00001011101: data <= 32'hbd63bf07;
    11'b00001011110: data <= 32'hbb4ec10b;
    11'b00001011111: data <= 32'hb94bbc8d;
    11'b00001100000: data <= 32'hba98358e;
    11'b00001100001: data <= 32'hb67135c8;
    11'b00001100010: data <= 32'h39caaed9;
    11'b00001100011: data <= 32'h3bc837cc;
    11'b00001100100: data <= 32'hb8893ead;
    11'b00001100101: data <= 32'hc0753f55;
    11'b00001100110: data <= 32'hbf223aad;
    11'b00001100111: data <= 32'h35671e05;
    11'b00001101000: data <= 32'h3e6cadf0;
    11'b00001101001: data <= 32'h3c0db32b;
    11'b00001101010: data <= 32'h346cb8ea;
    11'b00001101011: data <= 32'h3b67b47a;
    11'b00001101100: data <= 32'h3fbe3c14;
    11'b00001101101: data <= 32'h3df33ea2;
    11'b00001101110: data <= 32'hb10834ee;
    11'b00001101111: data <= 32'hbc98bf0c;
    11'b00001110000: data <= 32'hba91c068;
    11'b00001110001: data <= 32'hb3debb68;
    11'b00001110010: data <= 32'hb012afd6;
    11'b00001110011: data <= 32'h2f58bad7;
    11'b00001110100: data <= 32'h3979bdf1;
    11'b00001110101: data <= 32'h37f0b5a9;
    11'b00001110110: data <= 32'hbbfc3e2a;
    11'b00001110111: data <= 32'hc0a53ff8;
    11'b00001111000: data <= 32'hbf3a3a23;
    11'b00001111001: data <= 32'hb146b5ac;
    11'b00001111010: data <= 32'h3701b579;
    11'b00001111011: data <= 32'hb56628ff;
    11'b00001111100: data <= 32'hb81c2f32;
    11'b00001111101: data <= 32'h3bed3750;
    11'b00001111110: data <= 32'h40ee3d96;
    11'b00001111111: data <= 32'h3f703f32;
    11'b00010000000: data <= 32'hb0c0399b;
    11'b00010000001: data <= 32'hbca2bab6;
    11'b00010000010: data <= 32'hb67cbc58;
    11'b00010000011: data <= 32'h38efb529;
    11'b00010000100: data <= 32'h3a04b6e5;
    11'b00010000101: data <= 32'h38b3bf0e;
    11'b00010000110: data <= 32'h3a3cc09a;
    11'b00010000111: data <= 32'h392fb997;
    11'b00010001000: data <= 32'hb7333da8;
    11'b00010001001: data <= 32'hbe4c3e56;
    11'b00010001010: data <= 32'hbde9ab42;
    11'b00010001011: data <= 32'hb99bbcd3;
    11'b00010001100: data <= 32'hba09b9f4;
    11'b00010001101: data <= 32'hbdf23065;
    11'b00010001110: data <= 32'hbc6234ce;
    11'b00010001111: data <= 32'h3ada3558;
    11'b00010010000: data <= 32'h407f3c2a;
    11'b00010010001: data <= 32'h3d1b3ef5;
    11'b00010010010: data <= 32'hba813d90;
    11'b00010010011: data <= 32'hbd8c37a4;
    11'b00010010100: data <= 32'haa0e327b;
    11'b00010010101: data <= 32'h3cb5355b;
    11'b00010010110: data <= 32'h3c22b6ad;
    11'b00010010111: data <= 32'h3869bf87;
    11'b00010011000: data <= 32'h3b12c03d;
    11'b00010011001: data <= 32'h3d70b588;
    11'b00010011010: data <= 32'h3a853dbe;
    11'b00010011011: data <= 32'hb5a43c0a;
    11'b00010011100: data <= 32'hbb66bb5a;
    11'b00010011101: data <= 32'hbb57bf38;
    11'b00010011110: data <= 32'hbd13bb35;
    11'b00010011111: data <= 32'hbf1328ae;
    11'b00010100000: data <= 32'hbc68b40d;
    11'b00010100001: data <= 32'h3997b9b4;
    11'b00010100010: data <= 32'h3e552933;
    11'b00010100011: data <= 32'h348b3daf;
    11'b00010100100: data <= 32'hbe4c3f9e;
    11'b00010100101: data <= 32'hbe653d81;
    11'b00010100110: data <= 32'h21953b27;
    11'b00010100111: data <= 32'h3b9c391d;
    11'b00010101000: data <= 32'h3588b148;
    11'b00010101001: data <= 32'hb0babd1f;
    11'b00010101010: data <= 32'h3a9abcd9;
    11'b00010101011: data <= 32'h404c3611;
    11'b00010101100: data <= 32'h400a3e48;
    11'b00010101101: data <= 32'h38ee399f;
    11'b00010101110: data <= 32'hb78fbc73;
    11'b00010101111: data <= 32'hb9b8be39;
    11'b00010110000: data <= 32'hbb14b820;
    11'b00010110001: data <= 32'hbc82ade2;
    11'b00010110010: data <= 32'hb8babcc9;
    11'b00010110011: data <= 32'h3935c02b;
    11'b00010110100: data <= 32'h3c0bbc2f;
    11'b00010110101: data <= 32'hb4e33bf8;
    11'b00010110110: data <= 32'hbef83fab;
    11'b00010110111: data <= 32'hbdeb3d5f;
    11'b00010111000: data <= 32'hb1b43907;
    11'b00010111001: data <= 32'h2a7436f3;
    11'b00010111010: data <= 32'hbbef2ed3;
    11'b00010111011: data <= 32'hbcc6b7e1;
    11'b00010111100: data <= 32'h387db58d;
    11'b00010111101: data <= 32'h40ff3aab;
    11'b00010111110: data <= 32'h40db3e69;
    11'b00010111111: data <= 32'h3a133a87;
    11'b00011000000: data <= 32'hb642b720;
    11'b00011000001: data <= 32'hb471b750;
    11'b00011000010: data <= 32'h2209357e;
    11'b00011000011: data <= 32'hb0e8aa7b;
    11'b00011000100: data <= 32'ha94dbf9a;
    11'b00011000101: data <= 32'h3961c1de;
    11'b00011000110: data <= 32'h3b63be42;
    11'b00011000111: data <= 32'h8ae139d2;
    11'b00011001000: data <= 32'hbc173ddb;
    11'b00011001001: data <= 32'hbb3c3809;
    11'b00011001010: data <= 32'hb5b0b481;
    11'b00011001011: data <= 32'hbb5ca84d;
    11'b00011001100: data <= 32'hc05b33fd;
    11'b00011001101: data <= 32'hbfefaeb6;
    11'b00011001110: data <= 32'h3389b3c4;
    11'b00011001111: data <= 32'h406c3832;
    11'b00011010000: data <= 32'h3f613d48;
    11'b00011010001: data <= 32'h2cca3c9a;
    11'b00011010010: data <= 32'hb950391a;
    11'b00011010011: data <= 32'h2edb3af9;
    11'b00011010100: data <= 32'h39df3cf7;
    11'b00011010101: data <= 32'h3564327a;
    11'b00011010110: data <= 32'ha32dbfad;
    11'b00011010111: data <= 32'h38afc18a;
    11'b00011011000: data <= 32'h3d2dbcee;
    11'b00011011001: data <= 32'h3c193a1b;
    11'b00011011010: data <= 32'h33893af4;
    11'b00011011011: data <= 32'had8ab7ca;
    11'b00011011100: data <= 32'hb4a7bc45;
    11'b00011011101: data <= 32'hbd3db449;
    11'b00011011110: data <= 32'hc0fc34dc;
    11'b00011011111: data <= 32'hc01db57c;
    11'b00011100000: data <= 32'h2ab0bc30;
    11'b00011100001: data <= 32'h3e16b806;
    11'b00011100010: data <= 32'h3a0239ce;
    11'b00011100011: data <= 32'hbacd3d66;
    11'b00011100100: data <= 32'hbbb23d8d;
    11'b00011100101: data <= 32'h34923e72;
    11'b00011100110: data <= 32'h3a5b3ea9;
    11'b00011100111: data <= 32'haf0d3836;
    11'b00011101000: data <= 32'hb9cbbd24;
    11'b00011101001: data <= 32'h3411bf24;
    11'b00011101010: data <= 32'h3effb5f2;
    11'b00011101011: data <= 32'h40203be2;
    11'b00011101100: data <= 32'h3d113789;
    11'b00011101101: data <= 32'h3848bb80;
    11'b00011101110: data <= 32'h288fbc39;
    11'b00011101111: data <= 32'hbb082eef;
    11'b00011110000: data <= 32'hbf3636ec;
    11'b00011110001: data <= 32'hbdc9bb8e;
    11'b00011110010: data <= 32'h2d59c078;
    11'b00011110011: data <= 32'h3b10bea5;
    11'b00011110100: data <= 32'hac5e2d97;
    11'b00011110101: data <= 32'hbd023cbe;
    11'b00011110110: data <= 32'hbafd3d29;
    11'b00011110111: data <= 32'h35483d4d;
    11'b00011111000: data <= 32'h33693d9e;
    11'b00011111001: data <= 32'hbd0439e9;
    11'b00011111010: data <= 32'hbf5fb724;
    11'b00011111011: data <= 32'hb41ab9bd;
    11'b00011111100: data <= 32'h3f8234fe;
    11'b00011111101: data <= 32'h40c53c49;
    11'b00011111110: data <= 32'h3dab3611;
    11'b00011111111: data <= 32'h38e8b8cb;
    11'b00100000000: data <= 32'h3724b123;
    11'b00100000001: data <= 32'h2bb03c26;
    11'b00100000010: data <= 32'hb93c39ef;
    11'b00100000011: data <= 32'hb96cbd90;
    11'b00100000100: data <= 32'h31c7c1f8;
    11'b00100000101: data <= 32'h38f7c06d;
    11'b00100000110: data <= 32'had19b37e;
    11'b00100000111: data <= 32'hb9fb39bd;
    11'b00100001000: data <= 32'hb3b0368f;
    11'b00100001001: data <= 32'h36e43456;
    11'b00100001010: data <= 32'hb74839e6;
    11'b00100001011: data <= 32'hc0a83a59;
    11'b00100001100: data <= 32'hc1632d65;
    11'b00100001101: data <= 32'hb985b4fb;
    11'b00100001110: data <= 32'h3e1b335f;
    11'b00100001111: data <= 32'h3f063a04;
    11'b00100010000: data <= 32'h38f636ff;
    11'b00100010001: data <= 32'h318531d0;
    11'b00100010010: data <= 32'h39ee3c2d;
    11'b00100010011: data <= 32'h3b314009;
    11'b00100010100: data <= 32'h2fa53c9e;
    11'b00100010101: data <= 32'hb693bd34;
    11'b00100010110: data <= 32'h2d68c188;
    11'b00100010111: data <= 32'h39d2bf36;
    11'b00100011000: data <= 32'h390cac89;
    11'b00100011001: data <= 32'h35fc3264;
    11'b00100011010: data <= 32'h3967b96e;
    11'b00100011011: data <= 32'h3998ba3b;
    11'b00100011100: data <= 32'hb98e3419;
    11'b00100011101: data <= 32'hc12b3a9d;
    11'b00100011110: data <= 32'hc1742da7;
    11'b00100011111: data <= 32'hba5bba5d;
    11'b00100100000: data <= 32'h3b23b924;
    11'b00100100001: data <= 32'h389c2b04;
    11'b00100100010: data <= 32'hb85f365a;
    11'b00100100011: data <= 32'hb5f339f3;
    11'b00100100100: data <= 32'h3afd3ee4;
    11'b00100100101: data <= 32'h3cb440e1;
    11'b00100100110: data <= 32'h9ed23dd0;
    11'b00100100111: data <= 32'hbb92b98a;
    11'b00100101000: data <= 32'hb573bed2;
    11'b00100101001: data <= 32'h3b61b9cc;
    11'b00100101010: data <= 32'h3dca363b;
    11'b00100101011: data <= 32'h3d5bb04a;
    11'b00100101100: data <= 32'h3d58bd4a;
    11'b00100101101: data <= 32'h3c3ebc58;
    11'b00100101110: data <= 32'hb40f36fb;
    11'b00100101111: data <= 32'hbf4c3c1f;
    11'b00100110000: data <= 32'hbfb6b3cc;
    11'b00100110001: data <= 32'hb857bef1;
    11'b00100110010: data <= 32'h3539bee8;
    11'b00100110011: data <= 32'hb6aab941;
    11'b00100110100: data <= 32'hbd0e307f;
    11'b00100110101: data <= 32'hb80138c7;
    11'b00100110110: data <= 32'h3bc03d81;
    11'b00100110111: data <= 32'h3b0a4010;
    11'b00100111000: data <= 32'hbb113de7;
    11'b00100111001: data <= 32'hbfeb2ca9;
    11'b00100111010: data <= 32'hbb96b7b1;
    11'b00100111011: data <= 32'h3b3c3453;
    11'b00100111100: data <= 32'h3ebc39b4;
    11'b00100111101: data <= 32'h3dc0b3fe;
    11'b00100111110: data <= 32'h3d41bcf9;
    11'b00100111111: data <= 32'h3d4cb791;
    11'b00101000000: data <= 32'h38f83d0e;
    11'b00101000001: data <= 32'hb84a3dcc;
    11'b00101000010: data <= 32'hbaddb809;
    11'b00101000011: data <= 32'hb230c0ba;
    11'b00101000100: data <= 32'h2c4bc077;
    11'b00101000101: data <= 32'hb96abb68;
    11'b00101000110: data <= 32'hbc3bb382;
    11'b00101000111: data <= 32'h21a4b399;
    11'b00101001000: data <= 32'h3cb93254;
    11'b00101001001: data <= 32'h36893c54;
    11'b00101001010: data <= 32'hbf393d17;
    11'b00101001011: data <= 32'hc194389d;
    11'b00101001100: data <= 32'hbd813133;
    11'b00101001101: data <= 32'h38bb3806;
    11'b00101001110: data <= 32'h3c4b3855;
    11'b00101001111: data <= 32'h3842b4bd;
    11'b00101010000: data <= 32'h38f3b996;
    11'b00101010001: data <= 32'h3d7a3870;
    11'b00101010010: data <= 32'h3daa406a;
    11'b00101010011: data <= 32'h37633f98;
    11'b00101010100: data <= 32'hb434b65b;
    11'b00101010101: data <= 32'haeffc046;
    11'b00101010110: data <= 32'h2d8bbeec;
    11'b00101010111: data <= 32'hb2eab85f;
    11'b00101011000: data <= 32'hb070b831;
    11'b00101011001: data <= 32'h3b19bd1b;
    11'b00101011010: data <= 32'h3e17bc3f;
    11'b00101011011: data <= 32'h339c343d;
    11'b00101011100: data <= 32'hc00e3c61;
    11'b00101011101: data <= 32'hc17f3928;
    11'b00101011110: data <= 32'hbd3dac21;
    11'b00101011111: data <= 32'h30d7b07d;
    11'b00101100000: data <= 32'hab92aebd;
    11'b00101100001: data <= 32'hbaa6b6f6;
    11'b00101100010: data <= 32'hb432b402;
    11'b00101100011: data <= 32'h3d113cb3;
    11'b00101100100: data <= 32'h3eed4127;
    11'b00101100101: data <= 32'h38c24027;
    11'b00101100110: data <= 32'hb8522b87;
    11'b00101100111: data <= 32'hb767bc74;
    11'b00101101000: data <= 32'h3167b784;
    11'b00101101001: data <= 32'h372933c1;
    11'b00101101010: data <= 32'h39f5b8df;
    11'b00101101011: data <= 32'h3e11bfc0;
    11'b00101101100: data <= 32'h3f43be83;
    11'b00101101101: data <= 32'h3894311c;
    11'b00101101110: data <= 32'hbd2f3cca;
    11'b00101101111: data <= 32'hbf2536cd;
    11'b00101110000: data <= 32'hb9f9ba91;
    11'b00101110001: data <= 32'hb136bc77;
    11'b00101110010: data <= 32'hbc37ba65;
    11'b00101110011: data <= 32'hbf3ab967;
    11'b00101110100: data <= 32'hb99db572;
    11'b00101110101: data <= 32'h3ce83ac1;
    11'b00101110110: data <= 32'h3e28400f;
    11'b00101110111: data <= 32'haccf3f46;
    11'b00101111000: data <= 32'hbdc038a5;
    11'b00101111001: data <= 32'hbc3b2ea6;
    11'b00101111010: data <= 32'h2fd83a42;
    11'b00101111011: data <= 32'h39863b30;
    11'b00101111100: data <= 32'h3ac3b877;
    11'b00101111101: data <= 32'h3d89bfca;
    11'b00101111110: data <= 32'h3f5cbcf5;
    11'b00101111111: data <= 32'h3ce43a94;
    11'b00110000000: data <= 32'ha4ef3e65;
    11'b00110000001: data <= 32'hb769333b;
    11'b00110000010: data <= 32'haa1cbda5;
    11'b00110000011: data <= 32'hb33fbe71;
    11'b00110000100: data <= 32'hbd90bbeb;
    11'b00110000101: data <= 32'hbf5fbae6;
    11'b00110000110: data <= 32'hb633bbda;
    11'b00110000111: data <= 32'h3da1b51c;
    11'b00110001000: data <= 32'h3c9a3ab6;
    11'b00110001001: data <= 32'hbb5d3d07;
    11'b00110001010: data <= 32'hc0703aec;
    11'b00110001011: data <= 32'hbdbe3a7a;
    11'b00110001100: data <= 32'hab363d19;
    11'b00110001101: data <= 32'h338d3bb1;
    11'b00110001110: data <= 32'ha9ccb866;
    11'b00110001111: data <= 32'h3780bdfe;
    11'b00110010000: data <= 32'h3e25b529;
    11'b00110010001: data <= 32'h3f233ee1;
    11'b00110010010: data <= 32'h3c1d400b;
    11'b00110010011: data <= 32'h36843402;
    11'b00110010100: data <= 32'h34f3bd32;
    11'b00110010101: data <= 32'hafd9bc7b;
    11'b00110010110: data <= 32'hbc20b6af;
    11'b00110010111: data <= 32'hbc42ba9a;
    11'b00110011000: data <= 32'h36c0bf23;
    11'b00110011001: data <= 32'h3ef5be79;
    11'b00110011010: data <= 32'h3b8cb43b;
    11'b00110011011: data <= 32'hbce03a2a;
    11'b00110011100: data <= 32'hc0613a84;
    11'b00110011101: data <= 32'hbcd53979;
    11'b00110011110: data <= 32'hb2893a70;
    11'b00110011111: data <= 32'hb95f368e;
    11'b00110100000: data <= 32'hbdc4b97f;
    11'b00110100001: data <= 32'hb99dbc36;
    11'b00110100010: data <= 32'h3c613569;
    11'b00110100011: data <= 32'h3fcb4033;
    11'b00110100100: data <= 32'h3d094026;
    11'b00110100101: data <= 32'h355e374c;
    11'b00110100110: data <= 32'h2dabb7b7;
    11'b00110100111: data <= 32'ha85d3161;
    11'b00110101000: data <= 32'hb6723940;
    11'b00110101001: data <= 32'hb1aab872;
    11'b00110101010: data <= 32'h3c3ec089;
    11'b00110101011: data <= 32'h3fc8c08d;
    11'b00110101100: data <= 32'h3c4bb8d8;
    11'b00110101101: data <= 32'hb95e3993;
    11'b00110101110: data <= 32'hbcd23893;
    11'b00110101111: data <= 32'hb5f6a29e;
    11'b00110110000: data <= 32'hb11eb079;
    11'b00110110001: data <= 32'hbde3b499;
    11'b00110110010: data <= 32'hc102bb01;
    11'b00110110011: data <= 32'hbd9ebbe7;
    11'b00110110100: data <= 32'h3aaf3154;
    11'b00110110101: data <= 32'h3ed43e2a;
    11'b00110110110: data <= 32'h394f3e42;
    11'b00110110111: data <= 32'hb7e53905;
    11'b00110111000: data <= 32'hb7e73844;
    11'b00110111001: data <= 32'hab0f3e06;
    11'b00110111010: data <= 32'haab43e67;
    11'b00110111011: data <= 32'h2b37b3c5;
    11'b00110111100: data <= 32'h3b6fc067;
    11'b00110111101: data <= 32'h3f01bfe5;
    11'b00110111110: data <= 32'h3d93aa45;
    11'b00110111111: data <= 32'h366f3c3d;
    11'b00111000000: data <= 32'h327435cc;
    11'b00111000001: data <= 32'h3911b958;
    11'b00111000010: data <= 32'h2cdbb9e7;
    11'b00111000011: data <= 32'hbed3b7e1;
    11'b00111000100: data <= 32'hc145bb13;
    11'b00111000101: data <= 32'hbcf1bd51;
    11'b00111000110: data <= 32'h3b8fba60;
    11'b00111000111: data <= 32'h3d3f3460;
    11'b00111001000: data <= 32'hb2c83980;
    11'b00111001001: data <= 32'hbd6638aa;
    11'b00111001010: data <= 32'hbb2a3c74;
    11'b00111001011: data <= 32'hae4b4035;
    11'b00111001100: data <= 32'hb3e93f66;
    11'b00111001101: data <= 32'hb925afe9;
    11'b00111001110: data <= 32'haa5ebef5;
    11'b00111001111: data <= 32'h3c8abc37;
    11'b00111010000: data <= 32'h3e6f3b26;
    11'b00111010001: data <= 32'h3d393e09;
    11'b00111010010: data <= 32'h3cc034a1;
    11'b00111010011: data <= 32'h3ce1ba31;
    11'b00111010100: data <= 32'h355fb6d1;
    11'b00111010101: data <= 32'hbd493010;
    11'b00111010110: data <= 32'hbf87b86b;
    11'b00111010111: data <= 32'hb69ebf20;
    11'b00111011000: data <= 32'h3d31bfc0;
    11'b00111011001: data <= 32'h3c26bb9e;
    11'b00111011010: data <= 32'hb982ac6d;
    11'b00111011011: data <= 32'hbdef3542;
    11'b00111011100: data <= 32'hb91d3b91;
    11'b00111011101: data <= 32'h25293ebb;
    11'b00111011110: data <= 32'hba823d4c;
    11'b00111011111: data <= 32'hbf7db44a;
    11'b00111100000: data <= 32'hbd60bd01;
    11'b00111100001: data <= 32'h3649b406;
    11'b00111100010: data <= 32'h3e183db2;
    11'b00111100011: data <= 32'h3de53e37;
    11'b00111100100: data <= 32'h3cc23435;
    11'b00111100101: data <= 32'h3c4ab474;
    11'b00111100110: data <= 32'h3712398c;
    11'b00111100111: data <= 32'hb9523d4a;
    11'b00111101000: data <= 32'hbb1528b9;
    11'b00111101001: data <= 32'h35c2bfec;
    11'b00111101010: data <= 32'h3e10c107;
    11'b00111101011: data <= 32'h3bcabd8f;
    11'b00111101100: data <= 32'hb6feb446;
    11'b00111101101: data <= 32'hb95a280e;
    11'b00111101110: data <= 32'h34ee3345;
    11'b00111101111: data <= 32'h36423950;
    11'b00111110000: data <= 32'hbd39381b;
    11'b00111110001: data <= 32'hc1aeb7c4;
    11'b00111110010: data <= 32'hc054bc1e;
    11'b00111110011: data <= 32'ha97eb0e4;
    11'b00111110100: data <= 32'h3cbc3c25;
    11'b00111110101: data <= 32'h3ad63b96;
    11'b00111110110: data <= 32'h351e2f34;
    11'b00111110111: data <= 32'h367a36a6;
    11'b00111111000: data <= 32'h36283fb4;
    11'b00111111001: data <= 32'hb23e40ce;
    11'b00111111010: data <= 32'hb6923897;
    11'b00111111011: data <= 32'h3676bf15;
    11'b00111111100: data <= 32'h3d00c05c;
    11'b00111111101: data <= 32'h3be8ba9b;
    11'b00111111110: data <= 32'h34f53090;
    11'b00111111111: data <= 32'h38fdb0b7;
    11'b01000000000: data <= 32'h3ddcb825;
    11'b01000000001: data <= 32'h3b24b0a2;
    11'b01000000010: data <= 32'hbd6a303a;
    11'b01000000011: data <= 32'hc1dcb73c;
    11'b01000000100: data <= 32'hc00abc5f;
    11'b01000000101: data <= 32'h2c4dba59;
    11'b01000000110: data <= 32'h3a67aeeb;
    11'b01000000111: data <= 32'hadd5ad8d;
    11'b01000001000: data <= 32'hb9bcb362;
    11'b01000001001: data <= 32'hb1623a30;
    11'b01000001010: data <= 32'h35ad40f4;
    11'b01000001011: data <= 32'hb0a3416c;
    11'b01000001100: data <= 32'hba6039f2;
    11'b01000001101: data <= 32'hb70cbd2c;
    11'b01000001110: data <= 32'h37adbccf;
    11'b01000001111: data <= 32'h3b0f3444;
    11'b01000010000: data <= 32'h3bae3a02;
    11'b01000010001: data <= 32'h3e3cb2c1;
    11'b01000010010: data <= 32'h404cbaab;
    11'b01000010011: data <= 32'h3d07b039;
    11'b01000010100: data <= 32'hbb5c38d4;
    11'b01000010101: data <= 32'hc0412483;
    11'b01000010110: data <= 32'hbc53bcdf;
    11'b01000010111: data <= 32'h387dbea2;
    11'b01000011000: data <= 32'h3865bd1c;
    11'b01000011001: data <= 32'hb9f7bbcd;
    11'b01000011010: data <= 32'hbc87b92c;
    11'b01000011011: data <= 32'hacaa3828;
    11'b01000011100: data <= 32'h38b24007;
    11'b01000011101: data <= 32'hb6404036;
    11'b01000011110: data <= 32'hbef137c6;
    11'b01000011111: data <= 32'hbeafbaa7;
    11'b01000100000: data <= 32'hb6b8b3ee;
    11'b01000100001: data <= 32'h38ab3c40;
    11'b01000100010: data <= 32'h3c043bc0;
    11'b01000100011: data <= 32'h3e1ab529;
    11'b01000100100: data <= 32'h3fdbb923;
    11'b01000100101: data <= 32'h3d293985;
    11'b01000100110: data <= 32'hb4933ee5;
    11'b01000100111: data <= 32'hbc013a3d;
    11'b01000101000: data <= 32'habc3bca3;
    11'b01000101001: data <= 32'h3bb1c025;
    11'b01000101010: data <= 32'h36debebe;
    11'b01000101011: data <= 32'hba38bcbb;
    11'b01000101100: data <= 32'hb8f1bb5d;
    11'b01000101101: data <= 32'h3a4bb225;
    11'b01000101110: data <= 32'h3c893b16;
    11'b01000101111: data <= 32'hb8c73c48;
    11'b01000110000: data <= 32'hc1062d49;
    11'b01000110001: data <= 32'hc0eeb8a6;
    11'b01000110010: data <= 32'hbb4c2f1a;
    11'b01000110011: data <= 32'h32ba3bcf;
    11'b01000110100: data <= 32'h35e1377f;
    11'b01000110101: data <= 32'h3885b925;
    11'b01000110110: data <= 32'h3c69b404;
    11'b01000110111: data <= 32'h3c373ed4;
    11'b01000111000: data <= 32'h321a4190;
    11'b01000111001: data <= 32'hb4a23daa;
    11'b01000111010: data <= 32'h3495bade;
    11'b01000111011: data <= 32'h3a96bec4;
    11'b01000111100: data <= 32'h34a2bc31;
    11'b01000111101: data <= 32'hb574b8f2;
    11'b01000111110: data <= 32'h3710bb85;
    11'b01000111111: data <= 32'h3fb1bb71;
    11'b01001000000: data <= 32'h3f16b05e;
    11'b01001000001: data <= 32'hb8013632;
    11'b01001000010: data <= 32'hc10da89b;
    11'b01001000011: data <= 32'hc087b81d;
    11'b01001000100: data <= 32'hb98bb303;
    11'b01001000101: data <= 32'haa112d42;
    11'b01001000110: data <= 32'hb88cb855;
    11'b01001000111: data <= 32'hb94bbc9a;
    11'b01001001000: data <= 32'h3384ad5c;
    11'b01001001001: data <= 32'h3acc404f;
    11'b01001001010: data <= 32'h3576421a;
    11'b01001001011: data <= 32'hb5f53e1b;
    11'b01001001100: data <= 32'hb4a5b76b;
    11'b01001001101: data <= 32'h2dbdb9bb;
    11'b01001001110: data <= 32'h16a432de;
    11'b01001001111: data <= 32'h2d253452;
    11'b01001010000: data <= 32'h3d00ba88;
    11'b01001010001: data <= 32'h412cbd45;
    11'b01001010010: data <= 32'h4042b6a5;
    11'b01001010011: data <= 32'hae7b3899;
    11'b01001010100: data <= 32'hbed735ff;
    11'b01001010101: data <= 32'hbcb3b741;
    11'b01001010110: data <= 32'h2b78ba99;
    11'b01001010111: data <= 32'haefdbb83;
    11'b01001011000: data <= 32'hbd17bdb5;
    11'b01001011001: data <= 32'hbd6cbe74;
    11'b01001011010: data <= 32'h2822b5ac;
    11'b01001011011: data <= 32'h3bf73eaa;
    11'b01001011100: data <= 32'h345a40a3;
    11'b01001011101: data <= 32'hbc213c2b;
    11'b01001011110: data <= 32'hbd66b1d9;
    11'b01001011111: data <= 32'hba8b345e;
    11'b01001100000: data <= 32'hb6483d1a;
    11'b01001100001: data <= 32'h2b023a60;
    11'b01001100010: data <= 32'h3cb3ba81;
    11'b01001100011: data <= 32'h409bbd24;
    11'b01001100100: data <= 32'h3fe92f7f;
    11'b01001100101: data <= 32'h35f43e01;
    11'b01001100110: data <= 32'hb8763c95;
    11'b01001100111: data <= 32'h2e46b42d;
    11'b01001101000: data <= 32'h3a33bc7c;
    11'b01001101001: data <= 32'hada1bd28;
    11'b01001101010: data <= 32'hbdc5be46;
    11'b01001101011: data <= 32'hbc8bbf04;
    11'b01001101100: data <= 32'h3967bb7d;
    11'b01001101101: data <= 32'h3e2c3820;
    11'b01001101110: data <= 32'h33393c30;
    11'b01001101111: data <= 32'hbe973526;
    11'b01001110000: data <= 32'hc023ae20;
    11'b01001110001: data <= 32'hbd193a00;
    11'b01001110010: data <= 32'hb9863df4;
    11'b01001110011: data <= 32'hb7df384c;
    11'b01001110100: data <= 32'h322abc78;
    11'b01001110101: data <= 32'h3ce8bc45;
    11'b01001110110: data <= 32'h3dbc3b86;
    11'b01001110111: data <= 32'h395e40ef;
    11'b01001111000: data <= 32'h340f3f18;
    11'b01001111001: data <= 32'h39fc259e;
    11'b01001111010: data <= 32'h3b3bba44;
    11'b01001111011: data <= 32'hb204b900;
    11'b01001111100: data <= 32'hbcbbba8c;
    11'b01001111101: data <= 32'hb4c0bdf5;
    11'b01001111110: data <= 32'h3ed0bdf9;
    11'b01001111111: data <= 32'h4062b8b9;
    11'b01010000000: data <= 32'h35b22b99;
    11'b01010000001: data <= 32'hbea2add6;
    11'b01010000010: data <= 32'hbf59ae3e;
    11'b01010000011: data <= 32'hbb3a38c0;
    11'b01010000100: data <= 32'hb99c3ab4;
    11'b01010000101: data <= 32'hbd07b585;
    11'b01010000110: data <= 32'hbc6cbe99;
    11'b01010000111: data <= 32'h2b86bbd3;
    11'b01010001000: data <= 32'h3b4d3d61;
    11'b01010001001: data <= 32'h39c54167;
    11'b01010001010: data <= 32'h35623f12;
    11'b01010001011: data <= 32'h36fd32f3;
    11'b01010001100: data <= 32'h35322952;
    11'b01010001101: data <= 32'hb806399a;
    11'b01010001110: data <= 32'hbb0235c3;
    11'b01010001111: data <= 32'h36e3bc25;
    11'b01010010000: data <= 32'h40a7bf02;
    11'b01010010001: data <= 32'h40f2bc17;
    11'b01010010010: data <= 32'h38dba901;
    11'b01010010011: data <= 32'hbbb8303c;
    11'b01010010100: data <= 32'hb984a4b8;
    11'b01010010101: data <= 32'h2fc23022;
    11'b01010010110: data <= 32'hb6f1ac42;
    11'b01010010111: data <= 32'hbf41bcc0;
    11'b01010011000: data <= 32'hbfc2c025;
    11'b01010011001: data <= 32'hb726bc9e;
    11'b01010011010: data <= 32'h3aad3b8f;
    11'b01010011011: data <= 32'h39333faa;
    11'b01010011100: data <= 32'hb1503c23;
    11'b01010011101: data <= 32'hb78c31ca;
    11'b01010011110: data <= 32'hb83d3b01;
    11'b01010011111: data <= 32'hbb243f91;
    11'b01010100000: data <= 32'hbae53cd0;
    11'b01010100001: data <= 32'h369aba31;
    11'b01010100010: data <= 32'h4000bec3;
    11'b01010100011: data <= 32'h4035b93c;
    11'b01010100100: data <= 32'h3a4d39a3;
    11'b01010100101: data <= 32'h28253aa9;
    11'b01010100110: data <= 32'h39a9322b;
    11'b01010100111: data <= 32'h3ca8b106;
    11'b01010101000: data <= 32'hafe2b70d;
    11'b01010101001: data <= 32'hbfb4bd2e;
    11'b01010101010: data <= 32'hbf8cc014;
    11'b01010101011: data <= 32'ha465bdea;
    11'b01010101100: data <= 32'h3d24ab85;
    11'b01010101101: data <= 32'h39103838;
    11'b01010101110: data <= 32'hb9d4a41e;
    11'b01010101111: data <= 32'hbcbaa9cc;
    11'b01010110000: data <= 32'hbbb43d15;
    11'b01010110001: data <= 32'hbc3f408c;
    11'b01010110010: data <= 32'hbcc83cc0;
    11'b01010110011: data <= 32'hb6fcbb98;
    11'b01010110100: data <= 32'h3a8dbe00;
    11'b01010110101: data <= 32'h3cf12d65;
    11'b01010110110: data <= 32'h3a123e83;
    11'b01010110111: data <= 32'h39f13dc4;
    11'b01010111000: data <= 32'h3e1d3649;
    11'b01010111001: data <= 32'h3e4624c5;
    11'b01010111010: data <= 32'hab572ef2;
    11'b01010111011: data <= 32'hbebdb748;
    11'b01010111100: data <= 32'hbca0bde0;
    11'b01010111101: data <= 32'h3b7ebed2;
    11'b01010111110: data <= 32'h3fa8bc32;
    11'b01010111111: data <= 32'h39c1b90f;
    11'b01011000000: data <= 32'hbad0b9e2;
    11'b01011000001: data <= 32'hbc2bb40c;
    11'b01011000010: data <= 32'hb8283c78;
    11'b01011000011: data <= 32'hba653f02;
    11'b01011000100: data <= 32'hbe923697;
    11'b01011000101: data <= 32'hbe72bdd0;
    11'b01011000110: data <= 32'hb829bd96;
    11'b01011000111: data <= 32'h3621386f;
    11'b01011001000: data <= 32'h38813fbb;
    11'b01011001001: data <= 32'h3a783d87;
    11'b01011001010: data <= 32'h3d7635ab;
    11'b01011001011: data <= 32'h3c88386c;
    11'b01011001100: data <= 32'hb53c3d3d;
    11'b01011001101: data <= 32'hbd8a3b1b;
    11'b01011001110: data <= 32'hb675b959;
    11'b01011001111: data <= 32'h3e71bebd;
    11'b01011010000: data <= 32'h4052bdc6;
    11'b01011010001: data <= 32'h3a3fbb2b;
    11'b01011010010: data <= 32'hb6a4b995;
    11'b01011010011: data <= 32'ha2e8b3e6;
    11'b01011010100: data <= 32'h39483960;
    11'b01011010101: data <= 32'hb1cb3add;
    11'b01011010110: data <= 32'hbf96b755;
    11'b01011010111: data <= 32'hc0c7bf71;
    11'b01011011000: data <= 32'hbcd2bdb7;
    11'b01011011001: data <= 32'h2cc535fc;
    11'b01011011010: data <= 32'h36193d0a;
    11'b01011011011: data <= 32'h353d3812;
    11'b01011011100: data <= 32'h3802a5f6;
    11'b01011011101: data <= 32'h346d3c4b;
    11'b01011011110: data <= 32'hb9b340dd;
    11'b01011011111: data <= 32'hbd133fb1;
    11'b01011100000: data <= 32'hb3b4b048;
    11'b01011100001: data <= 32'h3d8ebde1;
    11'b01011100010: data <= 32'h3eb1bc5c;
    11'b01011100011: data <= 32'h391fb353;
    11'b01011100100: data <= 32'h3455a794;
    11'b01011100101: data <= 32'h3d3aa8ce;
    11'b01011100110: data <= 32'h3f9e352b;
    11'b01011100111: data <= 32'h37013579;
    11'b01011101000: data <= 32'hbf43b956;
    11'b01011101001: data <= 32'hc0aebeef;
    11'b01011101010: data <= 32'hbb0dbdda;
    11'b01011101011: data <= 32'h373fb542;
    11'b01011101100: data <= 32'h35a0aa37;
    11'b01011101101: data <= 32'hb44ab9fd;
    11'b01011101110: data <= 32'hb4fcb8af;
    11'b01011101111: data <= 32'hb3f83cf6;
    11'b01011110000: data <= 32'hba90419c;
    11'b01011110001: data <= 32'hbd694015;
    11'b01011110010: data <= 32'hba75b221;
    11'b01011110011: data <= 32'h34b1bcfb;
    11'b01011110100: data <= 32'h38cdb564;
    11'b01011110101: data <= 32'h341b3a16;
    11'b01011110110: data <= 32'h39ce3944;
    11'b01011110111: data <= 32'h403a301e;
    11'b01011111000: data <= 32'h40f134b1;
    11'b01011111001: data <= 32'h395a3910;
    11'b01011111010: data <= 32'hbe092d34;
    11'b01011111011: data <= 32'hbe6cbbca;
    11'b01011111100: data <= 32'h2ea3bd52;
    11'b01011111101: data <= 32'h3c91bc2c;
    11'b01011111110: data <= 32'h36c8bcc0;
    11'b01011111111: data <= 32'hb86dbea2;
    11'b01100000000: data <= 32'hb66fbc08;
    11'b01100000001: data <= 32'h2e273be7;
    11'b01100000010: data <= 32'hb6434092;
    11'b01100000011: data <= 32'hbdcd3d12;
    11'b01100000100: data <= 32'hbec7b9d5;
    11'b01100000101: data <= 32'hbc13bc8d;
    11'b01100000110: data <= 32'hb77d3421;
    11'b01100000111: data <= 32'hb2783d11;
    11'b01100001000: data <= 32'h393f399f;
    11'b01100001001: data <= 32'h3fd3a9e5;
    11'b01100001010: data <= 32'h40273801;
    11'b01100001011: data <= 32'h36633e2f;
    11'b01100001100: data <= 32'hbcd23d90;
    11'b01100001101: data <= 32'hba102b58;
    11'b01100001110: data <= 32'h3b9bbc04;
    11'b01100001111: data <= 32'h3dfbbd10;
    11'b01100010000: data <= 32'h3619bdd9;
    11'b01100010001: data <= 32'hb697bed0;
    11'b01100010010: data <= 32'h3589bc2f;
    11'b01100010011: data <= 32'h3cee383b;
    11'b01100010100: data <= 32'h37613d4b;
    11'b01100010101: data <= 32'hbd7b340b;
    11'b01100010110: data <= 32'hc08abcfa;
    11'b01100010111: data <= 32'hbedebc63;
    11'b01100011000: data <= 32'hbb38356a;
    11'b01100011001: data <= 32'hb7ac3ae6;
    11'b01100011010: data <= 32'h308baf78;
    11'b01100011011: data <= 32'h3c2eb934;
    11'b01100011100: data <= 32'h3c6c3963;
    11'b01100011101: data <= 32'hadb040e3;
    11'b01100011110: data <= 32'hbc2d40e0;
    11'b01100011111: data <= 32'hb5e43a11;
    11'b01100100000: data <= 32'h3be4b91c;
    11'b01100100001: data <= 32'h3c4cbad2;
    11'b01100100010: data <= 32'h27c0ba1f;
    11'b01100100011: data <= 32'hacd2bbae;
    11'b01100100100: data <= 32'h3db5b9ff;
    11'b01100100101: data <= 32'h40fb30f9;
    11'b01100100110: data <= 32'h3d1f38ea;
    11'b01100100111: data <= 32'hbc58b270;
    11'b01100101000: data <= 32'hc042bccf;
    11'b01100101001: data <= 32'hbd84bb8f;
    11'b01100101010: data <= 32'hb7e1a5d7;
    11'b01100101011: data <= 32'hb738b251;
    11'b01100101100: data <= 32'hb77cbd8c;
    11'b01100101101: data <= 32'h2c83bdc3;
    11'b01100101110: data <= 32'h359a38bc;
    11'b01100101111: data <= 32'hb4cb4165;
    11'b01100110000: data <= 32'hbbcb411d;
    11'b01100110001: data <= 32'hb8de39bc;
    11'b01100110010: data <= 32'h30a9b6e9;
    11'b01100110011: data <= 32'h9d8bad68;
    11'b01100110100: data <= 32'hb8c935b7;
    11'b01100110101: data <= 32'h2e04abfb;
    11'b01100110110: data <= 32'h402db77a;
    11'b01100110111: data <= 32'h42251ec4;
    11'b01100111000: data <= 32'h3e4f38d0;
    11'b01100111001: data <= 32'hba003498;
    11'b01100111010: data <= 32'hbd7ab72e;
    11'b01100111011: data <= 32'hb493b87e;
    11'b01100111100: data <= 32'h3611b6ce;
    11'b01100111101: data <= 32'hb423bcb1;
    11'b01100111110: data <= 32'hbab9c0a8;
    11'b01100111111: data <= 32'hb4c2bfeb;
    11'b01101000000: data <= 32'h36e93423;
    11'b01101000001: data <= 32'h2e854045;
    11'b01101000010: data <= 32'hbaa43ecc;
    11'b01101000011: data <= 32'hbcac2777;
    11'b01101000100: data <= 32'hbbe1b6ff;
    11'b01101000101: data <= 32'hbc793899;
    11'b01101000110: data <= 32'hbce23c74;
    11'b01101000111: data <= 32'haee133dc;
    11'b01101001000: data <= 32'h3f7db8b6;
    11'b01101001001: data <= 32'h413da000;
    11'b01101001010: data <= 32'h3cca3cba;
    11'b01101001011: data <= 32'hb8533d97;
    11'b01101001100: data <= 32'hb78b3910;
    11'b01101001101: data <= 32'h3a4ea7f2;
    11'b01101001110: data <= 32'h3bf3b777;
    11'b01101001111: data <= 32'hb32dbd7b;
    11'b01101010000: data <= 32'hbb26c0b0;
    11'b01101010001: data <= 32'h2fc7bfd2;
    11'b01101010010: data <= 32'h3d6bb04a;
    11'b01101010011: data <= 32'h3c013c84;
    11'b01101010100: data <= 32'hb82137af;
    11'b01101010101: data <= 32'hbe13b9eb;
    11'b01101010110: data <= 32'hbe5bb7e6;
    11'b01101010111: data <= 32'hbe363a93;
    11'b01101011000: data <= 32'hbdf83c1e;
    11'b01101011001: data <= 32'hb8beb58e;
    11'b01101011010: data <= 32'h3b5dbcea;
    11'b01101011011: data <= 32'h3de1ad4c;
    11'b01101011100: data <= 32'h37803f47;
    11'b01101011101: data <= 32'hb7de40ac;
    11'b01101011110: data <= 32'h2b783d73;
    11'b01101011111: data <= 32'h3c883634;
    11'b01101100000: data <= 32'h3a82a896;
    11'b01101100001: data <= 32'hb8bbb90c;
    11'b01101100010: data <= 32'hba73bdcd;
    11'b01101100011: data <= 32'h3b5ebdc4;
    11'b01101100100: data <= 32'h40f9b63a;
    11'b01101100101: data <= 32'h3f7d34da;
    11'b01101100110: data <= 32'hafe7b45d;
    11'b01101100111: data <= 32'hbd3fbba1;
    11'b01101101000: data <= 32'hbccfb599;
    11'b01101101001: data <= 32'hbc1d399d;
    11'b01101101010: data <= 32'hbd223440;
    11'b01101101011: data <= 32'hbc5cbde9;
    11'b01101101100: data <= 32'hb0d9c02b;
    11'b01101101101: data <= 32'h36d8b51d;
    11'b01101101110: data <= 32'ha21f3fd8;
    11'b01101101111: data <= 32'hb75440cb;
    11'b01101110000: data <= 32'h29cd3cf8;
    11'b01101110001: data <= 32'h38cb3763;
    11'b01101110010: data <= 32'haf1a391e;
    11'b01101110011: data <= 32'hbd2d3899;
    11'b01101110100: data <= 32'hbaa3b48e;
    11'b01101110101: data <= 32'h3db8bb0c;
    11'b01101110110: data <= 32'h4204b791;
    11'b01101110111: data <= 32'h40412d3f;
    11'b01101111000: data <= 32'h304bae64;
    11'b01101111001: data <= 32'hb8e9b609;
    11'b01101111010: data <= 32'ha8742eae;
    11'b01101111011: data <= 32'h2db33827;
    11'b01101111100: data <= 32'hba87b82e;
    11'b01101111101: data <= 32'hbd80c0b5;
    11'b01101111110: data <= 32'hb9a6c13e;
    11'b01101111111: data <= 32'h3207b90d;
    11'b01110000000: data <= 32'h31f63db4;
    11'b01110000001: data <= 32'hb41d3de2;
    11'b01110000010: data <= 32'hb4723564;
    11'b01110000011: data <= 32'hb50a3248;
    11'b01110000100: data <= 32'hbc9b3ccb;
    11'b01110000101: data <= 32'hbfcd3dfe;
    11'b01110000110: data <= 32'hbc44358a;
    11'b01110000111: data <= 32'h3cd1ba2e;
    11'b01110001000: data <= 32'h40fab828;
    11'b01110001001: data <= 32'h3e4136bb;
    11'b01110001010: data <= 32'h2f0b3a25;
    11'b01110001011: data <= 32'h31d738f9;
    11'b01110001100: data <= 32'h3cc33996;
    11'b01110001101: data <= 32'h3c193888;
    11'b01110001110: data <= 32'hb837b965;
    11'b01110001111: data <= 32'hbdbac0a0;
    11'b01110010000: data <= 32'hb832c0e8;
    11'b01110010001: data <= 32'h3ac5ba9f;
    11'b01110010010: data <= 32'h3be1381b;
    11'b01110010011: data <= 32'h30682f34;
    11'b01110010100: data <= 32'hb7e1b9fd;
    11'b01110010101: data <= 32'hbab3b03b;
    11'b01110010110: data <= 32'hbe283daf;
    11'b01110010111: data <= 32'hc0403e92;
    11'b01110011000: data <= 32'hbd9c28df;
    11'b01110011001: data <= 32'h3544bd26;
    11'b01110011010: data <= 32'h3cdab970;
    11'b01110011011: data <= 32'h383c3b19;
    11'b01110011100: data <= 32'hafe23e5d;
    11'b01110011101: data <= 32'h39543d3e;
    11'b01110011110: data <= 32'h3f063c47;
    11'b01110011111: data <= 32'h3c973b38;
    11'b01110100000: data <= 32'hb9ee20b1;
    11'b01110100001: data <= 32'hbdb0bd3a;
    11'b01110100010: data <= 32'h2d0abe9e;
    11'b01110100011: data <= 32'h3f54ba68;
    11'b01110100100: data <= 32'h3f44b402;
    11'b01110100101: data <= 32'h3839bad3;
    11'b01110100110: data <= 32'hb52fbd22;
    11'b01110100111: data <= 32'hb7b0b187;
    11'b01110101000: data <= 32'hbb5b3d75;
    11'b01110101001: data <= 32'hbea83c5c;
    11'b01110101010: data <= 32'hbe86bb59;
    11'b01110101011: data <= 32'hb95cc033;
    11'b01110101100: data <= 32'ha848bb9b;
    11'b01110101101: data <= 32'hb49d3c0d;
    11'b01110101110: data <= 32'hb4e73e9e;
    11'b01110101111: data <= 32'h39923c75;
    11'b01110110000: data <= 32'h3dc73b79;
    11'b01110110001: data <= 32'h36cc3d59;
    11'b01110110010: data <= 32'hbd903c8f;
    11'b01110110011: data <= 32'hbe062ae8;
    11'b01110110100: data <= 32'h3834b9fa;
    11'b01110110101: data <= 32'h40a8b919;
    11'b01110110110: data <= 32'h4007b7e1;
    11'b01110110111: data <= 32'h3900bb4b;
    11'b01110111000: data <= 32'h3189bb82;
    11'b01110111001: data <= 32'h38f232bb;
    11'b01110111010: data <= 32'h360e3d08;
    11'b01110111011: data <= 32'hbace3670;
    11'b01110111100: data <= 32'hbe96befb;
    11'b01110111101: data <= 32'hbce4c131;
    11'b01110111110: data <= 32'hb815bc9b;
    11'b01110111111: data <= 32'hb5ae3911;
    11'b01111000000: data <= 32'hb28b3a47;
    11'b01111000001: data <= 32'h374b29b3;
    11'b01111000010: data <= 32'h394f3564;
    11'b01111000011: data <= 32'hb8593e78;
    11'b01111000100: data <= 32'hc00b4016;
    11'b01111000101: data <= 32'hbeb93b68;
    11'b01111000110: data <= 32'h3689b574;
    11'b01111000111: data <= 32'h3f6ab865;
    11'b01111001000: data <= 32'h3d39b371;
    11'b01111001001: data <= 32'h34b3b297;
    11'b01111001010: data <= 32'h3990a907;
    11'b01111001011: data <= 32'h3f403a4e;
    11'b01111001100: data <= 32'h3e393d28;
    11'b01111001101: data <= 32'hb38a3208;
    11'b01111001110: data <= 32'hbe1fbef1;
    11'b01111001111: data <= 32'hbc6ec09e;
    11'b01111010000: data <= 32'ha90bbc4d;
    11'b01111010001: data <= 32'h34faa599;
    11'b01111010010: data <= 32'h3184b84f;
    11'b01111010011: data <= 32'h3432bd20;
    11'b01111010100: data <= 32'h2fe4b56c;
    11'b01111010101: data <= 32'hbb9c3e8a;
    11'b01111010110: data <= 32'hc037407a;
    11'b01111010111: data <= 32'hbf273a9a;
    11'b01111011000: data <= 32'hb375b97c;
    11'b01111011001: data <= 32'h38e8b96b;
    11'b01111011010: data <= 32'h28c331f8;
    11'b01111011011: data <= 32'hb4c738be;
    11'b01111011100: data <= 32'h3b94393f;
    11'b01111011101: data <= 32'h40d43c67;
    11'b01111011110: data <= 32'h3f9e3dc9;
    11'b01111011111: data <= 32'hb3b0395b;
    11'b01111100000: data <= 32'hbddbba23;
    11'b01111100001: data <= 32'hb887bd28;
    11'b01111100010: data <= 32'h3b16b982;
    11'b01111100011: data <= 32'h3c85b84b;
    11'b01111100100: data <= 32'h383dbe20;
    11'b01111100101: data <= 32'h34e0c01f;
    11'b01111100110: data <= 32'h3507b908;
    11'b01111100111: data <= 32'hb5eb3df6;
    11'b01111101000: data <= 32'hbdca3f04;
    11'b01111101001: data <= 32'hbeaca8cb;
    11'b01111101010: data <= 32'hbbcdbdda;
    11'b01111101011: data <= 32'hb939bb76;
    11'b01111101100: data <= 32'hbc2b363e;
    11'b01111101101: data <= 32'hba2b3a44;
    11'b01111101110: data <= 32'h3adc37fb;
    11'b01111101111: data <= 32'h40583a62;
    11'b01111110000: data <= 32'h3d3b3e3d;
    11'b01111110001: data <= 32'hba9b3e2f;
    11'b01111110010: data <= 32'hbe2738d8;
    11'b01111110011: data <= 32'had26aee3;
    11'b01111110100: data <= 32'h3de1b264;
    11'b01111110101: data <= 32'h3d78b900;
    11'b01111110110: data <= 32'h37eabea1;
    11'b01111110111: data <= 32'h3826bf7f;
    11'b01111111000: data <= 32'h3cafb585;
    11'b01111111001: data <= 32'h3b773d7c;
    11'b01111111010: data <= 32'hb5b93c3b;
    11'b01111111011: data <= 32'hbd54bb5a;
    11'b01111111100: data <= 32'hbd60bffb;
    11'b01111111101: data <= 32'hbcc9bc25;
    11'b01111111110: data <= 32'hbd3633ff;
    11'b01111111111: data <= 32'hba7d3056;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    