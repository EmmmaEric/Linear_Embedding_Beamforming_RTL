
    module interp_rom_1(
    CLK, rst,
    Addr, CEB, Q
    );

    input CLK, rst;
    input [9:0] Addr;
    input CEB;		
    output [20:0] Q;

    (*rom_style = "block" *) reg [20:0] data;

    always @(posedge CLK) begin
    if (rst) begin
        data <= 20'd0;
    end else begin
    if (CEB)
    case(Addr)
            10'b00000000: data <= 20'b10111101000101001000;
        10'b00000001: data <= 20'b11001000011100101111;
        10'b00000010: data <= 20'b01001000101100100101;
        10'b00000011: data <= 20'b10111010101100111110;
        10'b00000100: data <= 20'b10111001101100100010;
        10'b00000101: data <= 20'b01001011011100100011;
        10'b00000110: data <= 20'b11001000001100101011;
        10'b00000111: data <= 20'b00110111100100000101;
        10'b00001000: data <= 20'b11010010100101000001;
        10'b00001001: data <= 20'b00111110011100100010;
        10'b00001010: data <= 20'b01010000101100101010;
        10'b00001011: data <= 20'b11000111001100110010;
        10'b00001100: data <= 20'b01000111001100100101;
        10'b00001101: data <= 20'b00111010011100111110;
        10'b00001110: data <= 20'b11000011111100011011;
        10'b00001111: data <= 20'b01000110010100001010;
        10'b00010000: data <= 20'b11001100001100110111;
        10'b00010001: data <= 20'b01000110010100000001;
        10'b00010010: data <= 20'b11010110111101011001;
        10'b00010011: data <= 20'b00111011101100101010;
        10'b00010100: data <= 20'b01001100111100110111;
        10'b00010101: data <= 20'b11000111101100101111;
        10'b00010110: data <= 20'b00111101111100010101;
        10'b00010111: data <= 20'b01001111101100101000;
        10'b00011000: data <= 20'b11000110001100100000;
        10'b00011001: data <= 20'b01000011110100010110;
        10'b00011010: data <= 20'b11001110011101000001;
        10'b00011011: data <= 20'b01001011001100100001;
        10'b00011100: data <= 20'b11000110111101000110;
        10'b00011101: data <= 20'b11000000101100100111;
        10'b00011110: data <= 20'b01001010101100100000;
        10'b00011111: data <= 20'b11001001001100110111;
        10'b00100000: data <= 20'b11000000101100010100;
        10'b00100001: data <= 20'b01001001010100010011;
        10'b00100010: data <= 20'b00100000101100100100;
        10'b00100011: data <= 20'b01001110010100100111;
        10'b00100100: data <= 20'b11001001111100110111;
        10'b00100101: data <= 20'b01000111011100011110;
        10'b00100110: data <= 20'b01001001101101001101;
        10'b00100111: data <= 20'b11000110001100100111;
        10'b00101000: data <= 20'b01000100011100010000;
        10'b00101001: data <= 20'b01001000011101000000;
        10'b00101010: data <= 20'b10110111001100001100;
        10'b00101011: data <= 20'b01001100100100110011;
        10'b00101100: data <= 20'b00111100001100101000;
        10'b00101101: data <= 20'b01010000101011010111;
        10'b00101110: data <= 20'b11001011111100110110;
        10'b00101111: data <= 20'b10110101101100100000;
        10'b00110000: data <= 20'b01001100011100100110;
        10'b00110001: data <= 20'b11000110001100101111;
        10'b00110010: data <= 20'b01000001001100001101;
        10'b00110011: data <= 20'b01001101111100110001;
        10'b00110100: data <= 20'b01000100110011111000;
        10'b00110101: data <= 20'b11010100000101100010;
        10'b00110110: data <= 20'b11000110101100101001;
        10'b00110111: data <= 20'b01001001101100011001;
        10'b00111000: data <= 20'b11000111101101000011;
        10'b00111001: data <= 20'b11000001011100100100;
        10'b00111010: data <= 20'b01001000001100011111;
        10'b00111011: data <= 20'b11000011111100101010;
        10'b00111100: data <= 20'b01000010110100010011;
        10'b00111101: data <= 20'b11010011001100110100;
        10'b00111110: data <= 20'b01000010111100010110;
        10'b00111111: data <= 20'b01010100010100100100;
        10'b01000000: data <= 20'b11001001001100110000;
        10'b01000001: data <= 20'b01000010111100100010;
        10'b01000010: data <= 20'b01000111101100110111;
        10'b01000011: data <= 20'b11000000101100100000;
        10'b01000100: data <= 20'b01001001000011101111;
        10'b01000101: data <= 20'b11001000111100101110;
        10'b01000110: data <= 20'b01000101000100011110;
        10'b01000111: data <= 20'b11010011011100101111;
        10'b01001000: data <= 20'b11000000111100100111;
        10'b01001001: data <= 20'b01001011111100100111;
        10'b01001010: data <= 20'b11000101111100110100;
        10'b01001011: data <= 20'b01000000111100011111;
        10'b01001100: data <= 20'b01001011111100110111;
        10'b01001101: data <= 20'b11000100111100010100;
        10'b01001110: data <= 20'b01000000100100101000;
        10'b01001111: data <= 20'b11001100111100101111;
        10'b01010000: data <= 20'b01001000001100010111;
        10'b01010001: data <= 20'b01001011101101001100;
        10'b01010010: data <= 20'b11000001001100101011;
        10'b01010011: data <= 20'b01001001001100101001;
        10'b01010100: data <= 20'b11000110011100110010;
        10'b01010101: data <= 20'b10111010101100000110;
        10'b01010110: data <= 20'b01001100010100110010;
        10'b01010111: data <= 20'b11000011101100011101;
        10'b01011000: data <= 20'b01001010110100101011;
        10'b01011001: data <= 20'b11001100101100111001;
        10'b01011010: data <= 20'b01000100111100101000;
        10'b01011011: data <= 20'b01000111011101000000;
        10'b01011100: data <= 20'b11000100011100100101;
        10'b01011101: data <= 20'b01000111011100001011;
        10'b01011110: data <= 20'b11000110011101000001;
        10'b01011111: data <= 20'b11000000011100000000;
        10'b01100000: data <= 20'b01000010100100110110;
        10'b01100001: data <= 20'b11000100111100110000;
        10'b01100010: data <= 20'b01001101101100101000;
        10'b01100011: data <= 20'b11001000001100111000;
        10'b01100100: data <= 20'b00111111001100100001;
        10'b01100101: data <= 20'b01001101111100110100;
        10'b01100110: data <= 20'b11000111111100101000;
        10'b01100111: data <= 20'b00111011101011110101;
        10'b01101000: data <= 20'b01010001010101000000;
        10'b01101001: data <= 20'b01000101001100001101;
        10'b01101010: data <= 20'b01010111000100101101;
        10'b01101011: data <= 20'b11000001001100101110;
        10'b01101100: data <= 20'b01001011101100100101;
        10'b01101101: data <= 20'b11001010001100111100;
        10'b01101110: data <= 20'b11000001101100100000;
        10'b01101111: data <= 20'b01001000111100000101;
        10'b01110000: data <= 20'b11000111011100110011;
        10'b01110001: data <= 20'b01000001010011110001;
        10'b01110010: data <= 20'b11011001000101110001;
        10'b01110011: data <= 20'b01001000001100100010;
        10'b01110100: data <= 20'b01010000111101001101;
        10'b01110101: data <= 20'b11000111111100101100;
        10'b01110110: data <= 20'b01000100101100011000;
        10'b01110111: data <= 20'b01001100001101000010;
        10'b01111000: data <= 20'b11000100011100100001;
        10'b01111001: data <= 20'b01000101110010101110;
        10'b01111010: data <= 20'b01000000101100110101;
        10'b01111011: data <= 20'b01001100010100011111;
        10'b01111100: data <= 20'b11001110111101000010;
        10'b01111101: data <= 20'b10110010011100100011;
        10'b01111110: data <= 20'b01001101111100100100;
        10'b01111111: data <= 20'b11001001011100110011;
        10'b10000000: data <= 20'b00101000001100011101;
        10'b10000001: data <= 20'b01001010111100100011;
        10'b10000010: data <= 20'b10111110001100010111;
        10'b10000011: data <= 20'b01001010000100101101;
        10'b10000100: data <= 20'b11001001011100110010;
        10'b10000101: data <= 20'b01001001111011111001;
        10'b10000110: data <= 20'b11010000101101010000;
        10'b10000111: data <= 20'b11000101001100101000;
        10'b10001000: data <= 20'b01000111101100100000;
        10'b10001001: data <= 20'b10111110101100110111;
        10'b10001010: data <= 20'b00110111101100010100;
        10'b10001011: data <= 20'b01001101100011110001;
        10'b10001100: data <= 20'b10111100101100010011;
        10'b10001101: data <= 20'b01001011110100111010;
        10'b10001110: data <= 20'b11001100011100110010;
        10'b10001111: data <= 20'b01000001111100100001;
        10'b10010000: data <= 20'b01001101001100111001;
        10'b10010001: data <= 20'b11000100111100101010;
        10'b10010010: data <= 20'b01000110001100011101;
        10'b10010011: data <= 20'b10111100101100110110;
        10'b10010100: data <= 20'b10111011000011010110;
        10'b10010101: data <= 20'b11001000000101000100;
        10'b10010110: data <= 20'b11000100101100100110;
        10'b10010111: data <= 20'b01001100011100001001;
        10'b10011000: data <= 20'b11001010001101000000;
        10'b10011001: data <= 20'b00110000101100100101;
        10'b10011010: data <= 20'b01001001111100110010;
        10'b10011011: data <= 20'b11000101101100100110;
        10'b10011100: data <= 20'b01000010100011101011;
        10'b10011101: data <= 20'b11010101001101011011;
        10'b10011110: data <= 20'b01000000101011110011;
        10'b10011111: data <= 20'b01001111000101010001;
        10'b10100000: data <= 20'b11000111001100101111;
        10'b10100001: data <= 20'b01001000101100101000;
        10'b10100010: data <= 20'b11000010001100111010;
        10'b10100011: data <= 20'b10111100111100011110;
        10'b10100100: data <= 20'b01001100001100010010;
        10'b10100101: data <= 20'b11001000111100101011;
        10'b10100110: data <= 20'b00110100100100010000;
        10'b10100111: data <= 20'b11010010000100110001;
        10'b10101000: data <= 20'b01000000111100100110;
        10'b10101001: data <= 20'b01001110111100111001;
        10'b10101010: data <= 20'b11000101001100110000;
        10'b10101011: data <= 20'b01000110101100100001;
        10'b10101100: data <= 20'b00111101011101000001;
        10'b10101101: data <= 20'b11000100101100011010;
        10'b10101110: data <= 20'b01000011000100010010;
        10'b10101111: data <= 20'b11001101011100110100;
        10'b10110000: data <= 20'b01001001111010000110;
        10'b10110001: data <= 20'b11001101101101010001;
        10'b10110010: data <= 20'b00111110011100101000;
        10'b10110011: data <= 20'b01001101001100110110;
        10'b10110100: data <= 20'b11001000011100110000;
        10'b10110101: data <= 20'b00111001101100010010;
        10'b10110110: data <= 20'b01001110101100001001;
        10'b10110111: data <= 20'b11000101001100011101;
        10'b10111000: data <= 20'b01000111000100100001;
        10'b10111001: data <= 20'b11001010111100111101;
        10'b10111010: data <= 20'b01001011111100100011;
        10'b10111011: data <= 20'b11001001001101000011;
        10'b10111100: data <= 20'b11000010101100100100;
        10'b10111101: data <= 20'b01001001111100010111;
        10'b10111110: data <= 20'b11001000111100111001;
        10'b10111111: data <= 20'b10111111101100010010;
        10'b11000000: data <= 20'b01001001010100011101;
        10'b11000001: data <= 20'b01000000111100100011;
        10'b11000010: data <= 20'b01010001010100100111;
        10'b11000011: data <= 20'b11001001011100110011;
        10'b11000100: data <= 20'b01000101111100011110;
        10'b11000101: data <= 20'b01001101111101000101;
        10'b11000110: data <= 20'b11000111011100101001;
        10'b11000111: data <= 20'b01000010001100010010;
        10'b11001000: data <= 20'b01001011011100111000;
        10'b11001001: data <= 20'b01000000101011110111;
        10'b11001010: data <= 20'b01010001010101001010;
        10'b11001011: data <= 20'b10111000101100100101;
        10'b11001100: data <= 20'b01001111101100000010;
        10'b11001101: data <= 20'b11001011111100111000;
        10'b11001110: data <= 20'b10111100001100100001;
        10'b11001111: data <= 20'b01001010111100100100;
        10'b11010000: data <= 20'b11000101001100101100;
        10'b11010001: data <= 20'b01000011011011111011;
        10'b11010010: data <= 20'b01010000001101000110;
        10'b11010011: data <= 20'b01000110000100000010;
        10'b11010100: data <= 20'b11011000100101010010;
        10'b11010101: data <= 20'b11000110101100101001;
        10'b11010110: data <= 20'b01001000011100011111;
        10'b11010111: data <= 20'b00111100111101000010;
        10'b11011000: data <= 20'b11000000101100100010;
        10'b11011001: data <= 20'b01001001001100011101;
        10'b11011010: data <= 20'b11000101011100100111;
        10'b11011011: data <= 20'b01000001100100100000;
        10'b11011100: data <= 20'b11010001011100101010;
        10'b11011101: data <= 20'b01000001111100011101;
        10'b11011110: data <= 20'b01010010001100101101;
        10'b11011111: data <= 20'b11001000011100110010;
        10'b11100000: data <= 20'b01000010111100100010;
        10'b11100001: data <= 20'b01000110111100110111;
        10'b11100010: data <= 20'b11000000101100011000;
        10'b11100011: data <= 20'b01001001000100011011;
        10'b11100100: data <= 20'b11001001001100101101;
        10'b11100101: data <= 20'b01001000010100011000;
        10'b11100110: data <= 20'b11010010101101000011;
        10'b11100111: data <= 20'b10111111011100101000;
        10'b11101000: data <= 20'b01001010101100101100;
        10'b11101001: data <= 20'b11000101011100110001;
        10'b11101010: data <= 20'b01000000101100011000;
        10'b11101011: data <= 20'b01001110101100110100;
        10'b11101100: data <= 20'b11000101001100010001;
        10'b11101101: data <= 20'b00111101110100101101;
        10'b11101110: data <= 20'b11001100111100110000;
        10'b11101111: data <= 20'b01001000011100100001;
        10'b11110000: data <= 20'b01000110111101000010;
        10'b11110001: data <= 20'b10111111111100101001;
        10'b11110010: data <= 20'b01001001111100100111;
        10'b11110011: data <= 20'b11000111101100110011;
        10'b11110100: data <= 20'b10111110011100000001;
        10'b11110101: data <= 20'b01001000010100110100;
        10'b11110110: data <= 20'b11000001011100100010;
        10'b11110111: data <= 20'b01001101010100100001;
        10'b11111000: data <= 20'b11001011101100111001;
        10'b11111001: data <= 20'b01000101111100101000;
        10'b11111010: data <= 20'b01000110001100111110;
        10'b11111011: data <= 20'b11000100111100100100;
        10'b11111100: data <= 20'b01000101011100000000;
        10'b11111101: data <= 20'b11000010111101001001;
        10'b11111110: data <= 20'b10111100001011110011;
        10'b11111111: data <= 20'b01000100110101000000;
        10'b100000000: data <= 20'b11000000101100110000;
        10'b100000001: data <= 20'b01001101011100110001;
        10'b100000010: data <= 20'b11001000011100110101;
        10'b100000011: data <= 20'b00111010111100011111;
        10'b100000100: data <= 20'b01001101111100101100;
        10'b100000101: data <= 20'b11001000001100101001;
        10'b100000110: data <= 20'b00111011111011100110;
        10'b100000111: data <= 20'b01010000100101001010;
        10'b100001000: data <= 20'b01001000011100010110;
        10'b100001001: data <= 20'b01010100001101010101;
        10'b100001010: data <= 20'b11000011111100101100;
        10'b100001011: data <= 20'b01001010011100100000;
        10'b100001100: data <= 20'b11001001111101000000;
        10'b100001101: data <= 20'b11000010101100011110;
        10'b100001110: data <= 20'b01000111111011111011;
        10'b100001111: data <= 20'b11000100101100110011;
        10'b100010000: data <= 20'b01000110100100010000;
        10'b100010001: data <= 20'b11010001001101001001;
        10'b100010010: data <= 20'b01000110101100100000;
        10'b100010011: data <= 20'b01010001111101001011;
        10'b100010100: data <= 20'b11001000101100101101;
        10'b100010101: data <= 20'b01000001111100011001;
        10'b100010110: data <= 20'b01001101011100111001;
        10'b100010111: data <= 20'b11000010101100100000;
        10'b100011000: data <= 20'b01000111010011111000;
        10'b100011001: data <= 20'b10111000101100110101;
        10'b100011010: data <= 20'b01001100100100100010;
        10'b100011011: data <= 20'b11001111001100111100;
        10'b100011100: data <= 20'b10111100001100100011;
        10'b100011101: data <= 20'b01001100111100100100;
        10'b100011110: data <= 20'b11001000001100110011;
        10'b100011111: data <= 20'b00110111101100011100;
        10'b100100000: data <= 20'b01001011101100100101;
        10'b100100001: data <= 20'b10111101111100010000;
        10'b100100010: data <= 20'b01001001000100110111;
        10'b100100011: data <= 20'b11001001111100101111;
        10'b100100100: data <= 20'b01001000111100010010;
        10'b100100101: data <= 20'b11000111001101010001;
        10'b100100110: data <= 20'b11000100101100101000;
        10'b100100111: data <= 20'b01000111001100100001;
        10'b100101000: data <= 20'b11000001011100110100;
        10'b100101001: data <= 20'b00111010101100000100;
        10'b100101010: data <= 20'b01010000000100110110;
        10'b100101011: data <= 20'b10110100101100010101;
        10'b100101100: data <= 20'b01001110010100111001;
        10'b100101101: data <= 20'b11001100011100110100;
        10'b100101110: data <= 20'b01000000011100100011;
        10'b100101111: data <= 20'b01001011011100110111;
        10'b100110000: data <= 20'b11000100001100100111;
        10'b100110001: data <= 20'b01000110111100010011;
        10'b100110010: data <= 20'b11000011101100111011;
        10'b100110011: data <= 20'b10111011100011111100;
        10'b100110100: data <= 20'b11001101000101000011;
        10'b100110101: data <= 20'b11000101011100101001;
        10'b100110110: data <= 20'b01001011101100011011;
        10'b100110111: data <= 20'b11001000111100111101;
        10'b100111000: data <= 20'b00111101101100100101;
        10'b100111001: data <= 20'b01001010001100110011;
        10'b100111010: data <= 20'b11000110001100100101;
        10'b100111011: data <= 20'b00111111010100000100;
        10'b100111100: data <= 20'b11010100100100100100;
        10'b100111101: data <= 20'b01000010101100001010;
        10'b100111110: data <= 20'b01010100110101000100;
        10'b100111111: data <= 20'b11000110011100110000;
        10'b101000000: data <= 20'b01001000101100101001;
        10'b101000001: data <= 20'b11000100111100111000;
        10'b101000010: data <= 20'b10111110011100011011;
        10'b101000011: data <= 20'b01001010110011011011;
        10'b101000100: data <= 20'b11001001011100101011;
        10'b101000101: data <= 20'b01000000010100010011;
        10'b101000110: data <= 20'b11010100001011110101;
        10'b101000111: data <= 20'b01000010101100101001;
        10'b101001000: data <= 20'b01001100111100111101;
        10'b101001001: data <= 20'b11000110001100101101;
        10'b101001010: data <= 20'b01000110001100011000;
        10'b101001011: data <= 20'b01000011101101000011;
        10'b101001100: data <= 20'b11000101011100011000;
        10'b101001101: data <= 20'b01000010000100011000;
        10'b101001110: data <= 20'b11001100011100110111;
        10'b101001111: data <= 20'b01001011111100010001;
        10'b101010000: data <= 20'b11001001101101000111;
        10'b101010001: data <= 20'b00111101011100100110;
        10'b101010010: data <= 20'b01001101011100110010;
        10'b101010011: data <= 20'b11001000111100110000;
        10'b101010100: data <= 20'b10101101001100010011;
        10'b101010101: data <= 20'b01001101000011100111;
        10'b101010110: data <= 20'b11000010101100011100;
        10'b101010111: data <= 20'b01001001100100101001;
        10'b101011000: data <= 20'b11001001011100110111;
        10'b101011001: data <= 20'b01001011011100100011;
        10'b101011010: data <= 20'b11001000111101000011;
        10'b101011011: data <= 20'b11000100011100100100;
        10'b101011100: data <= 20'b01001000101100010011;
        10'b101011101: data <= 20'b11000110001100111100;
        10'b101011110: data <= 20'b10111010111100001100;
        10'b101011111: data <= 20'b01001011110100100111;
        10'b101100000: data <= 20'b01000101101100100001;
        10'b101100001: data <= 20'b01010011100100011000;
        10'b101100010: data <= 20'b11001010001100110010;
        10'b101100011: data <= 20'b01000011011100011111;
        10'b101100100: data <= 20'b01001110111100111110;
        10'b101100101: data <= 20'b11000110011100101000;
        10'b101100110: data <= 20'b01000010001100010001;
        10'b101100111: data <= 20'b01001010101100110100;
        10'b101101000: data <= 20'b01000011100100000000;
        10'b101101001: data <= 20'b11010110100101011110;
        10'b101101010: data <= 20'b10111111001100100110;
        10'b101101011: data <= 20'b01001110001100010001;
        10'b101101100: data <= 20'b11001011011100111001;
        10'b101101101: data <= 20'b10111100011100100001;
        10'b101101110: data <= 20'b01001010001100100101;
        10'b101101111: data <= 20'b11000100101100101000;
        10'b101110000: data <= 20'b01000100110011111011;
        10'b101110001: data <= 20'b11001110111101001011;
        10'b101110010: data <= 20'b01000111000011100100;
        10'b101110011: data <= 20'b11011101100100110000;
        10'b101110100: data <= 20'b11000111011100101010;
        10'b101110101: data <= 20'b01000110111100100000;
        10'b101110110: data <= 20'b01000000101100111111;
        10'b101110111: data <= 20'b10111101111100100001;
        10'b101111000: data <= 20'b01001010001100010111;
        10'b101111001: data <= 20'b11000100111100100101;
        10'b101111010: data <= 20'b01000100010100100100;
        10'b101111011: data <= 20'b11010000101100110010;
        10'b101111100: data <= 20'b00111110101100100011;
        10'b101111101: data <= 20'b01001111101100101111;
        10'b101111110: data <= 20'b11000111001100110001;
        10'b101111111: data <= 20'b01000011111100100010;
        10'b110000000: data <= 20'b01000101101100111000;
        10'b110000001: data <= 20'b11000010001100010011;
        10'b110000010: data <= 20'b01000110100100101000;
        10'b110000011: data <= 20'b11001001111100101100;
        10'b110000100: data <= 20'b01001001100100000100;
        10'b110000101: data <= 20'b11010000111101001000;
        10'b110000110: data <= 20'b10111111001100101001;
        10'b110000111: data <= 20'b01001001111100101110;
        10'b110001000: data <= 20'b11000101011100110001;
        10'b110001001: data <= 20'b01000000101100001111;
        10'b110001010: data <= 20'b01010000101100110000;
        10'b110001011: data <= 20'b11000100001100010001;
        10'b110001100: data <= 20'b01000100110100110010;
        10'b110001101: data <= 20'b11001011011100110010;
        10'b110001110: data <= 20'b01000111011100100110;
        10'b110001111: data <= 20'b01000101001101000001;
        10'b110010000: data <= 20'b11000000011100100110;
        10'b110010001: data <= 20'b01001010001100100000;
        10'b110010010: data <= 20'b11001000101100110100;
        10'b110010011: data <= 20'b10111110011011111101;
        10'b110010100: data <= 20'b01000101100100110111;
        10'b110010101: data <= 20'b10110111111100101000;
        10'b110010110: data <= 20'b01001111011100001010;
        10'b110010111: data <= 20'b11001000111100110110;
        10'b110011000: data <= 20'b01000101111100100100;
        10'b110011001: data <= 20'b01000111011101000001;
        10'b110011010: data <= 20'b11000101011100100100;
        10'b110011011: data <= 20'b01000011101011110011;
        10'b110011100: data <= 20'b01001100001101010010;
        10'b110011101: data <= 20'b00111111111011110011;
        10'b110011110: data <= 20'b01010000100101001110;
        10'b110011111: data <= 20'b10111001101100101110;
        10'b110100000: data <= 20'b01001101101100110001;
        10'b110100001: data <= 20'b11001001001100110101;
        10'b110100010: data <= 20'b10100000001100011100;
        10'b110100011: data <= 20'b01001101001100011101;
        10'b110100100: data <= 20'b11001000001100101011;
        10'b110100101: data <= 20'b00111110110011010000;
        10'b110100110: data <= 20'b01010100000101100000;
        10'b110100111: data <= 20'b01001001101100011010;
        10'b110101000: data <= 20'b01000100111101010011;
        10'b110101001: data <= 20'b11000100101100101001;
        10'b110101010: data <= 20'b01001001011100011100;
        10'b110101011: data <= 20'b11001000011101000001;
        10'b110101100: data <= 20'b11000010101100011101;
        10'b110101101: data <= 20'b01000111111011110011;
        10'b110101110: data <= 20'b10111110111100101111;
        10'b110101111: data <= 20'b01001001100100100000;
        10'b110110000: data <= 20'b11001101111101000000;
        10'b110110001: data <= 20'b01000101011100100001;
        10'b110110010: data <= 20'b01010001001101000011;
        10'b110110011: data <= 20'b11001000001100101101;
        10'b110110100: data <= 20'b00111111111100011001;
        10'b110110101: data <= 20'b01001100011100110011;
        10'b110110110: data <= 20'b11000001101100011100;
        10'b110110111: data <= 20'b01001001000100011011;
        10'b110111000: data <= 20'b11000100101100110000;
        10'b110111001: data <= 20'b01001100110100011001;
        10'b110111010: data <= 20'b11001110111100111110;
        10'b110111011: data <= 20'b11000000011100100100;
        10'b110111100: data <= 20'b01001011011100100001;
        10'b110111101: data <= 20'b11000111101100110100;
        10'b110111110: data <= 20'b00111100111100011000;
        10'b110111111: data <= 20'b01001100001100100110;
        10'b111000000: data <= 20'b10111100111100000010;
        10'b111000001: data <= 20'b01000111010101000000;
        10'b111000010: data <= 20'b11001001111100101110;
        10'b111000011: data <= 20'b01000111111100011010;
        10'b111000100: data <= 20'b01001010101101001010;
        10'b111000101: data <= 20'b11000100011100101001;
        10'b111000110: data <= 20'b01000110101100100001;
        10'b111000111: data <= 20'b11000001111100110010;
        10'b111001000: data <= 20'b00111000011011011110;
        10'b111001001: data <= 20'b01001001100101001011;
        10'b111001010: data <= 20'b10110010011100011011;
        10'b111001011: data <= 20'b01001111010100101110;
        10'b111001100: data <= 20'b11001011111100110101;
        10'b111001101: data <= 20'b00111111111100100101;
        10'b111001110: data <= 20'b01001001101100110110;
        10'b111001111: data <= 20'b11000011011100100101;
        10'b111010000: data <= 20'b01000110111100000001;
        10'b111010001: data <= 20'b11000111111101000000;
        10'b111010010: data <= 20'b00111001000100000010;
        10'b111010011: data <= 20'b11010000000101001011;
        10'b111010100: data <= 20'b11000101101100101010;
        10'b111010101: data <= 20'b01001010111100100111;
        10'b111010110: data <= 20'b11000110001100111000;
        10'b111010111: data <= 20'b00111101011100100001;
        10'b111011000: data <= 20'b01001100001100110001;
        10'b111011001: data <= 20'b11000111011100100100;
        10'b111011010: data <= 20'b00111010010100001110;
        10'b111011011: data <= 20'b11010010010100010111;
        10'b111011100: data <= 20'b01000101001100011000;
        10'b111011101: data <= 20'b01010100011101000001;
        10'b111011110: data <= 20'b11000100011100101111;
        10'b111011111: data <= 20'b01001001001100100111;
        10'b111100000: data <= 20'b11000110111100111000;
        10'b111100001: data <= 20'b11000000101100011000;
        10'b111100010: data <= 20'b01001001100100010011;
        10'b111100011: data <= 20'b11000111111100101011;
        10'b111100100: data <= 20'b01000110110100010011;
        10'b111100101: data <= 20'b11010010011101000110;
        10'b111100110: data <= 20'b01000011011100101001;
        10'b111100111: data <= 20'b01001100111101000000;
        10'b111101000: data <= 20'b11000110011100101011;
        10'b111101001: data <= 20'b01000100111100010100;
        10'b111101010: data <= 20'b01001011011101000100;
        10'b111101011: data <= 20'b11000100011100010110;
        10'b111101100: data <= 20'b01000100010100100000;
        10'b111101101: data <= 20'b11001010001100110111;
        10'b111101110: data <= 20'b01001100111100011100;
        10'b111101111: data <= 20'b11001010101101000000;
        10'b111110000: data <= 20'b00101111011100100011;
        10'b111110001: data <= 20'b01001101001100101001;
        10'b111110010: data <= 20'b11001001001100110001;
        10'b111110011: data <= 20'b10110110111100010000;
        10'b111110100: data <= 20'b01001100010100010011;
        10'b111110101: data <= 20'b00111011011100011001;
        10'b111110110: data <= 20'b01001111010100110100;
        10'b111110111: data <= 20'b11001000001100110001;
        10'b111111000: data <= 20'b01001010011100100000;
        10'b111111001: data <= 20'b11001001001101000101;
        10'b111111010: data <= 20'b11000100111100100100;
        10'b111111011: data <= 20'b01000111001100010000;
        10'b111111100: data <= 20'b11000000101100111100;
        10'b111111101: data <= 20'b00110111111100001000;
        10'b111111110: data <= 20'b01001110010100110010;
        10'b111111111: data <= 20'b01000100111100100001;
        10'b1000000000: data <= 20'b01010100000011100010;
        10'b1000000001: data <= 20'b11001010001100110001;
        10'b1000000010: data <= 20'b01000000101100011101;
        10'b1000000011: data <= 20'b01001110101100110111;
        10'b1000000100: data <= 20'b11000101111100100111;
        10'b1000000101: data <= 20'b01000011011100001110;
        10'b1000000110: data <= 20'b01001010001100110111;
        10'b1000000111: data <= 20'b01000101000100010001;
        10'b1000001000: data <= 20'b11010110110100100110;
        10'b1000001001: data <= 20'b11000001011100100101;
        10'b1000001010: data <= 20'b01001100111100010100;
        10'b1000001011: data <= 20'b11001010101100111011;
        10'b1000001100: data <= 20'b10111101001100100010;
        10'b1000001101: data <= 20'b01001001101100100100;
        10'b1000001110: data <= 20'b11000100011100100101;
        10'b1000001111: data <= 20'b01000101000100010100;
        10'b1000010000: data <= 20'b11010000001100111101;
        10'b1000010001: data <= 20'b01000110111100000000;
        10'b1000010010: data <= 20'b01011010011101110010;
        10'b1000010011: data <= 20'b11000111101100101100;
        10'b1000010100: data <= 20'b01000110001100100010;
        10'b1000010101: data <= 20'b01000001101100111010;
        10'b1000010110: data <= 20'b10111100001100011101;
        10'b1000010111: data <= 20'b01001011011011111011;
        10'b1000011000: data <= 20'b11000101011100100011;
        10'b1000011001: data <= 20'b01000101110100101001;
        10'b1000011010: data <= 20'b11010000011100110010;
        10'b1000011011: data <= 20'b00111000011100100100;
        10'b1000011100: data <= 20'b01001101101100110011;
        10'b1000011101: data <= 20'b11000101101100110000;
        10'b1000011110: data <= 20'b01000100101100100000;
        10'b1000011111: data <= 20'b01000101101100111010;
        10'b1000100000: data <= 20'b11000010011100010000;
        10'b1000100001: data <= 20'b01000100000100101110;
        10'b1000100010: data <= 20'b11001010001100101110;
        10'b1000100011: data <= 20'b01001010001100000011;
        10'b1000100100: data <= 20'b11001011011101001000;
        10'b1000100101: data <= 20'b10111011111100101000;
        10'b1000100110: data <= 20'b01001010011100110000;
        10'b1000100111: data <= 20'b11000110101100101111;
        10'b1000101000: data <= 20'b00111101001100000110;
        10'b1000101001: data <= 20'b01010001010100101000;
        10'b1000101010: data <= 20'b11000000011100010010;
        10'b1000101011: data <= 20'b01001010000100110101;
        10'b1000101100: data <= 20'b11001010001100110100;
        10'b1000101101: data <= 20'b01000111101100101010;
        10'b1000101110: data <= 20'b00011101111100111111;
        10'b1000101111: data <= 20'b11000000011100100011;
        10'b1000110000: data <= 20'b01001001101100010100;
        10'b1000110001: data <= 20'b11001001001100110101;
        10'b1000110010: data <= 20'b10111101011011011111;
        10'b1000110011: data <= 20'b11000000100100111111;
        10'b1000110100: data <= 20'b00110111101100101001;
        10'b1000110101: data <= 20'b01001111101100110001;
        10'b1000110110: data <= 20'b11000111111100110100;
        10'b1000110111: data <= 20'b01000101001100100001;
        10'b1000111000: data <= 20'b01001010001101000010;
        10'b1000111001: data <= 20'b11000110101100100011;
        10'b1000111010: data <= 20'b01000001001011101010;
        10'b1000111011: data <= 20'b01010101111101001000;
        10'b1000111100: data <= 20'b01000101111011110000;
        10'b1000111101: data <= 20'b01011100001101000001;
        10'b1000111110: data <= 20'b10111000001100101011;
        10'b1000111111: data <= 20'b01001101101100101110;
        10'b1001000000: data <= 20'b11001001101100110101;
        10'b1001000001: data <= 20'b10111010001100011011;
        10'b1001000010: data <= 20'b01001100001100010001;
        10'b1001000011: data <= 20'b11000110111100101001;
        10'b1001000100: data <= 20'b01000010110011111110;
        10'b1001000101: data <= 20'b11010100011101011101;
        10'b1001000110: data <= 20'b01001010011100011010;
        10'b1001000111: data <= 20'b11000100101101010010;
        10'b1001001000: data <= 20'b11000101101100101000;
        10'b1001001001: data <= 20'b01001000001100011001;
        10'b1001001010: data <= 20'b10111110001101000010;
        10'b1001001011: data <= 20'b11000010111100011110;
        10'b1001001100: data <= 20'b01000111011011100010;
        10'b1001001101: data <= 20'b00111100111100101011;
        10'b1001001110: data <= 20'b01001100100100101100;
        10'b1001001111: data <= 20'b11001100111100111001;
        10'b1001010000: data <= 20'b01000010011100100000;
        10'b1001010001: data <= 20'b01010000011100111001;
        10'b1001010010: data <= 20'b11001000101100101111;
        10'b1001010011: data <= 20'b01000000011100011001;
        10'b1001010100: data <= 20'b01001011001100110010;
        10'b1001010101: data <= 20'b10111101111100010011;
        10'b1001010110: data <= 20'b01001010110100101111;
        10'b1001010111: data <= 20'b11000101011100101011;
        10'b1001011000: data <= 20'b01001100100100001001;
        10'b1001011001: data <= 20'b11001110011101000001;
        10'b1001011010: data <= 20'b11000010001100100100;
        10'b1001011011: data <= 20'b01001001111100100010;
        10'b1001011100: data <= 20'b11000101001100110011;
        10'b1001011101: data <= 20'b00111111001100010010;
        10'b1001011110: data <= 20'b01001110101100100110;
        10'b1001011111: data <= 20'b10101110101011110001;
        10'b1001100000: data <= 20'b01000110000101000110;
        10'b1001100001: data <= 20'b11001001111100101110;
        10'b1001100010: data <= 20'b01000110001100100000;
        10'b1001100011: data <= 20'b01001011001101000011;
        10'b1001100100: data <= 20'b11000011011100100111;
        10'b1001100101: data <= 20'b01000111111100100000;
        10'b1001100110: data <= 20'b11000100101100110011;
        10'b1001100111: data <= 20'b00110111010011111101;
        10'b1001101000: data <= 20'b11010000010101001010;
        10'b1001101001: data <= 20'b10111101011100100001;
        10'b1001101010: data <= 20'b01001111000100000010;
        10'b1001101011: data <= 20'b11001010001100110111;
        10'b1001101100: data <= 20'b01000000111100100100;
        10'b1001101101: data <= 20'b01001000001100110111;
        10'b1001101110: data <= 20'b11000100001100100010;
        10'b1001101111: data <= 20'b01000110100011110110;
        10'b1001110000: data <= 20'b11001100101101000000;
        10'b1001110001: data <= 20'b01000000100011111100;
        10'b1001110010: data <= 20'b11010001110101010100;
        10'b1001110011: data <= 20'b11000100111100101101;
        10'b1001110100: data <= 20'b01001010011100101011;
        10'b1001110101: data <= 20'b11000101111100110101;
        10'b1001110110: data <= 20'b00111000101100011110;
        10'b1001110111: data <= 20'b01001101001100100101;
        10'b1001111000: data <= 20'b11000111101100100010;
        10'b1001111001: data <= 20'b00111100010100010111;
        10'b1001111010: data <= 20'b11010001001100100010;
        10'b1001111011: data <= 20'b01000101111100100010;
        10'b1001111100: data <= 20'b01001111011101000110;
        10'b1001111101: data <= 20'b11000011111100101100;
        10'b1001111110: data <= 20'b01001001001100100011;
        10'b1001111111: data <= 20'b11000111101100111011;
        10'b1010000000: data <= 20'b11000001101100010100;
        10'b1010000001: data <= 20'b01001000000100011010;
        10'b1010000010: data <= 20'b11001000001100101110;
        10'b1010000011: data <= 20'b01001001100100010011;
        10'b1010000100: data <= 20'b11001110011101000101;
        10'b1010000101: data <= 20'b01000100101100100111;
        10'b1010000110: data <= 20'b01001011101101000001;
        10'b1010000111: data <= 20'b11000111001100101001;
        10'b1010001000: data <= 20'b01000010011100001111;
        10'b1010001001: data <= 20'b01010000101101000001;
        10'b1010001010: data <= 20'b11000010101100010011;
        10'b1010001011: data <= 20'b01000110010100100111;
        10'b1010001100: data <= 20'b11001000011100110100;
        10'b1010001101: data <= 20'b01001101011100100010;
        10'b1010001110: data <= 20'b11001011001100111101;
        10'b1010001111: data <= 20'b10111011111100100010;
        10'b1010010000: data <= 20'b01001100101100100001;
        10'b1010010001: data <= 20'b11001000111100110010;
        10'b1010010010: data <= 20'b10111000111100001101;
        10'b1010010011: data <= 20'b01001100010100100001;
        10'b1010010100: data <= 20'b01000011111100010110;
        10'b1010010101: data <= 20'b01010011010100111000;
        10'b1010010110: data <= 20'b11000110101100110000;
        10'b1010010111: data <= 20'b01001000111100011100;
        10'b1010011000: data <= 20'b11000110011101000111;
        10'b1010011001: data <= 20'b11000101001100100100;
        10'b1010011010: data <= 20'b01000110001100010000;
        10'b1010011011: data <= 20'b00111000101100110111;
        10'b1010011100: data <= 20'b01000001011011100101;
        10'b1010011101: data <= 20'b01010100110101010010;
        10'b1010011110: data <= 20'b01000010011100100001;
        10'b1010011111: data <= 20'b01010010111100000011;
        10'b1010100000: data <= 20'b11001010001100110001;
        10'b1010100001: data <= 20'b00111100111100011111;
        10'b1010100010: data <= 20'b01001100111100101111;
        10'b1010100011: data <= 20'b11000101001100100111;
        10'b1010100100: data <= 20'b01000101011100000010;
        10'b1010100101: data <= 20'b01000100101100111011;
        10'b1010100110: data <= 20'b01000111000100010111;
        10'b1010100111: data <= 20'b11010101001100110111;
        10'b1010101000: data <= 20'b11000011111100100110;
        10'b1010101001: data <= 20'b01001010111100011110;
        10'b1010101010: data <= 20'b11001000011100111101;
        10'b1010101011: data <= 20'b10111011111100100001;
        10'b1010101100: data <= 20'b01001001011100100010;
        10'b1010101101: data <= 20'b11000100101100100001;
        10'b1010101110: data <= 20'b01000011100100100100;
        10'b1010101111: data <= 20'b11001110101100110000;
        10'b1010110000: data <= 20'b01000110001100010010;
        10'b1010110001: data <= 20'b01010101011101010101;
        10'b1010110010: data <= 20'b11000110011100101110;
        10'b1010110011: data <= 20'b01000101001100100011;
        10'b1010110100: data <= 20'b00111101101100110111;
        10'b1010110101: data <= 20'b10111100001100010100;
        10'b1010110110: data <= 20'b01001100000100011101;
        10'b1010110111: data <= 20'b11000101101100100010;
        10'b1010111000: data <= 20'b01001000100100101000;
        10'b1010111001: data <= 20'b11010000001100111000;
        10'b1010111010: data <= 20'b00110110101100100110;
        10'b1010111011: data <= 20'b01001100001100110011;
        10'b1010111100: data <= 20'b11000100111100101111;
        10'b1010111101: data <= 20'b01000100101100011001;
        10'b1010111110: data <= 20'b01001000001100111111;
        10'b1010111111: data <= 20'b11000011101100000111;
        10'b1011000000: data <= 20'b00111100010100110010;
        10'b1011000001: data <= 20'b11001001011100101110;
        10'b1011000010: data <= 20'b01001010001100011010;
        10'b1011000011: data <= 20'b11000110011101000100;
        10'b1011000100: data <= 20'b00110000011100100110;
        10'b1011000101: data <= 20'b01001011001100110000;
        10'b1011000110: data <= 20'b11000111101100101101;
        10'b1011000111: data <= 20'b00110010111011111000;
        10'b1011001000: data <= 20'b01001101110101000001;
        10'b1011001001: data <= 20'b10111011101100010101;
        10'b1011001010: data <= 20'b01001101100100110100;
        10'b1011001011: data <= 20'b11001001101100110100;
        10'b1011001100: data <= 20'b01001000001100101000;
        10'b1011001101: data <= 20'b10110110111101000000;
        10'b1011001110: data <= 20'b11000010111100100010;
        10'b1011001111: data <= 20'b01001000111100000010;
        10'b1011010000: data <= 20'b11001001101100110110;
        10'b1011010001: data <= 20'b10111001111011001011;
        10'b1011010010: data <= 20'b11000000010101000011;
        10'b1011010011: data <= 20'b00111111101100101011;
        10'b1011010100: data <= 20'b01001111001100111001;
        10'b1011010101: data <= 20'b11001000001100110010;
        10'b1011010110: data <= 20'b01000011101100011110;
        10'b1011010111: data <= 20'b01001101001100111111;
        10'b1011011000: data <= 20'b11000110101100100011;
        10'b1011011001: data <= 20'b01000001000011100110;
        10'b1011011010: data <= 20'b01000011011101100011;
        10'b1011011011: data <= 20'b01001001011100000110;
        10'b1011011100: data <= 20'b01001000001101010110;
        10'b1011011101: data <= 20'b10111101111100101000;
        10'b1011011110: data <= 20'b01001100111100100111;
        10'b1011011111: data <= 20'b11001001111100110110;
        10'b1011100000: data <= 20'b10111110001100011011;
        10'b1011100001: data <= 20'b01001010011011111110;
        10'b1011100010: data <= 20'b11000101011100101000;
        10'b1011100011: data <= 20'b01000110010100010110;
        10'b1011100100: data <= 20'b11001110001101000000;
        10'b1011100101: data <= 20'b01001001111100011110;
        10'b1011100110: data <= 20'b11000001111101010001;
        10'b1011100111: data <= 20'b11000110101100101000;
        10'b1011101000: data <= 20'b01000101111100011000;
        10'b1011101001: data <= 20'b01000100111101000001;
        10'b1011101010: data <= 20'b11000001011100011100;
        10'b1011101011: data <= 20'b01001000100011111000;
        10'b1011101100: data <= 20'b00111011101100100100;
        10'b1011101101: data <= 20'b01001110000100110011;
        10'b1011101110: data <= 20'b11001101001100110110;
        10'b1011101111: data <= 20'b00111111001100100001;
        10'b1011110000: data <= 20'b01001110101100110001;
        10'b1011110001: data <= 20'b11001000001100110000;
        10'b1011110010: data <= 20'b01000000001100011001;
        10'b1011110011: data <= 20'b01001010011100110000;
        10'b1011110100: data <= 20'b10110110101100000011;
        10'b1011110101: data <= 20'b01001010010101000000;
        10'b1011110110: data <= 20'b11000110001100101001;
        10'b1011110111: data <= 20'b01001100001011111001;
        10'b1011111000: data <= 20'b11001101001101000010;
        10'b1011111001: data <= 20'b11000001011100100101;
        10'b1011111010: data <= 20'b01001000111100100101;
        10'b1011111011: data <= 20'b11000100011100110000;
        10'b1011111100: data <= 20'b01000000101100000010;
        10'b1011111101: data <= 20'b01010100001100001000;
        10'b1011111110: data <= 20'b00111011011011111111;
        10'b1011111111: data <= 20'b01001100110101001000;
        10'b1100000000: data <= 20'b11001010001100110001;
        10'b1100000001: data <= 20'b01000100101100100010;
        10'b1100000010: data <= 20'b01001001101101000000;
        10'b1100000011: data <= 20'b11000001101100100110;
        10'b1100000100: data <= 20'b01001000101100011011;
        10'b1100000101: data <= 20'b11000110011100110001;
        10'b1100000110: data <= 20'b00110010010100001010;
        10'b1100000111: data <= 20'b11010001100101000001;
        10'b1100001000: data <= 20'b10111100111100100100;
        10'b1100001001: data <= 20'b01001110011100011010;
        10'b1100001010: data <= 20'b11001001001100110101;
        10'b1100001011: data <= 20'b01000010001100100100;
        10'b1100001100: data <= 20'b01001001011100110110;
        10'b1100001101: data <= 20'b11000100101100100000;
        10'b1100001110: data <= 20'b01000100110100010000;
        10'b1100001111: data <= 20'b11010000001100110101;
        10'b1100010000: data <= 20'b01000101010011011001;
        10'b1100010001: data <= 20'b11100000110110010010;
        10'b1100010010: data <= 20'b11000010111100101110;
        10'b1100010011: data <= 20'b01001001111100101101;
        10'b1100010100: data <= 20'b11000110101100110100;
        10'b1100010101: data <= 20'b00110000001100011000;
        10'b1100010110: data <= 20'b01001101101100010000;
        10'b1100010111: data <= 20'b11001000001100100010;
        10'b1100011000: data <= 20'b00111111110100011100;
        10'b1100011001: data <= 20'b11010000111100110001;
        10'b1100011010: data <= 20'b01000110011100100110;
        10'b1100011011: data <= 20'b01001010101101000101;
        10'b1100011100: data <= 20'b11000011111100101010;
        10'b1100011101: data <= 20'b01001000111100011101;
        10'b1100011110: data <= 20'b11000111001100111101;
        10'b1100011111: data <= 20'b11000010101100010100;
        10'b1100100000: data <= 20'b01000110000100100000;
        10'b1100100001: data <= 20'b11000110011100101110;
        10'b1100100010: data <= 20'b01001100100100000100;
        10'b1100100011: data <= 20'b11001011101101000000;
        10'b1100100100: data <= 20'b01000011111100100101;
        10'b1100100101: data <= 20'b01001100111101000000;
        10'b1100100110: data <= 20'b11000111101100101010;
        10'b1100100111: data <= 20'b00111111011100001011;
        10'b1100101000: data <= 20'b01010000111100101100;
        10'b1100101001: data <= 20'b10111101111100010100;
        10'b1100101010: data <= 20'b01001011010100110000;
        10'b1100101011: data <= 20'b11000001111100110010;
        10'b1100101100: data <= 20'b01001101011100100100;
        10'b1100101101: data <= 20'b11001011011100111011;
        10'b1100101110: data <= 20'b10111110111100100001;
        10'b1100101111: data <= 20'b01001011001100011001;
        10'b1100110000: data <= 20'b11001000011100110010;
        10'b1100110001: data <= 20'b10110101101100000111;
        10'b1100110010: data <= 20'b01001100100100101011;
        10'b1100110011: data <= 20'b01000111101100010000;
        10'b1100110100: data <= 20'b01011001101100110001;
        10'b1100110101: data <= 20'b11001000001100101111;
        10'b1100110110: data <= 20'b01000111011100011101;
        10'b1100110111: data <= 20'b01000110101101000111;
        10'b1100111000: data <= 20'b11000100011100100100;
        10'b1100111001: data <= 20'b01000101011100010001;
        10'b1100111010: data <= 20'b00111111011100110110;
        10'b1100111011: data <= 20'b01000100100100000111;
        10'b1100111100: data <= 20'b11011000101100111111;
        10'b1100111101: data <= 20'b00111110001100100001;
        10'b1100111110: data <= 20'b01010001001100010101;
        10'b1100111111: data <= 20'b11001010001100110011;
        10'b1101000000: data <= 20'b00111001101100100000;
        10'b1101000001: data <= 20'b01001011011100101101;
        10'b1101000010: data <= 20'b11000011101100100101;
        10'b1101000011: data <= 20'b01000110110011101000;
        10'b1101000100: data <= 20'b11000110111100111100;
        10'b1101000101: data <= 20'b01001000010100010110;
        10'b1101000110: data <= 20'b11010100011100111100;
        10'b1101000111: data <= 20'b11000100111100100111;
        10'b1101001000: data <= 20'b01001001101100100000;
        10'b1101001001: data <= 20'b11000101101100111011;
        10'b1101001010: data <= 20'b10101000011100100001;
        10'b1101001011: data <= 20'b01001010011100100100;
        10'b1101001100: data <= 20'b11000100011100011011;
        10'b1101001101: data <= 20'b01000011010100101011;
        10'b1101001110: data <= 20'b11001110011100110001;
        10'b1101001111: data <= 20'b01000100101100011101;
        10'b1101010000: data <= 20'b01010001011101000010;
        10'b1101010001: data <= 20'b11000101101100101110;
        10'b1101010010: data <= 20'b01000110001100100010;
        10'b1101010011: data <= 20'b10111110111100110111;
        10'b1101010100: data <= 20'b10111110111100001110;
        10'b1101010101: data <= 20'b01001001110100101111;
        10'b1101010110: data <= 20'b11000101001100100010;
        10'b1101010111: data <= 20'b01001011000100100011;
        10'b1101011000: data <= 20'b11001110111100111110;
        10'b1101011001: data <= 20'b00110010001100100111;
        10'b1101011010: data <= 20'b01001010001100110011;
        10'b1101011011: data <= 20'b11000100111100101100;
        10'b1101011100: data <= 20'b01000100011100010000;
        10'b1101011101: data <= 20'b01001100101101000110;
        10'b1101011110: data <= 20'b11000001111100000011;
        10'b1101011111: data <= 20'b00111110100100110111;
        10'b1101100000: data <= 20'b11001001001100110000;
        10'b1101100001: data <= 20'b01001001101100100100;
        10'b1101100010: data <= 20'b11000100111100111111;
        10'b1101100011: data <= 20'b00110000101100100100;
        10'b1101100100: data <= 20'b01001100001100101010;
        10'b1101100101: data <= 20'b11001000111100101100;
        10'b1101100110: data <= 20'b10110011001011100011;
        10'b1101100111: data <= 20'b01000110100101000100;
        10'b1101101000: data <= 20'b00111111111100011110;
        10'b1101101001: data <= 20'b01010001010100010001;
        10'b1101101010: data <= 20'b11000111011100110011;
        10'b1101101011: data <= 20'b01001000011100100110;
        10'b1101101100: data <= 20'b11000000011101000000;
        10'b1101101101: data <= 20'b11000011111100100000;
        10'b1101101110: data <= 20'b01000111011011100000;
        10'b1101101111: data <= 20'b11001001111100111101;
        10'b1101110000: data <= 20'b00111111100011110100;
        10'b1101110001: data <= 20'b11010000110101011001;
        10'b1101110010: data <= 20'b01000000011100101011;
        10'b1101110011: data <= 20'b01001110001100111011;
        10'b1101110100: data <= 20'b11001000011100110001;
        10'b1101110101: data <= 20'b01000001001100011011;
        10'b1101110110: data <= 20'b01001110101100110101;
        10'b1101110111: data <= 20'b11000110101100100011;
        10'b1101111000: data <= 20'b01000001100011111011;
        10'b1101111001: data <= 20'b11010001001101010011;
        10'b1101111010: data <= 20'b01001011001100000100;
        10'b1101111011: data <= 20'b11001101011101010000;
        10'b1101111100: data <= 20'b11000000001100100110;
        10'b1101111101: data <= 20'b01001100001100100001;
        10'b1101111110: data <= 20'b11001001111100111000;
        10'b1101111111: data <= 20'b10111111101100011011;
        10'b1110000000: data <= 20'b01001001011011111000;
        10'b1110000001: data <= 20'b11000011001100100110;
        10'b1110000010: data <= 20'b01001001100100100011;
        10'b1110000011: data <= 20'b11001100001100111010;
        10'b1110000100: data <= 20'b01001000111100011010;
        10'b1110000101: data <= 20'b01000101111101010010;
        10'b1110000110: data <= 20'b11000110101100101001;
        10'b1110000111: data <= 20'b01000100101100011000;
        10'b1110001000: data <= 20'b01001000001100111110;
        10'b1110001001: data <= 20'b10111100111100010110;
        10'b1110001010: data <= 20'b01001010110100010110;
        10'b1110001011: data <= 20'b10110100011100100101;
        10'b1110001100: data <= 20'b01001110100100101110;
        10'b1110001101: data <= 20'b11001100111100111000;
        10'b1110001110: data <= 20'b00111010101100100010;
        10'b1110001111: data <= 20'b01001100111100101111;
        10'b1110010000: data <= 20'b11000111011100101111;
        10'b1110010001: data <= 20'b01000001011100011000;
        10'b1110010010: data <= 20'b01001010111100110100;
        10'b1110010011: data <= 20'b10110111000011001010;
        10'b1110010100: data <= 20'b11000100110101000110;
        10'b1110010101: data <= 20'b11000111111100101001;
        10'b1110010110: data <= 20'b01001010101100001111;
        10'b1110010111: data <= 20'b11001010111101000101;
        10'b1110011000: data <= 20'b11000000111100100110;
        10'b1110011001: data <= 20'b01001000101100100100;
        10'b1110011010: data <= 20'b11000101001100101110;
        10'b1110011011: data <= 20'b01000001010011100101;
        10'b1110011100: data <= 20'b11011011000101110000;
        10'b1110011101: data <= 20'b00111110111100001010;
        10'b1110011110: data <= 20'b01010000110101000100;
        10'b1110011111: data <= 20'b11001001101100110001;
        10'b1110100000: data <= 20'b01000100101100100100;
        10'b1110100001: data <= 20'b01000111001100111010;
        10'b1110100010: data <= 20'b11000000011100100011;
        10'b1110100011: data <= 20'b01001001001100001010;
        10'b1110100100: data <= 20'b11001000111100110010;
        10'b1110100101: data <= 20'b00111001110100010000;
        10'b1110100110: data <= 20'b11010010010100111101;
        10'b1110100111: data <= 20'b11000000011100100111;
        10'b1110101000: data <= 20'b01001101001100101001;
        10'b1110101001: data <= 20'b11000110111100110100;
        10'b1110101010: data <= 20'b01000010101100100010;
        10'b1110101011: data <= 20'b01001010011100111000;
        10'b1110101100: data <= 20'b11000101101100011101;
        10'b1110101101: data <= 20'b01000000110100010111;
        10'b1110101110: data <= 20'b11001111101100101101;
        10'b1110101111: data <= 20'b01001000001100000011;
        10'b1110110000: data <= 20'b01001111011101011100;
        10'b1110110001: data <= 20'b11000001001100101100;
        10'b1110110010: data <= 20'b01001010001100101101;
        10'b1110110011: data <= 20'b11000111101100110100;
        10'b1110110100: data <= 20'b10111000011100010100;
        10'b1110110101: data <= 20'b01001100110100000101;
        10'b1110110110: data <= 20'b11000110101100100001;
        10'b1110110111: data <= 20'b01000101100100100001;
        10'b1110111000: data <= 20'b11001111101100111101;
        10'b1110111001: data <= 20'b01000110111100101000;
        10'b1110111010: data <= 20'b01001000001101000011;
        10'b1110111011: data <= 20'b11000100101100100111;
        10'b1110111100: data <= 20'b01001000001100010011;
        10'b1110111101: data <= 20'b11000110011101000000;
        10'b1110111110: data <= 20'b11000001101100010001;
        10'b1110111111: data <= 20'b01000110100100100101;
        10'b1111000000: data <= 20'b11000001011100110000;
        10'b1111000001: data <= 20'b01001110101100010011;
        10'b1111000010: data <= 20'b11001010011100111001;
        10'b1111000011: data <= 20'b01000010011100100010;
        10'b1111000100: data <= 20'b01001101111100111001;
        10'b1111000101: data <= 20'b11001000011100101011;
        10'b1111000110: data <= 20'b00111100111100001011;
        10'b1111000111: data <= 20'b01001111101100001101;
        10'b1111001000: data <= 20'b00110111111100001111;
        10'b1111001001: data <= 20'b01001110100100111101;
        10'b1111001010: data <= 20'b11000100011100110000;
        10'b1111001011: data <= 20'b01001100101100011101;
        10'b1111001100: data <= 20'b11001011111100111110;
        10'b1111001101: data <= 20'b11000001011100100001;
        10'b1111001110: data <= 20'b01001001101100010100;
        10'b1111001111: data <= 20'b11000111001100110100;
        10'b1111010000: data <= 20'b00111100011100000000;
        10'b1111010001: data <= 20'b01010000100100110111;
        10'b1111010010: data <= 20'b01001000001100010001;
        10'b1111010011: data <= 20'b01011001011101001001;
        10'b1111010100: data <= 20'b11001000101100101100;
        10'b1111010101: data <= 20'b01000101101100011100;
        10'b1111010110: data <= 20'b01001010011101000011;
        10'b1111010111: data <= 20'b11000100101100100101;
        10'b1111011000: data <= 20'b01000101111100001111;
        10'b1111011001: data <= 20'b00111011011100110010;
        10'b1111011010: data <= 20'b01000110000100011100;
        10'b1111011011: data <= 20'b11010011001100111000;
        10'b1111011100: data <= 20'b00110011001100100011;
        10'b1111011101: data <= 20'b01001111101100011111;
        10'b1111011110: data <= 20'b11001001101100110100;
        10'b1111011111: data <= 20'b00111000111100100000;
        10'b1111100000: data <= 20'b01001001111100101100;
        10'b1111100001: data <= 20'b11000011101100100001;
        10'b1111100010: data <= 20'b01000111010100010111;
        10'b1111100011: data <= 20'b11001011101100110101;
        10'b1111100100: data <= 20'b01001000110100000011;
        10'b1111100101: data <= 20'b11010101101101010000;
        10'b1111100110: data <= 20'b11000100101100100111;
        10'b1111100111: data <= 20'b01001000101100100011;
        10'b1111101000: data <= 20'b11000010101100111000;
        10'b1111101001: data <= 20'b00111001011100011100;
        10'b1111101010: data <= 20'b01001100011100100001;
        10'b1111101011: data <= 20'b11000100101100010110;
        10'b1111101100: data <= 20'b01000011100100110000;
        10'b1111101101: data <= 20'b11001101101100110001;
        10'b1111101110: data <= 20'b01000011011100100001;
        10'b1111101111: data <= 20'b01001110111101000000;
        10'b1111110000: data <= 20'b11000100101100101100;
        10'b1111110001: data <= 20'b01000110111100100010;
        10'b1111110010: data <= 20'b11000001111100110110;
        10'b1111110011: data <= 20'b11000000001100000100;
        10'b1111110100: data <= 20'b01000101110100110101;
        10'b1111110101: data <= 20'b11000110001100100110;
        10'b1111110110: data <= 20'b01001100000100000110;
        10'b1111110111: data <= 20'b11001100101101000001;
        10'b1111111000: data <= 20'b00111100111100100111;
        10'b1111111001: data <= 20'b01001010011100110110;
        10'b1111111010: data <= 20'b11000101101100101000;
        10'b1111111011: data <= 20'b01000011101011111011;
        10'b1111111100: data <= 20'b01001111111101010101;
    
    endcase
    end
    end

    assign Q = data;

    endmodule

        