
module memory_rom_44(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h32153e47;
    11'b00000000001: data <= 32'h317a3b30;
    11'b00000000010: data <= 32'had3cbb43;
    11'b00000000011: data <= 32'h38f9bf10;
    11'b00000000100: data <= 32'h3eb7b63e;
    11'b00000000101: data <= 32'h3f133e2d;
    11'b00000000110: data <= 32'h3c0c3e41;
    11'b00000000111: data <= 32'h3822b178;
    11'b00000001000: data <= 32'h355fbd3d;
    11'b00000001001: data <= 32'hb6c5babf;
    11'b00000001010: data <= 32'hbe07b48d;
    11'b00000001011: data <= 32'hbd6bbb9b;
    11'b00000001100: data <= 32'h359ebf7e;
    11'b00000001101: data <= 32'h3e55bdf0;
    11'b00000001110: data <= 32'h38f9ad10;
    11'b00000001111: data <= 32'hbd713acc;
    11'b00000010000: data <= 32'hbf9b3b96;
    11'b00000010001: data <= 32'hba2f3c34;
    11'b00000010010: data <= 32'hac113ce6;
    11'b00000010011: data <= 32'hba763891;
    11'b00000010100: data <= 32'hbdd1ba11;
    11'b00000010101: data <= 32'hb6ddbc48;
    11'b00000010110: data <= 32'h3d953678;
    11'b00000010111: data <= 32'h40253fcb;
    11'b00000011000: data <= 32'h3d723e67;
    11'b00000011001: data <= 32'h38b62788;
    11'b00000011010: data <= 32'h3523b81a;
    11'b00000011011: data <= 32'hae033594;
    11'b00000011100: data <= 32'hb98038d0;
    11'b00000011101: data <= 32'hb672bb37;
    11'b00000011110: data <= 32'h3b60c113;
    11'b00000011111: data <= 32'h3ea4c087;
    11'b00000100000: data <= 32'h3913b83e;
    11'b00000100001: data <= 32'hbb513914;
    11'b00000100010: data <= 32'hbc3a3864;
    11'b00000100011: data <= 32'hb0a03416;
    11'b00000100100: data <= 32'hb40234f3;
    11'b00000100101: data <= 32'hbf212839;
    11'b00000100110: data <= 32'hc133b9cf;
    11'b00000100111: data <= 32'hbca6ba72;
    11'b00000101000: data <= 32'h3c623624;
    11'b00000101001: data <= 32'h3f1d3e1e;
    11'b00000101010: data <= 32'h3a193d0d;
    11'b00000101011: data <= 32'hb0103624;
    11'b00000101100: data <= 32'ha82238ff;
    11'b00000101101: data <= 32'h310f3ecb;
    11'b00000101110: data <= 32'haee53de8;
    11'b00000101111: data <= 32'ha531b950;
    11'b00000110000: data <= 32'h3b1cc10a;
    11'b00000110001: data <= 32'h3e3dc00f;
    11'b00000110010: data <= 32'h3c2db037;
    11'b00000110011: data <= 32'h323839f0;
    11'b00000110100: data <= 32'h34822bbf;
    11'b00000110101: data <= 32'h39a2b8dc;
    11'b00000110110: data <= 32'hb1f2b625;
    11'b00000110111: data <= 32'hc04ab1f8;
    11'b00000111000: data <= 32'hc1acb9ca;
    11'b00000111001: data <= 32'hbc93bc84;
    11'b00000111010: data <= 32'h3bd9b82c;
    11'b00000111011: data <= 32'h3c96366b;
    11'b00000111100: data <= 32'hb42838ca;
    11'b00000111101: data <= 32'hbbef387b;
    11'b00000111110: data <= 32'hb5763d77;
    11'b00000111111: data <= 32'h338f40ca;
    11'b00001000000: data <= 32'hb2093f4a;
    11'b00001000001: data <= 32'hb8bcb675;
    11'b00001000010: data <= 32'h2da0bfa1;
    11'b00001000011: data <= 32'h3cabbc30;
    11'b00001000100: data <= 32'h3de439d5;
    11'b00001000101: data <= 32'h3cf13bfa;
    11'b00001000110: data <= 32'h3d45b349;
    11'b00001000111: data <= 32'h3d35bb1f;
    11'b00001001000: data <= 32'h2ea6b327;
    11'b00001001001: data <= 32'hbedf3440;
    11'b00001001010: data <= 32'hc034b8a4;
    11'b00001001011: data <= 32'hb78cbef6;
    11'b00001001100: data <= 32'h3c4ebeed;
    11'b00001001101: data <= 32'h38d3ba56;
    11'b00001001110: data <= 32'hbb7aac94;
    11'b00001001111: data <= 32'hbcff3624;
    11'b00001010000: data <= 32'hb1f73d06;
    11'b00001010001: data <= 32'h33f4401f;
    11'b00001010010: data <= 32'hbaa13de8;
    11'b00001010011: data <= 32'hbf36b484;
    11'b00001010100: data <= 32'hbc54bc9b;
    11'b00001010101: data <= 32'h38d1ac8b;
    11'b00001010110: data <= 32'h3e303d45;
    11'b00001010111: data <= 32'h3e163c29;
    11'b00001011000: data <= 32'h3dbbb42e;
    11'b00001011001: data <= 32'h3d47b6b4;
    11'b00001011010: data <= 32'h36e63a64;
    11'b00001011011: data <= 32'hbad13d13;
    11'b00001011100: data <= 32'hbbffb346;
    11'b00001011101: data <= 32'h3460c047;
    11'b00001011110: data <= 32'h3cbac0de;
    11'b00001011111: data <= 32'h36a5bd43;
    11'b00001100000: data <= 32'hba5fb5fc;
    11'b00001100001: data <= 32'hb8a4aa77;
    11'b00001100010: data <= 32'h386236b9;
    11'b00001100011: data <= 32'h35fd3c1b;
    11'b00001100100: data <= 32'hbe0d3a42;
    11'b00001100101: data <= 32'hc1b7b4b7;
    11'b00001100110: data <= 32'hbfa9b9c3;
    11'b00001100111: data <= 32'h31183258;
    11'b00001101000: data <= 32'h3cb23c55;
    11'b00001101001: data <= 32'h3b1038ea;
    11'b00001101010: data <= 32'h390db2ef;
    11'b00001101011: data <= 32'h3ab3369c;
    11'b00001101100: data <= 32'h390e401a;
    11'b00001101101: data <= 32'hb05c4088;
    11'b00001101110: data <= 32'hb58c3291;
    11'b00001101111: data <= 32'h36f7bffe;
    11'b00001110000: data <= 32'h3c12c050;
    11'b00001110001: data <= 32'h383bbaf4;
    11'b00001110010: data <= 32'h94b5b1ae;
    11'b00001110011: data <= 32'h3934b7e8;
    11'b00001110100: data <= 32'h3e25b86c;
    11'b00001110101: data <= 32'h396b2d7e;
    11'b00001110110: data <= 32'hbed835c1;
    11'b00001110111: data <= 32'hc218b42b;
    11'b00001111000: data <= 32'hbf8dba26;
    11'b00001111001: data <= 32'h2d6cb63e;
    11'b00001111010: data <= 32'h388c2cc7;
    11'b00001111011: data <= 32'hb367b251;
    11'b00001111100: data <= 32'hb747b504;
    11'b00001111101: data <= 32'h35303ba6;
    11'b00001111110: data <= 32'h39b24166;
    11'b00001111111: data <= 32'h27c54149;
    11'b00010000000: data <= 32'hb8d237a7;
    11'b00010000001: data <= 32'hb356bd89;
    11'b00010000010: data <= 32'h37b8bc5f;
    11'b00010000011: data <= 32'h394931eb;
    11'b00010000100: data <= 32'h3a7f345e;
    11'b00010000101: data <= 32'h3e8eba19;
    11'b00010000110: data <= 32'h4069bc37;
    11'b00010000111: data <= 32'h3c25ac1f;
    11'b00010001000: data <= 32'hbd01393f;
    11'b00010001001: data <= 32'hc07d2120;
    11'b00010001010: data <= 32'hbc37bc4b;
    11'b00010001011: data <= 32'h35b9bd64;
    11'b00010001100: data <= 32'h2b4fbc46;
    11'b00010001101: data <= 32'hbc65bbd2;
    11'b00010001110: data <= 32'hbc0fb8ed;
    11'b00010001111: data <= 32'h34db3a39;
    11'b00010010000: data <= 32'h3a9d409d;
    11'b00010010001: data <= 32'hb4e64059;
    11'b00010010010: data <= 32'hbe2b3736;
    11'b00010010011: data <= 32'hbd5eb94f;
    11'b00010010100: data <= 32'hb3162b0f;
    11'b00010010101: data <= 32'h38733c45;
    11'b00010010110: data <= 32'h3bf73812;
    11'b00010010111: data <= 32'h3ed5baf5;
    11'b00010011000: data <= 32'h404bbb00;
    11'b00010011001: data <= 32'h3d043965;
    11'b00010011010: data <= 32'hb6a23e5a;
    11'b00010011011: data <= 32'hbbe63825;
    11'b00010011100: data <= 32'ha6edbcff;
    11'b00010011101: data <= 32'h3959bfa9;
    11'b00010011110: data <= 32'hb1abbe3b;
    11'b00010011111: data <= 32'hbcf4bd05;
    11'b00010100000: data <= 32'hb91fbbee;
    11'b00010100001: data <= 32'h3b9aa960;
    11'b00010100010: data <= 32'h3c723c8d;
    11'b00010100011: data <= 32'hb9e73cde;
    11'b00010100100: data <= 32'hc0de3339;
    11'b00010100101: data <= 32'hc04cb2b4;
    11'b00010100110: data <= 32'hb98638b3;
    11'b00010100111: data <= 32'h31ea3c8c;
    11'b00010101000: data <= 32'h35a0322c;
    11'b00010101001: data <= 32'h3a57bbd2;
    11'b00010101010: data <= 32'h3dbab50a;
    11'b00010101011: data <= 32'h3cfd3ef4;
    11'b00010101100: data <= 32'h34de4121;
    11'b00010101101: data <= 32'had903c16;
    11'b00010101110: data <= 32'h3731bc38;
    11'b00010101111: data <= 32'h3922be6d;
    11'b00010110000: data <= 32'hb272bc12;
    11'b00010110001: data <= 32'hb9d1baeb;
    11'b00010110010: data <= 32'h361fbcfc;
    11'b00010110011: data <= 32'h3faebc06;
    11'b00010110100: data <= 32'h3e18a863;
    11'b00010110101: data <= 32'hbaa2378e;
    11'b00010110110: data <= 32'hc1222e0c;
    11'b00010110111: data <= 32'hc019b089;
    11'b00010111000: data <= 32'hb8f2349d;
    11'b00010111001: data <= 32'hb43c35bb;
    11'b00010111010: data <= 32'hba04b8c3;
    11'b00010111011: data <= 32'hb80ebcd9;
    11'b00010111100: data <= 32'h38c72ced;
    11'b00010111101: data <= 32'h3c8c409e;
    11'b00010111110: data <= 32'h387d41c9;
    11'b00010111111: data <= 32'haaa73ccd;
    11'b00011000000: data <= 32'h28f4b86f;
    11'b00011000001: data <= 32'h309eb861;
    11'b00011000010: data <= 32'hb3343364;
    11'b00011000011: data <= 32'hae86aea3;
    11'b00011000100: data <= 32'h3d17bd3c;
    11'b00011000101: data <= 32'h4120be4b;
    11'b00011000110: data <= 32'h3f5eb78f;
    11'b00011000111: data <= 32'hb6fe37d6;
    11'b00011001000: data <= 32'hbf0834d5;
    11'b00011001001: data <= 32'hbc2ab493;
    11'b00011001010: data <= 32'hab19b733;
    11'b00011001011: data <= 32'hb889b953;
    11'b00011001100: data <= 32'hbeabbd7a;
    11'b00011001101: data <= 32'hbd66be1c;
    11'b00011001110: data <= 32'h3467ad3c;
    11'b00011001111: data <= 32'h3ca13f9a;
    11'b00011010000: data <= 32'h3610408d;
    11'b00011010001: data <= 32'hb9fd3b4e;
    11'b00011010010: data <= 32'hbb73a862;
    11'b00011010011: data <= 32'hb8863918;
    11'b00011010100: data <= 32'hb6433d90;
    11'b00011010101: data <= 32'h2ab4373d;
    11'b00011010110: data <= 32'h3d43bd29;
    11'b00011010111: data <= 32'h40c6be23;
    11'b00011011000: data <= 32'h3f5d1e50;
    11'b00011011001: data <= 32'h32f83d02;
    11'b00011011010: data <= 32'hb78b3a88;
    11'b00011011011: data <= 32'h3415b5c8;
    11'b00011011100: data <= 32'h38b5bb88;
    11'b00011011101: data <= 32'hb92fbc79;
    11'b00011011110: data <= 32'hbfb9be43;
    11'b00011011111: data <= 32'hbcffbef1;
    11'b00011100000: data <= 32'h39c8b9fc;
    11'b00011100001: data <= 32'h3dc039a4;
    11'b00011100010: data <= 32'h2cb33c3e;
    11'b00011100011: data <= 32'hbe19359a;
    11'b00011100100: data <= 32'hbec133d6;
    11'b00011100101: data <= 32'hbbe63d1d;
    11'b00011100110: data <= 32'hb9383efd;
    11'b00011100111: data <= 32'hb79635db;
    11'b00011101000: data <= 32'h3609bd80;
    11'b00011101001: data <= 32'h3dbebc75;
    11'b00011101010: data <= 32'h3e033b5d;
    11'b00011101011: data <= 32'h39fb4054;
    11'b00011101100: data <= 32'h38363d35;
    11'b00011101101: data <= 32'h3c1fb30d;
    11'b00011101110: data <= 32'h3a99b9ae;
    11'b00011101111: data <= 32'hb8ffb875;
    11'b00011110000: data <= 32'hbe43bbc0;
    11'b00011110001: data <= 32'hb678beb9;
    11'b00011110010: data <= 32'h3e72be14;
    11'b00011110011: data <= 32'h3f69b86c;
    11'b00011110100: data <= 32'ha59b1f53;
    11'b00011110101: data <= 32'hbec5acf0;
    11'b00011110110: data <= 32'hbe463388;
    11'b00011110111: data <= 32'hb9f63c83;
    11'b00011111000: data <= 32'hba9f3cb2;
    11'b00011111001: data <= 32'hbd92b518;
    11'b00011111010: data <= 32'hbbfcbe7f;
    11'b00011111011: data <= 32'h34a2ba16;
    11'b00011111100: data <= 32'h3c463df5;
    11'b00011111101: data <= 32'h3b2c40f2;
    11'b00011111110: data <= 32'h39a83d66;
    11'b00011111111: data <= 32'h3ad92a79;
    11'b00100000000: data <= 32'h376231d4;
    11'b00100000001: data <= 32'hb9503a12;
    11'b00100000010: data <= 32'hbc0d2e3f;
    11'b00100000011: data <= 32'h3732bd9c;
    11'b00100000100: data <= 32'h4078bfce;
    11'b00100000101: data <= 32'h4029bc87;
    11'b00100000110: data <= 32'h321bb3ae;
    11'b00100000111: data <= 32'hbc1ba958;
    11'b00100001000: data <= 32'hb8012e3f;
    11'b00100001001: data <= 32'h2ee637d2;
    11'b00100001010: data <= 32'hba4b3305;
    11'b00100001011: data <= 32'hc04fbc49;
    11'b00100001100: data <= 32'hbfe8bf8c;
    11'b00100001101: data <= 32'hb52dba53;
    11'b00100001110: data <= 32'h3b003cca;
    11'b00100001111: data <= 32'h399a3f38;
    11'b00100010000: data <= 32'h30243a5f;
    11'b00100010001: data <= 32'ha11a339d;
    11'b00100010010: data <= 32'hb3013cd2;
    11'b00100010011: data <= 32'hba7c4019;
    11'b00100010100: data <= 32'hba3b3bba;
    11'b00100010101: data <= 32'h38aabc85;
    11'b00100010110: data <= 32'h400bbf7e;
    11'b00100010111: data <= 32'h3f63ba47;
    11'b00100011000: data <= 32'h3846361b;
    11'b00100011001: data <= 32'h2e5736c7;
    11'b00100011010: data <= 32'h3b622677;
    11'b00100011011: data <= 32'h3c51a89d;
    11'b00100011100: data <= 32'hb8a2b4bf;
    11'b00100011101: data <= 32'hc0b4bcfc;
    11'b00100011110: data <= 32'hc008bf9d;
    11'b00100011111: data <= 32'haae5bcb5;
    11'b00100100000: data <= 32'h3c4f310d;
    11'b00100100001: data <= 32'h3686377f;
    11'b00100100010: data <= 32'hb91eae91;
    11'b00100100011: data <= 32'hba6a327a;
    11'b00100100100: data <= 32'hb9113f0b;
    11'b00100100101: data <= 32'hbb69411c;
    11'b00100100110: data <= 32'hbc433c61;
    11'b00100100111: data <= 32'hb2a5bc67;
    11'b00100101000: data <= 32'h3bafbddb;
    11'b00100101001: data <= 32'h3cb32dd7;
    11'b00100101010: data <= 32'h39dd3d32;
    11'b00100101011: data <= 32'h3bf33b46;
    11'b00100101100: data <= 32'h3f6e2c2f;
    11'b00100101101: data <= 32'h3e481368;
    11'b00100101110: data <= 32'hb66b3020;
    11'b00100101111: data <= 32'hbff4b877;
    11'b00100110000: data <= 32'hbcf1be22;
    11'b00100110001: data <= 32'h3a74be74;
    11'b00100110010: data <= 32'h3df6bbe0;
    11'b00100110011: data <= 32'h33f6ba03;
    11'b00100110100: data <= 32'hbbaaba94;
    11'b00100110101: data <= 32'hba6c9bdc;
    11'b00100110110: data <= 32'hb5253e64;
    11'b00100110111: data <= 32'hba884024;
    11'b00100111000: data <= 32'hbea23797;
    11'b00100111001: data <= 32'hbdd6bd5a;
    11'b00100111010: data <= 32'hb5afbc4c;
    11'b00100111011: data <= 32'h36ad3a27;
    11'b00100111100: data <= 32'h39273ed8;
    11'b00100111101: data <= 32'h3c963b47;
    11'b00100111110: data <= 32'h3f2f2dbf;
    11'b00100111111: data <= 32'h3d3f38b5;
    11'b00101000000: data <= 32'hb6913d45;
    11'b00101000001: data <= 32'hbdae3965;
    11'b00101000010: data <= 32'hb4edbb49;
    11'b00101000011: data <= 32'h3e15bf16;
    11'b00101000100: data <= 32'h3ec6be14;
    11'b00101000101: data <= 32'h341cbc8d;
    11'b00101000110: data <= 32'hb88abb84;
    11'b00101000111: data <= 32'h306bb273;
    11'b00101001000: data <= 32'h39803ba1;
    11'b00101001001: data <= 32'hb6ce3c4e;
    11'b00101001010: data <= 32'hc03eb599;
    11'b00101001011: data <= 32'hc0c2be62;
    11'b00101001100: data <= 32'hbc85bb87;
    11'b00101001101: data <= 32'h254d39c8;
    11'b00101001110: data <= 32'h35973cae;
    11'b00101001111: data <= 32'h388b32f5;
    11'b00101010000: data <= 32'h3b69ac2d;
    11'b00101010001: data <= 32'h38b03d35;
    11'b00101010010: data <= 32'hb8834114;
    11'b00101010011: data <= 32'hbc3f3ee4;
    11'b00101010100: data <= 32'h290bb635;
    11'b00101010101: data <= 32'h3dbcbe35;
    11'b00101010110: data <= 32'h3d60bcac;
    11'b00101010111: data <= 32'h346bb861;
    11'b00101011000: data <= 32'h33eab768;
    11'b00101011001: data <= 32'h3df3b43e;
    11'b00101011010: data <= 32'h3f693570;
    11'b00101011011: data <= 32'h2ca7360e;
    11'b00101011100: data <= 32'hc047b938;
    11'b00101011101: data <= 32'hc0d0be19;
    11'b00101011110: data <= 32'hbb69bc1f;
    11'b00101011111: data <= 32'h3216a289;
    11'b00101100000: data <= 32'h2adbad87;
    11'b00101100001: data <= 32'hb434bb10;
    11'b00101100010: data <= 32'ha3a7b6c3;
    11'b00101100011: data <= 32'h29d83e90;
    11'b00101100100: data <= 32'hb8fe420e;
    11'b00101100101: data <= 32'hbc593fd0;
    11'b00101100110: data <= 32'hb755b46b;
    11'b00101100111: data <= 32'h375ebc77;
    11'b00101101000: data <= 32'h3790b3f8;
    11'b00101101001: data <= 32'h304037c4;
    11'b00101101010: data <= 32'h3b2f3073;
    11'b00101101011: data <= 32'h40ceb408;
    11'b00101101100: data <= 32'h40f530f4;
    11'b00101101101: data <= 32'h362b3837;
    11'b00101101110: data <= 32'hbedeac23;
    11'b00101101111: data <= 32'hbe62bbbf;
    11'b00101110000: data <= 32'h23b2bc77;
    11'b00101110001: data <= 32'h399dbb21;
    11'b00101110010: data <= 32'haf3ebd25;
    11'b00101110011: data <= 32'hba1fbf17;
    11'b00101110100: data <= 32'hb45dba87;
    11'b00101110101: data <= 32'h33cb3d8c;
    11'b00101110110: data <= 32'hb5a5410b;
    11'b00101110111: data <= 32'hbd583d27;
    11'b00101111000: data <= 32'hbdbbb8af;
    11'b00101111001: data <= 32'hbaa6b9d1;
    11'b00101111010: data <= 32'hb7c138a5;
    11'b00101111011: data <= 32'hb2353c89;
    11'b00101111100: data <= 32'h3b6b343e;
    11'b00101111101: data <= 32'h40a8b5bc;
    11'b00101111110: data <= 32'h407036ac;
    11'b00101111111: data <= 32'h35713dbb;
    11'b00110000000: data <= 32'hbc963c8a;
    11'b00110000001: data <= 32'hb858b019;
    11'b00110000010: data <= 32'h3b8bbbf5;
    11'b00110000011: data <= 32'h3c27bd14;
    11'b00110000100: data <= 32'hb286beac;
    11'b00110000101: data <= 32'hb965bfbd;
    11'b00110000110: data <= 32'h362abc18;
    11'b00110000111: data <= 32'h3cd539db;
    11'b00110001000: data <= 32'h342f3db4;
    11'b00110001001: data <= 32'hbdf43460;
    11'b00110001010: data <= 32'hc055bbd7;
    11'b00110001011: data <= 32'hbe70b831;
    11'b00110001100: data <= 32'hbbcc3a72;
    11'b00110001101: data <= 32'hb8693af9;
    11'b00110001110: data <= 32'h351bb5e1;
    11'b00110001111: data <= 32'h3d82b9d6;
    11'b00110010000: data <= 32'h3d543a6a;
    11'b00110010001: data <= 32'h2abe40e4;
    11'b00110010010: data <= 32'hb9f64063;
    11'b00110010011: data <= 32'h2a553845;
    11'b00110010100: data <= 32'h3c87b93d;
    11'b00110010101: data <= 32'h3a22baeb;
    11'b00110010110: data <= 32'hb627bc13;
    11'b00110010111: data <= 32'hb22bbd58;
    11'b00110011000: data <= 32'h3e0abbbf;
    11'b00110011001: data <= 32'h40c52de7;
    11'b00110011010: data <= 32'h3b7f3811;
    11'b00110011011: data <= 32'hbd53b4d3;
    11'b00110011100: data <= 32'hc03abc0a;
    11'b00110011101: data <= 32'hbd79b701;
    11'b00110011110: data <= 32'hb9d63668;
    11'b00110011111: data <= 32'hba10b0bc;
    11'b00110100000: data <= 32'hb83abdeb;
    11'b00110100001: data <= 32'h33ccbd2c;
    11'b00110100010: data <= 32'h38373b60;
    11'b00110100011: data <= 32'hb02741a8;
    11'b00110100100: data <= 32'hb8fc40d0;
    11'b00110100101: data <= 32'hb01238f9;
    11'b00110100110: data <= 32'h3686b448;
    11'b00110100111: data <= 32'haef32cb0;
    11'b00110101000: data <= 32'hba0531c5;
    11'b00110101001: data <= 32'h327eb7c0;
    11'b00110101010: data <= 32'h4098ba89;
    11'b00110101011: data <= 32'h4208b2b2;
    11'b00110101100: data <= 32'h3d1d3597;
    11'b00110101101: data <= 32'hbb492656;
    11'b00110101110: data <= 32'hbd19b771;
    11'b00110101111: data <= 32'hb490b4ad;
    11'b00110110000: data <= 32'h1f4cb23e;
    11'b00110110001: data <= 32'hba3ebccf;
    11'b00110110010: data <= 32'hbc7ac0c8;
    11'b00110110011: data <= 32'hb4dfbf14;
    11'b00110110100: data <= 32'h373838f3;
    11'b00110110101: data <= 32'h2eb9408f;
    11'b00110110110: data <= 32'hb92c3e7f;
    11'b00110110111: data <= 32'hba662fa8;
    11'b00110111000: data <= 32'hb9c5a3f7;
    11'b00110111001: data <= 32'hbc6b3bc6;
    11'b00110111010: data <= 32'hbcd93c67;
    11'b00110111011: data <= 32'h3041acd8;
    11'b00110111100: data <= 32'h4056badd;
    11'b00110111101: data <= 32'h4155b0f4;
    11'b00110111110: data <= 32'h3c543b8b;
    11'b00110111111: data <= 32'hb7583c2c;
    11'b00111000000: data <= 32'hb14336ba;
    11'b00111000001: data <= 32'h3b2d1c5b;
    11'b00111000010: data <= 32'h390ab6d6;
    11'b00111000011: data <= 32'hba3bbe13;
    11'b00111000100: data <= 32'hbcdac100;
    11'b00111000101: data <= 32'h28cfbf80;
    11'b00111000110: data <= 32'h3cda2aea;
    11'b00111000111: data <= 32'h3a153c88;
    11'b00111001000: data <= 32'hb8c135fd;
    11'b00111001001: data <= 32'hbd61b87a;
    11'b00111001010: data <= 32'hbdb02cb4;
    11'b00111001011: data <= 32'hbe4d3d6e;
    11'b00111001100: data <= 32'hbe193c9d;
    11'b00111001101: data <= 32'hb6beb7c6;
    11'b00111001110: data <= 32'h3caebd06;
    11'b00111001111: data <= 32'h3e45213f;
    11'b00111010000: data <= 32'h38293eef;
    11'b00111010001: data <= 32'hb1ec4005;
    11'b00111010010: data <= 32'h388c3c62;
    11'b00111010011: data <= 32'h3d9935c2;
    11'b00111010100: data <= 32'h38d2a841;
    11'b00111010101: data <= 32'hbbb9ba96;
    11'b00111010110: data <= 32'hbba4bee0;
    11'b00111010111: data <= 32'h3b51be44;
    11'b00111011000: data <= 32'h4092b73b;
    11'b00111011001: data <= 32'h3de52dfb;
    11'b00111011010: data <= 32'hb5d9b81a;
    11'b00111011011: data <= 32'hbd08bad8;
    11'b00111011100: data <= 32'hbc88307a;
    11'b00111011101: data <= 32'hbcbe3cb0;
    11'b00111011110: data <= 32'hbe0f366a;
    11'b00111011111: data <= 32'hbc90bde7;
    11'b00111100000: data <= 32'hac83bf7f;
    11'b00111100001: data <= 32'h374c21e4;
    11'b00111100010: data <= 32'h2a8a4014;
    11'b00111100011: data <= 32'haf294058;
    11'b00111100100: data <= 32'h38d13c51;
    11'b00111100101: data <= 32'h3bae389f;
    11'b00111100110: data <= 32'hb02a3a5b;
    11'b00111100111: data <= 32'hbd943789;
    11'b00111101000: data <= 32'hb9b8b895;
    11'b00111101001: data <= 32'h3e5abc76;
    11'b00111101010: data <= 32'h41bab96a;
    11'b00111101011: data <= 32'h3f03b438;
    11'b00111101100: data <= 32'habb0b7ce;
    11'b00111101101: data <= 32'hb802b7ac;
    11'b00111101110: data <= 32'h2888357c;
    11'b00111101111: data <= 32'hb1903a12;
    11'b00111110000: data <= 32'hbcf2b80e;
    11'b00111110001: data <= 32'hbe88c0ac;
    11'b00111110010: data <= 32'hba6cc0a7;
    11'b00111110011: data <= 32'h2c0db370;
    11'b00111110100: data <= 32'h2d743e2a;
    11'b00111110101: data <= 32'hadef3d41;
    11'b00111110110: data <= 32'h30313548;
    11'b00111110111: data <= 32'h1fea3857;
    11'b00111111000: data <= 32'hbc473e54;
    11'b00111111001: data <= 32'hbf793e3f;
    11'b00111111010: data <= 32'hba3d3141;
    11'b00111111011: data <= 32'h3de9bb61;
    11'b00111111100: data <= 32'h40e5b921;
    11'b00111111101: data <= 32'h3d602f95;
    11'b00111111110: data <= 32'h302a352f;
    11'b00111111111: data <= 32'h37f9356d;
    11'b01000000000: data <= 32'h3d823978;
    11'b01000000001: data <= 32'h3a433896;
    11'b01000000010: data <= 32'hbbc6ba7d;
    11'b01000000011: data <= 32'hbedfc0c7;
    11'b01000000100: data <= 32'hb964c086;
    11'b01000000101: data <= 32'h38b8b892;
    11'b01000000110: data <= 32'h393a37f3;
    11'b01000000111: data <= 32'h2579ad84;
    11'b01000001000: data <= 32'hb52bb977;
    11'b01000001001: data <= 32'hb933358c;
    11'b01000001010: data <= 32'hbe013fbd;
    11'b01000001011: data <= 32'hc01e3f4e;
    11'b01000001100: data <= 32'hbc9c2476;
    11'b01000001101: data <= 32'h388dbcd2;
    11'b01000001110: data <= 32'h3cd7b855;
    11'b01000001111: data <= 32'h37493a40;
    11'b01000010000: data <= 32'h2ed63cdd;
    11'b01000010001: data <= 32'h3cb53be0;
    11'b01000010010: data <= 32'h402e3bbc;
    11'b01000010011: data <= 32'h3c2f3ab1;
    11'b01000010100: data <= 32'hbc09b207;
    11'b01000010101: data <= 32'hbe13bdf1;
    11'b01000010110: data <= 32'h2a40be96;
    11'b01000010111: data <= 32'h3e3aba3b;
    11'b01000011000: data <= 32'h3d5db79c;
    11'b01000011001: data <= 32'h3324bcbc;
    11'b01000011010: data <= 32'hb505bd2e;
    11'b01000011011: data <= 32'hb6a13353;
    11'b01000011100: data <= 32'hbc093f2c;
    11'b01000011101: data <= 32'hbf173cfd;
    11'b01000011110: data <= 32'hbe57bab2;
    11'b01000011111: data <= 32'hb8c5bf2b;
    11'b01000100000: data <= 32'haf20b865;
    11'b01000100001: data <= 32'hb5a63c75;
    11'b01000100010: data <= 32'ha90f3da5;
    11'b01000100011: data <= 32'h3cf43b1d;
    11'b01000100100: data <= 32'h3f5d3b9c;
    11'b01000100101: data <= 32'h37b03d9b;
    11'b01000100110: data <= 32'hbd943c1c;
    11'b01000100111: data <= 32'hbd3fb05a;
    11'b01000101000: data <= 32'h39a8bab9;
    11'b01000101001: data <= 32'h404aba04;
    11'b01000101010: data <= 32'h3e41babd;
    11'b01000101011: data <= 32'h3580bd76;
    11'b01000101100: data <= 32'h32efbc7e;
    11'b01000101101: data <= 32'h396d35e1;
    11'b01000101110: data <= 32'h32313db7;
    11'b01000101111: data <= 32'hbc8c3643;
    11'b01000110000: data <= 32'hbf35bec0;
    11'b01000110001: data <= 32'hbd48c06b;
    11'b01000110010: data <= 32'hb9cdb943;
    11'b01000110011: data <= 32'hb8823a6d;
    11'b01000110100: data <= 32'haf5e38f8;
    11'b01000110101: data <= 32'h3a97a839;
    11'b01000110110: data <= 32'h3bcb388d;
    11'b01000110111: data <= 32'hb6d53f9d;
    11'b01000111000: data <= 32'hbf654031;
    11'b01000111001: data <= 32'hbd273aab;
    11'b01000111010: data <= 32'h39eeb5cb;
    11'b01000111011: data <= 32'h3f2ab8ac;
    11'b01000111100: data <= 32'h3c03b81e;
    11'b01000111101: data <= 32'h32bdb95e;
    11'b01000111110: data <= 32'h3b75b5d8;
    11'b01000111111: data <= 32'h3ff43994;
    11'b01001000000: data <= 32'h3d903cc9;
    11'b01001000001: data <= 32'hb869a45b;
    11'b01001000010: data <= 32'hbeddbf2f;
    11'b01001000011: data <= 32'hbcf4c00b;
    11'b01001000100: data <= 32'hb58ab9a6;
    11'b01001000101: data <= 32'hade82764;
    11'b01001000110: data <= 32'ha360b9f1;
    11'b01001000111: data <= 32'h35b8bd28;
    11'b01001001000: data <= 32'h34042711;
    11'b01001001001: data <= 32'hbb434019;
    11'b01001001010: data <= 32'hbfcc40cb;
    11'b01001001011: data <= 32'hbda53ae7;
    11'b01001001100: data <= 32'h2d4fb80b;
    11'b01001001101: data <= 32'h38bcb74a;
    11'b01001001110: data <= 32'haff9304e;
    11'b01001001111: data <= 32'hb18e33f0;
    11'b01001010000: data <= 32'h3d853520;
    11'b01001010001: data <= 32'h41753b61;
    11'b01001010010: data <= 32'h3f6c3d07;
    11'b01001010011: data <= 32'hb6783616;
    11'b01001010100: data <= 32'hbdd7bb7c;
    11'b01001010101: data <= 32'hb85abcb7;
    11'b01001010110: data <= 32'h38e2b864;
    11'b01001010111: data <= 32'h38f5b98f;
    11'b01001011000: data <= 32'h30f9bf74;
    11'b01001011001: data <= 32'h32c9c042;
    11'b01001011010: data <= 32'h34a4b521;
    11'b01001011011: data <= 32'hb7763f49;
    11'b01001011100: data <= 32'hbdd53f6b;
    11'b01001011101: data <= 32'hbdf42ae3;
    11'b01001011110: data <= 32'hba9abc5f;
    11'b01001011111: data <= 32'hb9fdb728;
    11'b01001100000: data <= 32'hbcbd38a1;
    11'b01001100001: data <= 32'hb8c138dd;
    11'b01001100010: data <= 32'h3d4a3488;
    11'b01001100011: data <= 32'h410b39e1;
    11'b01001100100: data <= 32'h3d7c3df5;
    11'b01001100101: data <= 32'hba143d5a;
    11'b01001100110: data <= 32'hbcf936d6;
    11'b01001100111: data <= 32'h320baea6;
    11'b01001101000: data <= 32'h3d55b2ac;
    11'b01001101001: data <= 32'h3b3ebb4b;
    11'b01001101010: data <= 32'h3082c02f;
    11'b01001101011: data <= 32'h371ec028;
    11'b01001101100: data <= 32'h3c87b403;
    11'b01001101101: data <= 32'h39ee3dc4;
    11'b01001101110: data <= 32'hb8633b9e;
    11'b01001101111: data <= 32'hbd73bb33;
    11'b01001110000: data <= 32'hbd7bbe4d;
    11'b01001110001: data <= 32'hbda9b74a;
    11'b01001110010: data <= 32'hbe3b3835;
    11'b01001110011: data <= 32'hba472b1c;
    11'b01001110100: data <= 32'h3b05b910;
    11'b01001110101: data <= 32'h3e882d88;
    11'b01001110110: data <= 32'h36463e89;
    11'b01001110111: data <= 32'hbd194069;
    11'b01001111000: data <= 32'hbc993dd0;
    11'b01001111001: data <= 32'h371438a0;
    11'b01001111010: data <= 32'h3ccc3004;
    11'b01001111011: data <= 32'h35d5b844;
    11'b01001111100: data <= 32'hb3b1bd97;
    11'b01001111101: data <= 32'h3a6bbd22;
    11'b01001111110: data <= 32'h4073301c;
    11'b01001111111: data <= 32'h3ffc3ca8;
    11'b01010000000: data <= 32'h346c35c6;
    11'b01010000001: data <= 32'hbc3bbcdb;
    11'b01010000010: data <= 32'hbcd8bdaf;
    11'b01010000011: data <= 32'hbc38b486;
    11'b01010000100: data <= 32'hbc5f2e44;
    11'b01010000101: data <= 32'hb942bc59;
    11'b01010000110: data <= 32'h3623bfc9;
    11'b01010000111: data <= 32'h3a18b9c6;
    11'b01010001000: data <= 32'hb4743e11;
    11'b01010001001: data <= 32'hbdb540cd;
    11'b01010001010: data <= 32'hbc563e13;
    11'b01010001011: data <= 32'h2f1f37d3;
    11'b01010001100: data <= 32'h332e3434;
    11'b01010001101: data <= 32'hba883069;
    11'b01010001110: data <= 32'hbb42b5cf;
    11'b01010001111: data <= 32'h3b9db6d7;
    11'b01010010000: data <= 32'h41ae36be;
    11'b01010010001: data <= 32'h41073c4a;
    11'b01010010010: data <= 32'h38383749;
    11'b01010010011: data <= 32'hb9ffb8a2;
    11'b01010010100: data <= 32'hb7dab849;
    11'b01010010101: data <= 32'ha2ba3137;
    11'b01010010110: data <= 32'hb395b4dd;
    11'b01010010111: data <= 32'hb691c020;
    11'b01010011000: data <= 32'h2fc5c1b5;
    11'b01010011001: data <= 32'h3835bce4;
    11'b01010011010: data <= 32'hac133cbf;
    11'b01010011011: data <= 32'hbb4a3f48;
    11'b01010011100: data <= 32'hbb093938;
    11'b01010011101: data <= 32'hb75fb2b0;
    11'b01010011110: data <= 32'hbba8324b;
    11'b01010011111: data <= 32'hbfd73959;
    11'b01010100000: data <= 32'hbe1c33ba;
    11'b01010100001: data <= 32'h39f2b3a1;
    11'b01010100010: data <= 32'h4128337f;
    11'b01010100011: data <= 32'h3fff3c2c;
    11'b01010100100: data <= 32'h2e873c4a;
    11'b01010100101: data <= 32'hb8ba38e7;
    11'b01010100110: data <= 32'h34ee390f;
    11'b01010100111: data <= 32'h3b6539f3;
    11'b01010101000: data <= 32'h3455b52e;
    11'b01010101001: data <= 32'hb660c072;
    11'b01010101010: data <= 32'h2fb9c19a;
    11'b01010101011: data <= 32'h3c21bc85;
    11'b01010101100: data <= 32'h3baf3ab8;
    11'b01010101101: data <= 32'h2def3ae8;
    11'b01010101110: data <= 32'hb7b6b7d1;
    11'b01010101111: data <= 32'hba26bb3b;
    11'b01010110000: data <= 32'hbe2c3074;
    11'b01010110001: data <= 32'hc0ba3a87;
    11'b01010110010: data <= 32'hbefe2203;
    11'b01010110011: data <= 32'h34c4bbac;
    11'b01010110100: data <= 32'h3e8fb7fb;
    11'b01010110101: data <= 32'h3adf3b30;
    11'b01010110110: data <= 32'hb8e43eac;
    11'b01010110111: data <= 32'hb8813e2f;
    11'b01010111000: data <= 32'h39d93d81;
    11'b01010111001: data <= 32'h3c643ca9;
    11'b01010111010: data <= 32'hac102e23;
    11'b01010111011: data <= 32'hbac4bdeb;
    11'b01010111100: data <= 32'h3200bf82;
    11'b01010111101: data <= 32'h3f55b897;
    11'b01010111110: data <= 32'h40383917;
    11'b01010111111: data <= 32'h3c063025;
    11'b01011000000: data <= 32'ha84ebc60;
    11'b01011000001: data <= 32'hb82fbbbe;
    11'b01011000010: data <= 32'hbc8935ac;
    11'b01011000011: data <= 32'hbf37395a;
    11'b01011000100: data <= 32'hbde9ba97;
    11'b01011000101: data <= 32'haffac04f;
    11'b01011000110: data <= 32'h392fbda7;
    11'b01011000111: data <= 32'had8f38b3;
    11'b01011001000: data <= 32'hbbee3eef;
    11'b01011001001: data <= 32'hb7b73e3d;
    11'b01011001010: data <= 32'h39503cef;
    11'b01011001011: data <= 32'h36f63cd1;
    11'b01011001100: data <= 32'hbc7439ac;
    11'b01011001101: data <= 32'hbe84b581;
    11'b01011001110: data <= 32'h2eb5ba1e;
    11'b01011001111: data <= 32'h408ca9d2;
    11'b01011010000: data <= 32'h41243873;
    11'b01011010001: data <= 32'h3cfba51b;
    11'b01011010010: data <= 32'h336cba34;
    11'b01011010011: data <= 32'h3149b34f;
    11'b01011010100: data <= 32'h9d4a3b54;
    11'b01011010101: data <= 32'hb9bb3835;
    11'b01011010110: data <= 32'hbbf7be61;
    11'b01011010111: data <= 32'hb596c202;
    11'b01011011000: data <= 32'h3220bfc5;
    11'b01011011001: data <= 32'hb21f33bb;
    11'b01011011010: data <= 32'hb9253c9a;
    11'b01011011011: data <= 32'hb17d38ed;
    11'b01011011100: data <= 32'h35df355a;
    11'b01011011101: data <= 32'hb8213b56;
    11'b01011011110: data <= 32'hc0653cbd;
    11'b01011011111: data <= 32'hc0a13753;
    11'b01011100000: data <= 32'hb1a1b41a;
    11'b01011100001: data <= 32'h3fe7a945;
    11'b01011100010: data <= 32'h3ff33711;
    11'b01011100011: data <= 32'h393d3510;
    11'b01011100100: data <= 32'h32413142;
    11'b01011100101: data <= 32'h3b3b3b00;
    11'b01011100110: data <= 32'h3c6e3e61;
    11'b01011100111: data <= 32'h2ecd390d;
    11'b01011101000: data <= 32'hba26bebd;
    11'b01011101001: data <= 32'hb684c1c8;
    11'b01011101010: data <= 32'h36babee8;
    11'b01011101011: data <= 32'h387c2ac5;
    11'b01011101100: data <= 32'h348e33f1;
    11'b01011101101: data <= 32'h358bb977;
    11'b01011101110: data <= 32'h3366b953;
    11'b01011101111: data <= 32'hbbfd3904;
    11'b01011110000: data <= 32'hc11a3d71;
    11'b01011110001: data <= 32'hc0eb37eb;
    11'b01011110010: data <= 32'hb813b980;
    11'b01011110011: data <= 32'h3c4fb96d;
    11'b01011110100: data <= 32'h39a23155;
    11'b01011110101: data <= 32'hb596399e;
    11'b01011110110: data <= 32'ha49e3bb4;
    11'b01011110111: data <= 32'h3d513e54;
    11'b01011111000: data <= 32'h3e243ff7;
    11'b01011111001: data <= 32'h2ce13bee;
    11'b01011111010: data <= 32'hbc60bbb3;
    11'b01011111011: data <= 32'hb778bf5c;
    11'b01011111100: data <= 32'h3bdfbb38;
    11'b01011111101: data <= 32'h3e2f2db4;
    11'b01011111110: data <= 32'h3cadb787;
    11'b01011111111: data <= 32'h3a8fbe1f;
    11'b01100000000: data <= 32'h3794bc30;
    11'b01100000001: data <= 32'hb8b6398a;
    11'b01100000010: data <= 32'hbf8a3d4d;
    11'b01100000011: data <= 32'hbfceada4;
    11'b01100000100: data <= 32'hb9a1bec6;
    11'b01100000101: data <= 32'h2f27be42;
    11'b01100000110: data <= 32'hb78fb2c4;
    11'b01100000111: data <= 32'hbc3b39b8;
    11'b01100001000: data <= 32'haf633b9d;
    11'b01100001001: data <= 32'h3d6c3d6a;
    11'b01100001010: data <= 32'h3c893f59;
    11'b01100001011: data <= 32'hba163d9b;
    11'b01100001100: data <= 32'hbf5f3092;
    11'b01100001101: data <= 32'hb92eb80f;
    11'b01100001110: data <= 32'h3d4ca8cc;
    11'b01100001111: data <= 32'h3fd632de;
    11'b01100010000: data <= 32'h3d62b987;
    11'b01100010001: data <= 32'h3b8cbde9;
    11'b01100010010: data <= 32'h3bf8b85d;
    11'b01100010011: data <= 32'h38173cd2;
    11'b01100010100: data <= 32'hb8bf3d32;
    11'b01100010101: data <= 32'hbc8ab9be;
    11'b01100010110: data <= 32'hb99cc0f1;
    11'b01100010111: data <= 32'hb650c01b;
    11'b01100011000: data <= 32'hbac8b783;
    11'b01100011001: data <= 32'hbbcd3405;
    11'b01100011010: data <= 32'h2ffc2769;
    11'b01100011011: data <= 32'h3cbc3459;
    11'b01100011100: data <= 32'h35b13ce9;
    11'b01100011101: data <= 32'hbeff3e8e;
    11'b01100011110: data <= 32'hc1023bcc;
    11'b01100011111: data <= 32'hbb243460;
    11'b01100100000: data <= 32'h3c61342f;
    11'b01100100001: data <= 32'h3d883265;
    11'b01100100010: data <= 32'h38c5b7ad;
    11'b01100100011: data <= 32'h38e6b9e9;
    11'b01100100100: data <= 32'h3dff370c;
    11'b01100100101: data <= 32'h3e8f3f7f;
    11'b01100100110: data <= 32'h38023daa;
    11'b01100100111: data <= 32'hb8b0baa3;
    11'b01100101000: data <= 32'hb900c0b5;
    11'b01100101001: data <= 32'hb482bed2;
    11'b01100101010: data <= 32'hb51fb66c;
    11'b01100101011: data <= 32'hb221b6e6;
    11'b01100101100: data <= 32'h391abd1d;
    11'b01100101101: data <= 32'h3c66bbf6;
    11'b01100101110: data <= 32'haebc38c7;
    11'b01100101111: data <= 32'hc02e3e96;
    11'b01100110000: data <= 32'hc1193c74;
    11'b01100110001: data <= 32'hbc0e2d93;
    11'b01100110010: data <= 32'h363fb259;
    11'b01100110011: data <= 32'h2e08ac11;
    11'b01100110100: data <= 32'hb953b1b0;
    11'b01100110101: data <= 32'h2a3398ba;
    11'b01100110110: data <= 32'h3eec3c7f;
    11'b01100110111: data <= 32'h404e4068;
    11'b01100111000: data <= 32'h39dc3e76;
    11'b01100111001: data <= 32'hb996b451;
    11'b01100111010: data <= 32'hb93bbd2f;
    11'b01100111011: data <= 32'h31b2b918;
    11'b01100111100: data <= 32'h3886a41d;
    11'b01100111101: data <= 32'h3940bb84;
    11'b01100111110: data <= 32'h3c4dc066;
    11'b01100111111: data <= 32'h3cf1be9c;
    11'b01101000000: data <= 32'h31af3695;
    11'b01101000001: data <= 32'hbdad3e37;
    11'b01101000010: data <= 32'hbf483925;
    11'b01101000011: data <= 32'hbafcba46;
    11'b01101000100: data <= 32'hb5babc1e;
    11'b01101000101: data <= 32'hbc97b6e0;
    11'b01101000110: data <= 32'hbea8af1e;
    11'b01101000111: data <= 32'hb55d2cc8;
    11'b01101001000: data <= 32'h3eac3b2b;
    11'b01101001001: data <= 32'h3f763f71;
    11'b01101001010: data <= 32'h2bd23edd;
    11'b01101001011: data <= 32'hbd7638f8;
    11'b01101001100: data <= 32'hbaae2e12;
    11'b01101001101: data <= 32'h38363839;
    11'b01101001110: data <= 32'h3c1c36d7;
    11'b01101001111: data <= 32'h3aafbc2a;
    11'b01101010000: data <= 32'h3c32c085;
    11'b01101010001: data <= 32'h3df3bd63;
    11'b01101010010: data <= 32'h3c4c3a7e;
    11'b01101010011: data <= 32'hace63e1d;
    11'b01101010100: data <= 32'hb99a293a;
    11'b01101010101: data <= 32'hb838be4c;
    11'b01101010110: data <= 32'hb9bfbe14;
    11'b01101010111: data <= 32'hbe8bb8a0;
    11'b01101011000: data <= 32'hbf3bb59d;
    11'b01101011001: data <= 32'hb3d2b951;
    11'b01101011010: data <= 32'h3df4b351;
    11'b01101011011: data <= 32'h3c913ba9;
    11'b01101011100: data <= 32'hbb403e64;
    11'b01101011101: data <= 32'hc00d3d24;
    11'b01101011110: data <= 32'hbc083be6;
    11'b01101011111: data <= 32'h37893c57;
    11'b01101100000: data <= 32'h38e238d5;
    11'b01101100001: data <= 32'h2ae8ba73;
    11'b01101100010: data <= 32'h371fbe61;
    11'b01101100011: data <= 32'h3e8cb6a2;
    11'b01101100100: data <= 32'h400a3de3;
    11'b01101100101: data <= 32'h3c813e6a;
    11'b01101100110: data <= 32'h305cb251;
    11'b01101100111: data <= 32'hb2dfbe5c;
    11'b01101101000: data <= 32'hb878bc9a;
    11'b01101101001: data <= 32'hbcccb445;
    11'b01101101010: data <= 32'hbc75b993;
    11'b01101101011: data <= 32'h33d0bf23;
    11'b01101101100: data <= 32'h3d8cbe66;
    11'b01101101101: data <= 32'h38c72416;
    11'b01101101110: data <= 32'hbd6b3d4e;
    11'b01101101111: data <= 32'hc0203d66;
    11'b01101110000: data <= 32'hbb623b40;
    11'b01101110001: data <= 32'h2cd53a0e;
    11'b01101110010: data <= 32'hb7e83645;
    11'b01101110011: data <= 32'hbd3ab7ff;
    11'b01101110100: data <= 32'hb710ba82;
    11'b01101110101: data <= 32'h3e3a35a4;
    11'b01101110110: data <= 32'h40de3f3a;
    11'b01101110111: data <= 32'h3de63e8c;
    11'b01101111000: data <= 32'h325a2d96;
    11'b01101111001: data <= 32'hb0f9b9ab;
    11'b01101111010: data <= 32'hae2d205d;
    11'b01101111011: data <= 32'hb4db3714;
    11'b01101111100: data <= 32'hb2c0bafb;
    11'b01101111101: data <= 32'h3997c12b;
    11'b01101111110: data <= 32'h3d97c0c4;
    11'b01101111111: data <= 32'h3925b630;
    11'b01110000000: data <= 32'hbad13c67;
    11'b01110000001: data <= 32'hbd053af2;
    11'b01110000010: data <= 32'hb7772b05;
    11'b01110000011: data <= 32'hb54dae36;
    11'b01110000100: data <= 32'hbe691ddf;
    11'b01110000101: data <= 32'hc0e2b590;
    11'b01110000110: data <= 32'hbc54b851;
    11'b01110000111: data <= 32'h3d423486;
    11'b01110001000: data <= 32'h403d3d9f;
    11'b01110001001: data <= 32'h3aca3dc6;
    11'b01110001010: data <= 32'hb741391b;
    11'b01110001011: data <= 32'hb5903853;
    11'b01110001100: data <= 32'h34e83d44;
    11'b01110001101: data <= 32'h35083cb6;
    11'b01110001110: data <= 32'h2f69ba07;
    11'b01110001111: data <= 32'h391cc134;
    11'b01110010000: data <= 32'h3d8dc04b;
    11'b01110010001: data <= 32'h3cd9a98c;
    11'b01110010010: data <= 32'h357e3c44;
    11'b01110010011: data <= 32'h210b3364;
    11'b01110010100: data <= 32'h325cbad5;
    11'b01110010101: data <= 32'hb6ecb9c3;
    11'b01110010110: data <= 32'hc010b047;
    11'b01110010111: data <= 32'hc15bb5db;
    11'b01110011000: data <= 32'hbc60bbc8;
    11'b01110011001: data <= 32'h3c63b984;
    11'b01110011010: data <= 32'h3d7b35cf;
    11'b01110011011: data <= 32'hb2893be9;
    11'b01110011100: data <= 32'hbcea3c0c;
    11'b01110011101: data <= 32'hb83d3d73;
    11'b01110011110: data <= 32'h36e63ffb;
    11'b01110011111: data <= 32'h31a73e09;
    11'b01110100000: data <= 32'hb814b715;
    11'b01110100001: data <= 32'hadacbfa9;
    11'b01110100010: data <= 32'h3ccdbca4;
    11'b01110100011: data <= 32'h3f6439a7;
    11'b01110100100: data <= 32'h3ddb3ca6;
    11'b01110100101: data <= 32'h3befb0cd;
    11'b01110100110: data <= 32'h39bebc79;
    11'b01110100111: data <= 32'hb0fdb812;
    11'b01110101000: data <= 32'hbe4b3475;
    11'b01110101001: data <= 32'hbfdcb637;
    11'b01110101010: data <= 32'hb85dbf17;
    11'b01110101011: data <= 32'h3c13bfdf;
    11'b01110101100: data <= 32'h39b7b9ef;
    11'b01110101101: data <= 32'hbafe376a;
    11'b01110101110: data <= 32'hbdb13b55;
    11'b01110101111: data <= 32'hb5ee3d05;
    11'b01110110000: data <= 32'h355d3eba;
    11'b01110110001: data <= 32'hb8e23d1a;
    11'b01110110010: data <= 32'hbf14b0df;
    11'b01110110011: data <= 32'hbc97bc30;
    11'b01110110100: data <= 32'h3a9eb264;
    11'b01110110101: data <= 32'h401e3cce;
    11'b01110110110: data <= 32'h3f203c99;
    11'b01110110111: data <= 32'h3c6fb054;
    11'b01110111000: data <= 32'h3a74b860;
    11'b01110111001: data <= 32'h34f33853;
    11'b01110111010: data <= 32'hb8e53ca5;
    11'b01110111011: data <= 32'hbb2cb3e1;
    11'b01110111100: data <= 32'h2c28c0ad;
    11'b01110111101: data <= 32'h3c0bc16e;
    11'b01110111110: data <= 32'h382ebcf2;
    11'b01110111111: data <= 32'hb95b30e1;
    11'b01111000000: data <= 32'hb9e4366d;
    11'b01111000001: data <= 32'h340535a4;
    11'b01111000010: data <= 32'h34233993;
    11'b01111000011: data <= 32'hbdd839f8;
    11'b01111000100: data <= 32'hc1b99bba;
    11'b01111000101: data <= 32'hbfaab88e;
    11'b01111000110: data <= 32'h371c2448;
    11'b01111000111: data <= 32'h3eb43b7a;
    11'b01111001000: data <= 32'h3c733a76;
    11'b01111001001: data <= 32'h35d12d67;
    11'b01111001010: data <= 32'h37eb36dc;
    11'b01111001011: data <= 32'h39913f38;
    11'b01111001100: data <= 32'h31b6401c;
    11'b01111001101: data <= 32'hb4c52c45;
    11'b01111001110: data <= 32'h30ffc07f;
    11'b01111001111: data <= 32'h3b0ac0e2;
    11'b01111010000: data <= 32'h3a27babb;
    11'b01111010001: data <= 32'h33ba3273;
    11'b01111010010: data <= 32'h37afb301;
    11'b01111010011: data <= 32'h3c64b99b;
    11'b01111010100: data <= 32'h3658b1bd;
    11'b01111010101: data <= 32'hbf013711;
    11'b01111010110: data <= 32'hc2252c41;
    11'b01111010111: data <= 32'hbfaeb995;
    11'b01111011000: data <= 32'h343db94f;
    11'b01111011001: data <= 32'h3b74aa24;
    11'b01111011010: data <= 32'hac0d3115;
    11'b01111011011: data <= 32'hb92331d0;
    11'b01111011100: data <= 32'h30823c53;
    11'b01111011101: data <= 32'h3b0640ee;
    11'b01111011110: data <= 32'h352240d9;
    11'b01111011111: data <= 32'hb907363a;
    11'b01111100000: data <= 32'hb7e7be32;
    11'b01111100001: data <= 32'h37f8bd68;
    11'b01111100010: data <= 32'h3c682f3a;
    11'b01111100011: data <= 32'h3cab3778;
    11'b01111100100: data <= 32'h3dd0b90e;
    11'b01111100101: data <= 32'h3ed1bce1;
    11'b01111100110: data <= 32'h39ecb439;
    11'b01111100111: data <= 32'hbd063a09;
    11'b01111101000: data <= 32'hc08b3330;
    11'b01111101001: data <= 32'hbcccbcb9;
    11'b01111101010: data <= 32'h357ebee6;
    11'b01111101011: data <= 32'h3426bc98;
    11'b01111101100: data <= 32'hbbb8b7fc;
    11'b01111101101: data <= 32'hbc86a8c2;
    11'b01111101110: data <= 32'h31b43b4f;
    11'b01111101111: data <= 32'h3b85402c;
    11'b01111110000: data <= 32'hb0c2401f;
    11'b01111110001: data <= 32'hbe9c385f;
    11'b01111110010: data <= 32'hbe30b964;
    11'b01111110011: data <= 32'ha956b1bd;
    11'b01111110100: data <= 32'h3c8d3b30;
    11'b01111110101: data <= 32'h3d9638c7;
    11'b01111110110: data <= 32'h3e1cb9ff;
    11'b01111110111: data <= 32'h3edabbaf;
    11'b01111111000: data <= 32'h3c6e3848;
    11'b01111111001: data <= 32'hb49d3e7d;
    11'b01111111010: data <= 32'hbc0e3871;
    11'b01111111011: data <= 32'hb4e3be1d;
    11'b01111111100: data <= 32'h37f7c0b7;
    11'b01111111101: data <= 32'ha8e5be7d;
    11'b01111111110: data <= 32'hbc41ba48;
    11'b01111111111: data <= 32'hb9adb800;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    