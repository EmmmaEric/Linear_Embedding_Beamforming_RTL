
module memory_rom_14(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hb3d73e46;
    11'b00000000001: data <= 32'hadef3aaf;
    11'b00000000010: data <= 32'h32d8bbc0;
    11'b00000000011: data <= 32'h3c99bded;
    11'b00000000100: data <= 32'h3ee332e9;
    11'b00000000101: data <= 32'h3cd84011;
    11'b00000000110: data <= 32'h38043ee4;
    11'b00000000111: data <= 32'h387aae77;
    11'b00000001000: data <= 32'h3978bcb0;
    11'b00000001001: data <= 32'hb345bb3e;
    11'b00000001010: data <= 32'hbd91b9bc;
    11'b00000001011: data <= 32'hbba7bd57;
    11'b00000001100: data <= 32'h3bbbbebd;
    11'b00000001101: data <= 32'h3fbdbb4d;
    11'b00000001110: data <= 32'h38173070;
    11'b00000001111: data <= 32'hbe7e36ba;
    11'b00000010000: data <= 32'hc02235e7;
    11'b00000010001: data <= 32'hbbe53a83;
    11'b00000010010: data <= 32'hb6ab3c97;
    11'b00000010011: data <= 32'hbbc333d7;
    11'b00000010100: data <= 32'hbc9dbcc5;
    11'b00000010101: data <= 32'ha814bc5d;
    11'b00000010110: data <= 32'h3d0b3b2d;
    11'b00000010111: data <= 32'h3da040fb;
    11'b00000011000: data <= 32'h3a8c3f66;
    11'b00000011001: data <= 32'h386e3026;
    11'b00000011010: data <= 32'h3706b623;
    11'b00000011011: data <= 32'hb36c3574;
    11'b00000011100: data <= 32'hbab03576;
    11'b00000011101: data <= 32'haafdbc3b;
    11'b00000011110: data <= 32'h3ebdc05e;
    11'b00000011111: data <= 32'h406dbe88;
    11'b00000100000: data <= 32'h3946b44f;
    11'b00000100001: data <= 32'hbc70359d;
    11'b00000100010: data <= 32'hbc8732d9;
    11'b00000100011: data <= 32'hb1bd32b4;
    11'b00000100100: data <= 32'hb60a32c0;
    11'b00000100101: data <= 32'hbf20b840;
    11'b00000100110: data <= 32'hc083bddd;
    11'b00000100111: data <= 32'hba47bc2c;
    11'b00000101000: data <= 32'h3bfa3a31;
    11'b00000101001: data <= 32'h3cf33ff7;
    11'b00000101010: data <= 32'h35293d7b;
    11'b00000101011: data <= 32'hb3af34e0;
    11'b00000101100: data <= 32'hb2a6391b;
    11'b00000101101: data <= 32'hb59c3ed2;
    11'b00000101110: data <= 32'hb8293d43;
    11'b00000101111: data <= 32'h336bb9fb;
    11'b00000110000: data <= 32'h3e87c05b;
    11'b00000110001: data <= 32'h401dbdb0;
    11'b00000110010: data <= 32'h3bc5339b;
    11'b00000110011: data <= 32'ha9ea3a0c;
    11'b00000110100: data <= 32'h34a72e85;
    11'b00000110101: data <= 32'h3ac9b635;
    11'b00000110110: data <= 32'hb0e8b6ce;
    11'b00000110111: data <= 32'hc026ba9e;
    11'b00000111000: data <= 32'hc0f0be1f;
    11'b00000111001: data <= 32'hb94cbd7d;
    11'b00000111010: data <= 32'h3c8bb0f0;
    11'b00000111011: data <= 32'h3b6f39d2;
    11'b00000111100: data <= 32'hb7b83792;
    11'b00000111101: data <= 32'hbc703448;
    11'b00000111110: data <= 32'hb98d3d1d;
    11'b00000111111: data <= 32'hb77640c4;
    11'b00001000000: data <= 32'hb9b23e6b;
    11'b00001000001: data <= 32'hb69eb949;
    11'b00001000010: data <= 32'h3980bf33;
    11'b00001000011: data <= 32'h3db8b89a;
    11'b00001000100: data <= 32'h3cb63cb4;
    11'b00001000101: data <= 32'h3b373d16;
    11'b00001000110: data <= 32'h3d6c2ebf;
    11'b00001000111: data <= 32'h3de8b7ac;
    11'b00001001000: data <= 32'h2c5cb15e;
    11'b00001001001: data <= 32'hbf21b446;
    11'b00001001010: data <= 32'hbf2abcd5;
    11'b00001001011: data <= 32'h30d7bf39;
    11'b00001001100: data <= 32'h3e2fbd3d;
    11'b00001001101: data <= 32'h39d0b87d;
    11'b00001001110: data <= 32'hbb7bb54f;
    11'b00001001111: data <= 32'hbd2429dc;
    11'b00001010000: data <= 32'hb8083cd9;
    11'b00001010001: data <= 32'hb60c401a;
    11'b00001010010: data <= 32'hbd0d3c5d;
    11'b00001010011: data <= 32'hbe86baef;
    11'b00001010100: data <= 32'hb91ebd88;
    11'b00001010101: data <= 32'h39253277;
    11'b00001010110: data <= 32'h3c6f3ef7;
    11'b00001010111: data <= 32'h3caa3d83;
    11'b00001011000: data <= 32'h3dd82f69;
    11'b00001011001: data <= 32'h3d6a2024;
    11'b00001011010: data <= 32'h2ed33b6b;
    11'b00001011011: data <= 32'hbcdb3b71;
    11'b00001011100: data <= 32'hba9fb8bc;
    11'b00001011101: data <= 32'h3badc003;
    11'b00001011110: data <= 32'h3f4abfd7;
    11'b00001011111: data <= 32'h3990bc69;
    11'b00001100000: data <= 32'hb988b892;
    11'b00001100001: data <= 32'hb7f9b205;
    11'b00001100010: data <= 32'h36e238cf;
    11'b00001100011: data <= 32'h124d3c59;
    11'b00001100100: data <= 32'hbf0733ec;
    11'b00001100101: data <= 32'hc14cbc9b;
    11'b00001100110: data <= 32'hbe2dbcca;
    11'b00001100111: data <= 32'h311d3510;
    11'b00001101000: data <= 32'h3a8a3d8c;
    11'b00001101001: data <= 32'h394a3a50;
    11'b00001101010: data <= 32'h3964a8b0;
    11'b00001101011: data <= 32'h395b39a7;
    11'b00001101100: data <= 32'ha7894064;
    11'b00001101101: data <= 32'hba604024;
    11'b00001101110: data <= 32'hb563a497;
    11'b00001101111: data <= 32'h3c34bf57;
    11'b00001110000: data <= 32'h3e54beec;
    11'b00001110001: data <= 32'h399eb913;
    11'b00001110010: data <= 32'h2a8eb169;
    11'b00001110011: data <= 32'h3a94b4a1;
    11'b00001110100: data <= 32'h3e89ac4f;
    11'b00001110101: data <= 32'h3832347a;
    11'b00001110110: data <= 32'hbf60b216;
    11'b00001110111: data <= 32'hc1aabca4;
    11'b00001111000: data <= 32'hbdf9bd01;
    11'b00001111001: data <= 32'h33f6b4cf;
    11'b00001111010: data <= 32'h3801336d;
    11'b00001111011: data <= 32'hb233b499;
    11'b00001111100: data <= 32'hb553b667;
    11'b00001111101: data <= 32'h2a3d3c6d;
    11'b00001111110: data <= 32'hafa041ad;
    11'b00001111111: data <= 32'hba0540ed;
    11'b00010000000: data <= 32'hb97d316a;
    11'b00010000001: data <= 32'h3327bdac;
    11'b00010000010: data <= 32'h3a3fbac6;
    11'b00010000011: data <= 32'h38883684;
    11'b00010000100: data <= 32'h39dd3778;
    11'b00010000101: data <= 32'h3f63b49f;
    11'b00010000110: data <= 32'h40ccb5b1;
    11'b00010000111: data <= 32'h3b31342b;
    11'b00010001000: data <= 32'hbde933be;
    11'b00010001001: data <= 32'hc03fb977;
    11'b00010001010: data <= 32'hb8e1bd5d;
    11'b00010001011: data <= 32'h3a0cbcb0;
    11'b00010001100: data <= 32'h34eabc0c;
    11'b00010001101: data <= 32'hba76bd0a;
    11'b00010001110: data <= 32'hba1aba9f;
    11'b00010001111: data <= 32'h2e693b72;
    11'b00010010000: data <= 32'h2e3740f6;
    11'b00010010001: data <= 32'hbbc63fac;
    11'b00010010010: data <= 32'hbe6fae82;
    11'b00010010011: data <= 32'hbc35bc0d;
    11'b00010010100: data <= 32'hb24b2c06;
    11'b00010010101: data <= 32'h33cd3cd0;
    11'b00010010110: data <= 32'h3acf39c1;
    11'b00010010111: data <= 32'h3fbcb602;
    11'b00010011000: data <= 32'h4092b1a2;
    11'b00010011001: data <= 32'h3b4e3c3c;
    11'b00010011010: data <= 32'hbb503d82;
    11'b00010011011: data <= 32'hbc353056;
    11'b00010011100: data <= 32'h3680bd00;
    11'b00010011101: data <= 32'h3cbcbe91;
    11'b00010011110: data <= 32'h32b2be29;
    11'b00010011111: data <= 32'hbac1be39;
    11'b00010100000: data <= 32'hb44bbc59;
    11'b00010100001: data <= 32'h3bad34ec;
    11'b00010100010: data <= 32'h396c3db8;
    11'b00010100011: data <= 32'hbc983b23;
    11'b00010100100: data <= 32'hc0d5b84d;
    11'b00010100101: data <= 32'hbfc9ba4b;
    11'b00010100110: data <= 32'hba4236df;
    11'b00010100111: data <= 32'hb02b3c8c;
    11'b00010101000: data <= 32'h34f53315;
    11'b00010101001: data <= 32'h3c4fb9bf;
    11'b00010101010: data <= 32'h3dd03233;
    11'b00010101011: data <= 32'h39164031;
    11'b00010101100: data <= 32'hb7a54104;
    11'b00010101101: data <= 32'hb55f3ad2;
    11'b00010101110: data <= 32'h3a40bb82;
    11'b00010101111: data <= 32'h3c35bd62;
    11'b00010110000: data <= 32'h29c7bc15;
    11'b00010110001: data <= 32'hb6e4bc2f;
    11'b00010110010: data <= 32'h3a75bc48;
    11'b00010110011: data <= 32'h404fb5dd;
    11'b00010110100: data <= 32'h3d8336c7;
    11'b00010110101: data <= 32'hbc2d31b0;
    11'b00010110110: data <= 32'hc102b96b;
    11'b00010110111: data <= 32'hbf71b992;
    11'b00010111000: data <= 32'hb9123051;
    11'b00010111001: data <= 32'hb5d533a2;
    11'b00010111010: data <= 32'hb862babd;
    11'b00010111011: data <= 32'hae83bd20;
    11'b00010111100: data <= 32'h388b35c1;
    11'b00010111101: data <= 32'h3659413b;
    11'b00010111110: data <= 32'hb51c41c4;
    11'b00010111111: data <= 32'hb5ff3c20;
    11'b00011000000: data <= 32'h3315b875;
    11'b00011000001: data <= 32'h346ab734;
    11'b00011000010: data <= 32'hb4da316c;
    11'b00011000011: data <= 32'ha427b14e;
    11'b00011000100: data <= 32'h3ebebb46;
    11'b00011000101: data <= 32'h41d6b9e8;
    11'b00011000110: data <= 32'h3f2f2f1e;
    11'b00011000111: data <= 32'hb9503548;
    11'b00011001000: data <= 32'hbf14b3d9;
    11'b00011001001: data <= 32'hbad0b896;
    11'b00011001010: data <= 32'h2dc1b71d;
    11'b00011001011: data <= 32'hb662bab9;
    11'b00011001100: data <= 32'hbce2bf51;
    11'b00011001101: data <= 32'hba72bf37;
    11'b00011001110: data <= 32'h354a2f8e;
    11'b00011001111: data <= 32'h3854406f;
    11'b00011010000: data <= 32'hb5694078;
    11'b00011010001: data <= 32'hbbec38a3;
    11'b00011010010: data <= 32'hbaf3b4c6;
    11'b00011010011: data <= 32'hb9cf3806;
    11'b00011010100: data <= 32'hba223ce2;
    11'b00011010101: data <= 32'ha3a93618;
    11'b00011010110: data <= 32'h3edbbb2c;
    11'b00011010111: data <= 32'h4176b9e7;
    11'b00011011000: data <= 32'h3eb138c6;
    11'b00011011001: data <= 32'hb3183d0a;
    11'b00011011010: data <= 32'hb94938ca;
    11'b00011011011: data <= 32'h3670b4e1;
    11'b00011011100: data <= 32'h3a81ba00;
    11'b00011011101: data <= 32'hb5f8bd2c;
    11'b00011011110: data <= 32'hbda6c02a;
    11'b00011011111: data <= 32'hb8fdbfeb;
    11'b00011100000: data <= 32'h3bb7b6ac;
    11'b00011100001: data <= 32'h3c8c3c85;
    11'b00011100010: data <= 32'hb50b3bef;
    11'b00011100011: data <= 32'hbe60b0aa;
    11'b00011100100: data <= 32'hbeb0b2da;
    11'b00011100101: data <= 32'hbd333c01;
    11'b00011100110: data <= 32'hbc763ddb;
    11'b00011100111: data <= 32'hb815301c;
    11'b00011101000: data <= 32'h3a95bcf2;
    11'b00011101001: data <= 32'h3ed2b89e;
    11'b00011101010: data <= 32'h3c7c3d99;
    11'b00011101011: data <= 32'h2bf54091;
    11'b00011101100: data <= 32'h31563d52;
    11'b00011101101: data <= 32'h3c56291b;
    11'b00011101110: data <= 32'h3b95b740;
    11'b00011101111: data <= 32'hb815b9e3;
    11'b00011110000: data <= 32'hbcd3bda5;
    11'b00011110001: data <= 32'h323bbedd;
    11'b00011110010: data <= 32'h4011bb83;
    11'b00011110011: data <= 32'h3f7b27a3;
    11'b00011110100: data <= 32'hb007a66e;
    11'b00011110101: data <= 32'hbe88b895;
    11'b00011110110: data <= 32'hbe2bb1b8;
    11'b00011110111: data <= 32'hbc1a3b40;
    11'b00011111000: data <= 32'hbc943ab8;
    11'b00011111001: data <= 32'hbce9ba55;
    11'b00011111010: data <= 32'hb6ffbf5f;
    11'b00011111011: data <= 32'h3834b84d;
    11'b00011111100: data <= 32'h389f3f4f;
    11'b00011111101: data <= 32'h305b4137;
    11'b00011111110: data <= 32'h350c3db0;
    11'b00011111111: data <= 32'h3a853446;
    11'b00100000000: data <= 32'h3569353a;
    11'b00100000001: data <= 32'hbb393835;
    11'b00100000010: data <= 32'hbb9bb406;
    11'b00100000011: data <= 32'h3b90bcf9;
    11'b00100000100: data <= 32'h417dbccd;
    11'b00100000101: data <= 32'h407ab748;
    11'b00100000110: data <= 32'h30fdb1b7;
    11'b00100000111: data <= 32'hbbd9b564;
    11'b00100001000: data <= 32'hb77da569;
    11'b00100001001: data <= 32'ha9d93811;
    11'b00100001010: data <= 32'hbafcad00;
    11'b00100001011: data <= 32'hbf17bee1;
    11'b00100001100: data <= 32'hbd31c0b4;
    11'b00100001101: data <= 32'ha7b8b9e6;
    11'b00100001110: data <= 32'h37e33de7;
    11'b00100001111: data <= 32'h30313f9a;
    11'b00100010000: data <= 32'haeb839f0;
    11'b00100010001: data <= 32'had5a33a6;
    11'b00100010010: data <= 32'hb8c43c95;
    11'b00100010011: data <= 32'hbd8c3ee2;
    11'b00100010100: data <= 32'hbbb038f7;
    11'b00100010101: data <= 32'h3be4bbc1;
    11'b00100010110: data <= 32'h4101bcbe;
    11'b00100010111: data <= 32'h3fb3b168;
    11'b00100011000: data <= 32'h3578383e;
    11'b00100011001: data <= 32'h98a436c0;
    11'b00100011010: data <= 32'h3b5b34a4;
    11'b00100011011: data <= 32'h3c053438;
    11'b00100011100: data <= 32'hb87bb815;
    11'b00100011101: data <= 32'hbfafbfb8;
    11'b00100011110: data <= 32'hbd41c0c2;
    11'b00100011111: data <= 32'h35afbc39;
    11'b00100100000: data <= 32'h3bd3380e;
    11'b00100100001: data <= 32'h329d3841;
    11'b00100100010: data <= 32'hb8dab4ef;
    11'b00100100011: data <= 32'hbaa924dc;
    11'b00100100100: data <= 32'hbc8b3e4e;
    11'b00100100101: data <= 32'hbe8a4051;
    11'b00100100110: data <= 32'hbd263923;
    11'b00100100111: data <= 32'h3246bcab;
    11'b00100101000: data <= 32'h3d75bc4b;
    11'b00100101001: data <= 32'h3c3d3802;
    11'b00100101010: data <= 32'h35033dde;
    11'b00100101011: data <= 32'h39ec3c7f;
    11'b00100101100: data <= 32'h3f2c38a6;
    11'b00100101101: data <= 32'h3dc23721;
    11'b00100101110: data <= 32'hb82aa83e;
    11'b00100101111: data <= 32'hbf02bca4;
    11'b00100110000: data <= 32'hb932bf4e;
    11'b00100110001: data <= 32'h3d3abd13;
    11'b00100110010: data <= 32'h3eb7b7f2;
    11'b00100110011: data <= 32'h361bb967;
    11'b00100110100: data <= 32'hb9a8bc3c;
    11'b00100110101: data <= 32'hba12b117;
    11'b00100110110: data <= 32'hba443e01;
    11'b00100110111: data <= 32'hbda43ed1;
    11'b00100111000: data <= 32'hbedcb018;
    11'b00100111001: data <= 32'hbbb1beed;
    11'b00100111010: data <= 32'h95b3bc32;
    11'b00100111011: data <= 32'h31813b89;
    11'b00100111100: data <= 32'h306e3f4a;
    11'b00100111101: data <= 32'h3b1b3ca0;
    11'b00100111110: data <= 32'h3ed638ca;
    11'b00100111111: data <= 32'h3c0e3bba;
    11'b00101000000: data <= 32'hbad43c82;
    11'b00101000001: data <= 32'hbe1f31a0;
    11'b00101000010: data <= 32'h2cc2bc00;
    11'b00101000011: data <= 32'h400cbd01;
    11'b00101000100: data <= 32'h4004bbaf;
    11'b00101000101: data <= 32'h3803bc1c;
    11'b00101000110: data <= 32'hb466bc2e;
    11'b00101000111: data <= 32'h3314ad9e;
    11'b00101001000: data <= 32'h35c33c96;
    11'b00101001001: data <= 32'hba4d3ac8;
    11'b00101001010: data <= 32'hbfd9bc29;
    11'b00101001011: data <= 32'hbf21c06f;
    11'b00101001100: data <= 32'hba22bc89;
    11'b00101001101: data <= 32'hb1983a23;
    11'b00101001110: data <= 32'h21f03ccb;
    11'b00101001111: data <= 32'h3818354f;
    11'b00101010000: data <= 32'h3b3a3391;
    11'b00101010001: data <= 32'h2fd13dee;
    11'b00101010010: data <= 32'hbd4c4089;
    11'b00101010011: data <= 32'hbde13d10;
    11'b00101010100: data <= 32'h33feb6d1;
    11'b00101010101: data <= 32'h3f6dbc4c;
    11'b00101010110: data <= 32'h3e48b9b0;
    11'b00101010111: data <= 32'h3617b711;
    11'b00101011000: data <= 32'h368db5c7;
    11'b00101011001: data <= 32'h3e3232c8;
    11'b00101011010: data <= 32'h3e883af5;
    11'b00101011011: data <= 32'hb09e3528;
    11'b00101011100: data <= 32'hbfa3bd43;
    11'b00101011101: data <= 32'hbf4ac04c;
    11'b00101011110: data <= 32'hb841bcba;
    11'b00101011111: data <= 32'h32402cd6;
    11'b00101100000: data <= 32'h2c24aee3;
    11'b00101100001: data <= 32'h2006bb87;
    11'b00101100010: data <= 32'h2e83b55d;
    11'b00101100011: data <= 32'hb7953eb8;
    11'b00101100100: data <= 32'hbe06416f;
    11'b00101100101: data <= 32'hbe473dd9;
    11'b00101100110: data <= 32'hb499b770;
    11'b00101100111: data <= 32'h3a42bb57;
    11'b00101101000: data <= 32'h37d3ab51;
    11'b00101101001: data <= 32'ha1333814;
    11'b00101101010: data <= 32'h3b29361e;
    11'b00101101011: data <= 32'h40d93772;
    11'b00101101100: data <= 32'h40883afa;
    11'b00101101101: data <= 32'h2e6a389a;
    11'b00101101110: data <= 32'hbea7b8eb;
    11'b00101101111: data <= 32'hbcbcbd94;
    11'b00101110000: data <= 32'h3661bc23;
    11'b00101110001: data <= 32'h3b55b940;
    11'b00101110010: data <= 32'h331cbd3e;
    11'b00101110011: data <= 32'hb338bfa9;
    11'b00101110100: data <= 32'ha43aba1b;
    11'b00101110101: data <= 32'hb2393df9;
    11'b00101110110: data <= 32'hbc6e4096;
    11'b00101110111: data <= 32'hbe9b39fb;
    11'b00101111000: data <= 32'hbcacbc15;
    11'b00101111001: data <= 32'hb898bb13;
    11'b00101111010: data <= 32'hb92137a0;
    11'b00101111011: data <= 32'hb7a33c18;
    11'b00101111100: data <= 32'h3b2e37dd;
    11'b00101111101: data <= 32'h40be357b;
    11'b00101111110: data <= 32'h3fba3c4d;
    11'b00101111111: data <= 32'hb20c3dd9;
    11'b00110000000: data <= 32'hbdb939a4;
    11'b00110000001: data <= 32'hb660b508;
    11'b00110000010: data <= 32'h3cf7b983;
    11'b00110000011: data <= 32'h3d4abb89;
    11'b00110000100: data <= 32'h3391bec8;
    11'b00110000101: data <= 32'haca6c00f;
    11'b00110000110: data <= 32'h399dba3a;
    11'b00110000111: data <= 32'h3b643c78;
    11'b00110001000: data <= 32'hb36c3d99;
    11'b00110001001: data <= 32'hbe2fb425;
    11'b00110001010: data <= 32'hbf21be53;
    11'b00110001011: data <= 32'hbd7fbb29;
    11'b00110001100: data <= 32'hbca13853;
    11'b00110001101: data <= 32'hb9ec3927;
    11'b00110001110: data <= 32'h37aeb4c4;
    11'b00110001111: data <= 32'h3e33b42e;
    11'b00110010000: data <= 32'h3bd33ced;
    11'b00110010001: data <= 32'hb9cd40c0;
    11'b00110010010: data <= 32'hbd4b3f51;
    11'b00110010011: data <= 32'ha5cb3779;
    11'b00110010100: data <= 32'h3d34b528;
    11'b00110010101: data <= 32'h3b74b8ff;
    11'b00110010110: data <= 32'haeb2bc73;
    11'b00110010111: data <= 32'h341bbd4a;
    11'b00110011000: data <= 32'h3f2ab6e2;
    11'b00110011001: data <= 32'h40753a80;
    11'b00110011010: data <= 32'h393239ae;
    11'b00110011011: data <= 32'hbd03b9f3;
    11'b00110011100: data <= 32'hbee5be4c;
    11'b00110011101: data <= 32'hbca0ba02;
    11'b00110011110: data <= 32'hba773209;
    11'b00110011111: data <= 32'hb95ab6b7;
    11'b00110100000: data <= 32'ha94bbe67;
    11'b00110100001: data <= 32'h38f1bc5f;
    11'b00110100010: data <= 32'h32253c96;
    11'b00110100011: data <= 32'hbbe14165;
    11'b00110100100: data <= 32'hbd0f401d;
    11'b00110100101: data <= 32'hb3c337f2;
    11'b00110100110: data <= 32'h3782b08c;
    11'b00110100111: data <= 32'hb1892a24;
    11'b00110101000: data <= 32'hba22abd0;
    11'b00110101001: data <= 32'h36e0b69a;
    11'b00110101010: data <= 32'h4107ada6;
    11'b00110101011: data <= 32'h41d0398c;
    11'b00110101100: data <= 32'h3c0a3961;
    11'b00110101101: data <= 32'hbb7cb492;
    11'b00110101110: data <= 32'hbc37ba7a;
    11'b00110101111: data <= 32'hb0e5b551;
    11'b00110110000: data <= 32'h2a39b2be;
    11'b00110110001: data <= 32'hb6bbbdd0;
    11'b00110110010: data <= 32'hb5d0c143;
    11'b00110110011: data <= 32'h33acbebc;
    11'b00110110100: data <= 32'h335b3ab5;
    11'b00110110101: data <= 32'hb8c54073;
    11'b00110110110: data <= 32'hbc5a3d2c;
    11'b00110110111: data <= 32'hba3eb116;
    11'b00110111000: data <= 32'hb9a0b213;
    11'b00110111001: data <= 32'hbd7b3929;
    11'b00110111010: data <= 32'hbdc33973;
    11'b00110111011: data <= 32'h342aac3b;
    11'b00110111100: data <= 32'h40cab1a9;
    11'b00110111101: data <= 32'h4118394c;
    11'b00110111110: data <= 32'h39503cde;
    11'b00110111111: data <= 32'hba193ab3;
    11'b00111000000: data <= 32'hb30c357d;
    11'b00111000001: data <= 32'h3b1c341c;
    11'b00111000010: data <= 32'h3978b475;
    11'b00111000011: data <= 32'hb594bf05;
    11'b00111000100: data <= 32'hb69ec17f;
    11'b00111000101: data <= 32'h3901bec3;
    11'b00111000110: data <= 32'h3c8f37d8;
    11'b00111000111: data <= 32'h358f3d27;
    11'b00111001000: data <= 32'hb9b72f45;
    11'b00111001001: data <= 32'hbc8cbb7c;
    11'b00111001010: data <= 32'hbd9db46d;
    11'b00111001011: data <= 32'hbfad3b0a;
    11'b00111001100: data <= 32'hbf0138f1;
    11'b00111001101: data <= 32'hb163b918;
    11'b00111001110: data <= 32'h3e21baac;
    11'b00111001111: data <= 32'h3dca3852;
    11'b00111010000: data <= 32'hac863f60;
    11'b00111010001: data <= 32'hb9f03f63;
    11'b00111010010: data <= 32'h34c13cbc;
    11'b00111010011: data <= 32'h3cfd39d2;
    11'b00111010100: data <= 32'h382c2e24;
    11'b00111010101: data <= 32'hb9c8bc82;
    11'b00111010110: data <= 32'hb5bcbfb5;
    11'b00111010111: data <= 32'h3da3bcaf;
    11'b00111011000: data <= 32'h40a2346b;
    11'b00111011001: data <= 32'h3d3c37b5;
    11'b00111011010: data <= 32'hb436b93a;
    11'b00111011011: data <= 32'hbbc8bcaa;
    11'b00111011100: data <= 32'hbc8aaffa;
    11'b00111011101: data <= 32'hbdf63a4f;
    11'b00111011110: data <= 32'hbe30b033;
    11'b00111011111: data <= 32'hb8dcbf30;
    11'b00111100000: data <= 32'h3805bf08;
    11'b00111100001: data <= 32'h365a340b;
    11'b00111100010: data <= 32'hb89b4007;
    11'b00111100011: data <= 32'hb99f4008;
    11'b00111100100: data <= 32'h35193cb0;
    11'b00111100101: data <= 32'h39e03a9b;
    11'b00111100110: data <= 32'hb6d439a9;
    11'b00111100111: data <= 32'hbdec1e0c;
    11'b00111101000: data <= 32'hb6bdba30;
    11'b00111101001: data <= 32'h3fc5b8a4;
    11'b00111101010: data <= 32'h41da327c;
    11'b00111101011: data <= 32'h3eab333b;
    11'b00111101100: data <= 32'h276db821;
    11'b00111101101: data <= 32'hb552b89b;
    11'b00111101110: data <= 32'habbc362c;
    11'b00111101111: data <= 32'hb6ae392c;
    11'b00111110000: data <= 32'hbc3abb8d;
    11'b00111110001: data <= 32'hbae5c183;
    11'b00111110010: data <= 32'hac69c0c4;
    11'b00111110011: data <= 32'h2f4badb1;
    11'b00111110100: data <= 32'hb6223e20;
    11'b00111110101: data <= 32'hb7323cbe;
    11'b00111110110: data <= 32'h2a4b3552;
    11'b00111110111: data <= 32'hb2223872;
    11'b00111111000: data <= 32'hbe313ce7;
    11'b00111111001: data <= 32'hc0723b59;
    11'b00111111010: data <= 32'hb96eaf05;
    11'b00111111011: data <= 32'h3f19b72f;
    11'b00111111100: data <= 32'h41032fb7;
    11'b00111111101: data <= 32'h3cb13803;
    11'b00111111110: data <= 32'h2222356e;
    11'b00111111111: data <= 32'h36c737dc;
    11'b01000000000: data <= 32'h3c873c46;
    11'b01000000001: data <= 32'h383839be;
    11'b01000000010: data <= 32'hb9f4bca5;
    11'b01000000011: data <= 32'hbb78c1a3;
    11'b01000000100: data <= 32'h2b33c091;
    11'b01000000101: data <= 32'h39e6b49d;
    11'b01000000110: data <= 32'h3754394b;
    11'b01000000111: data <= 32'h284cb025;
    11'b01000001000: data <= 32'haff9b9ef;
    11'b01000001001: data <= 32'hba3032ea;
    11'b01000001010: data <= 32'hc0193dd0;
    11'b01000001011: data <= 32'hc0f23c68;
    11'b01000001100: data <= 32'hbc08b612;
    11'b01000001101: data <= 32'h3bacbbd9;
    11'b01000001110: data <= 32'h3d22af48;
    11'b01000001111: data <= 32'h310a3b4b;
    11'b01000010000: data <= 32'hb3303cca;
    11'b01000010001: data <= 32'h3b4b3d2a;
    11'b01000010010: data <= 32'h3ee53e1f;
    11'b01000010011: data <= 32'h396d3c32;
    11'b01000010100: data <= 32'hbbbbb874;
    11'b01000010101: data <= 32'hbbd8bf8d;
    11'b01000010110: data <= 32'h38d0be09;
    11'b01000010111: data <= 32'h3eefb407;
    11'b01000011000: data <= 32'h3d86ae79;
    11'b01000011001: data <= 32'h3829bc77;
    11'b01000011010: data <= 32'h2af0bd30;
    11'b01000011011: data <= 32'hb80431ff;
    11'b01000011100: data <= 32'hbe1f3dc8;
    11'b01000011101: data <= 32'hc01938d0;
    11'b01000011110: data <= 32'hbcdcbd55;
    11'b01000011111: data <= 32'ha4cabf72;
    11'b01000100000: data <= 32'h2606b78f;
    11'b01000100001: data <= 32'hb9733c0c;
    11'b01000100010: data <= 32'hb64e3d57;
    11'b01000100011: data <= 32'h3bf63cd6;
    11'b01000100100: data <= 32'h3ddb3dd2;
    11'b01000100101: data <= 32'ha9143dd6;
    11'b01000100110: data <= 32'hbeae3831;
    11'b01000100111: data <= 32'hbc8db84f;
    11'b01000101000: data <= 32'h3c15b8a5;
    11'b01000101001: data <= 32'h4092add9;
    11'b01000101010: data <= 32'h3ebfb655;
    11'b01000101011: data <= 32'h3987bcf2;
    11'b01000101100: data <= 32'h384cbbb1;
    11'b01000101101: data <= 32'h383938ff;
    11'b01000101110: data <= 32'hb4713da5;
    11'b01000101111: data <= 32'hbcebaba2;
    11'b01000110000: data <= 32'hbcdfc06a;
    11'b01000110001: data <= 32'hb8dbc0e6;
    11'b01000110010: data <= 32'hb824b9f5;
    11'b01000110011: data <= 32'hba2d391b;
    11'b01000110100: data <= 32'hb3b0384b;
    11'b01000110101: data <= 32'h3ab132b4;
    11'b01000110110: data <= 32'h39c03afd;
    11'b01000110111: data <= 32'hbc353ee2;
    11'b01000111000: data <= 32'hc0c73dbd;
    11'b01000111001: data <= 32'hbd80361f;
    11'b01000111010: data <= 32'h3b48b071;
    11'b01000111011: data <= 32'h3f85a943;
    11'b01000111100: data <= 32'h3c38b334;
    11'b01000111101: data <= 32'h364eb8b1;
    11'b01000111110: data <= 32'h3c2fa738;
    11'b01000111111: data <= 32'h3ed43d2c;
    11'b01001000000: data <= 32'h3b5d3e06;
    11'b01001000001: data <= 32'hb8aab496;
    11'b01001000010: data <= 32'hbc7cc08b;
    11'b01001000011: data <= 32'hb895c07b;
    11'b01001000100: data <= 32'hafbab9a3;
    11'b01001000101: data <= 32'hae089e35;
    11'b01001000110: data <= 32'h333dba17;
    11'b01001000111: data <= 32'h39c7bc72;
    11'b01001001000: data <= 32'h317d31ec;
    11'b01001001001: data <= 32'hbe2b3eff;
    11'b01001001010: data <= 32'hc11d3ec4;
    11'b01001001011: data <= 32'hbe0d35b3;
    11'b01001001100: data <= 32'h34a4b78d;
    11'b01001001101: data <= 32'h3964b3d2;
    11'b01001001110: data <= 32'hb2482e74;
    11'b01001001111: data <= 32'hb246324a;
    11'b01001010000: data <= 32'h3d3f39f7;
    11'b01001010001: data <= 32'h40b63ed0;
    11'b01001010010: data <= 32'h3d503eca;
    11'b01001010011: data <= 32'hb88d310b;
    11'b01001010100: data <= 32'hbc73bd6c;
    11'b01001010101: data <= 32'haff9bcfb;
    11'b01001010110: data <= 32'h3a1bb521;
    11'b01001010111: data <= 32'h3a44b846;
    11'b01001011000: data <= 32'h3980bf2c;
    11'b01001011001: data <= 32'h3a84bfbe;
    11'b01001011010: data <= 32'h3526af62;
    11'b01001011011: data <= 32'hbc263e9e;
    11'b01001011100: data <= 32'hbfc23d2a;
    11'b01001011101: data <= 32'hbd90b743;
    11'b01001011110: data <= 32'hb736bd22;
    11'b01001011111: data <= 32'hb8fbb8c1;
    11'b01001100000: data <= 32'hbd43339d;
    11'b01001100001: data <= 32'hb95e369e;
    11'b01001100010: data <= 32'h3d1a396c;
    11'b01001100011: data <= 32'h40633ddd;
    11'b01001100100: data <= 32'h3a443f3e;
    11'b01001100101: data <= 32'hbcb33c08;
    11'b01001100110: data <= 32'hbd102608;
    11'b01001100111: data <= 32'h34a4a795;
    11'b01001101000: data <= 32'h3d6a3197;
    11'b01001101001: data <= 32'h3c68b96e;
    11'b01001101010: data <= 32'h39e0c003;
    11'b01001101011: data <= 32'h3c2cbf35;
    11'b01001101100: data <= 32'h3c8d3213;
    11'b01001101101: data <= 32'h339c3e71;
    11'b01001101110: data <= 32'hbaaa3950;
    11'b01001101111: data <= 32'hbc27bd52;
    11'b01001110000: data <= 32'hbae5bf85;
    11'b01001110001: data <= 32'hbd05ba3d;
    11'b01001110010: data <= 32'hbe8d2c61;
    11'b01001110011: data <= 32'hb984b243;
    11'b01001110100: data <= 32'h3c5fb562;
    11'b01001110101: data <= 32'h3e0438e8;
    11'b01001110110: data <= 32'hb2573ed7;
    11'b01001110111: data <= 32'hbf933ee2;
    11'b01001111000: data <= 32'hbdcc3c20;
    11'b01001111001: data <= 32'h355d3964;
    11'b01001111010: data <= 32'h3c703710;
    11'b01001111011: data <= 32'h376bb767;
    11'b01001111100: data <= 32'h3214bdb8;
    11'b01001111101: data <= 32'h3cccbb79;
    11'b01001111110: data <= 32'h40373ac3;
    11'b01001111111: data <= 32'h3e123eb5;
    11'b01010000000: data <= 32'h2e66353d;
    11'b01010000001: data <= 32'hb970be1b;
    11'b01010000010: data <= 32'hba08beb0;
    11'b01010000011: data <= 32'hbb8db82f;
    11'b01010000100: data <= 32'hbc41b3d7;
    11'b01010000101: data <= 32'hb420bd23;
    11'b01010000110: data <= 32'h3bbebeef;
    11'b01010000111: data <= 32'h3b1bb612;
    11'b01010001000: data <= 32'hba593dbf;
    11'b01010001001: data <= 32'hc0263f7f;
    11'b01010001010: data <= 32'hbda03c67;
    11'b01010001011: data <= 32'h237037c4;
    11'b01010001100: data <= 32'h2ec534e6;
    11'b01010001101: data <= 32'hbadfb039;
    11'b01010001110: data <= 32'hb9b1b8ec;
    11'b01010001111: data <= 32'h3c8bad42;
    11'b01010010000: data <= 32'h41413d1c;
    11'b01010010001: data <= 32'h400e3eea;
    11'b01010010010: data <= 32'h34ce3812;
    11'b01010010011: data <= 32'hb87bba6c;
    11'b01010010100: data <= 32'hb4bab8eb;
    11'b01010010101: data <= 32'hab9d316c;
    11'b01010010110: data <= 32'hb073b6d9;
    11'b01010010111: data <= 32'h336dc056;
    11'b01010011000: data <= 32'h3bafc156;
    11'b01010011001: data <= 32'h3a87bb40;
    11'b01010011010: data <= 32'hb7853cbd;
    11'b01010011011: data <= 32'hbda33dcb;
    11'b01010011100: data <= 32'hbbea3510;
    11'b01010011101: data <= 32'hb604b566;
    11'b01010011110: data <= 32'hbc1fac54;
    11'b01010011111: data <= 32'hc0302c7b;
    11'b01010100000: data <= 32'hbdcdb2f5;
    11'b01010100001: data <= 32'h3b2c24bd;
    11'b01010100010: data <= 32'h40d73c0e;
    11'b01010100011: data <= 32'h3e1f3e4a;
    11'b01010100100: data <= 32'hb46f3c10;
    11'b01010100101: data <= 32'hb9c73688;
    11'b01010100110: data <= 32'h311d39c7;
    11'b01010100111: data <= 32'h39603bae;
    11'b01010101000: data <= 32'h3551b53b;
    11'b01010101001: data <= 32'h3463c0a2;
    11'b01010101010: data <= 32'h3ba6c134;
    11'b01010101011: data <= 32'h3d39b962;
    11'b01010101100: data <= 32'h390f3c7e;
    11'b01010101101: data <= 32'hb1dd3a5a;
    11'b01010101110: data <= 32'hb518b952;
    11'b01010101111: data <= 32'hb80abc46;
    11'b01010110000: data <= 32'hbe53b44b;
    11'b01010110001: data <= 32'hc1042df7;
    11'b01010110010: data <= 32'hbe59b834;
    11'b01010110011: data <= 32'h3949ba8f;
    11'b01010110100: data <= 32'h3ed42a9a;
    11'b01010110101: data <= 32'h379b3c93;
    11'b01010110110: data <= 32'hbc6e3dad;
    11'b01010110111: data <= 32'hbb783d48;
    11'b01010111000: data <= 32'h35bc3e2a;
    11'b01010111001: data <= 32'h39943d97;
    11'b01010111010: data <= 32'hb024a436;
    11'b01010111011: data <= 32'hb5c8bedc;
    11'b01010111100: data <= 32'h3a50bec4;
    11'b01010111101: data <= 32'h3fcc2c56;
    11'b01010111110: data <= 32'h3f363ce5;
    11'b01010111111: data <= 32'h3b133567;
    11'b01011000000: data <= 32'h342dbc67;
    11'b01011000001: data <= 32'hb41fbc24;
    11'b01011000010: data <= 32'hbcf62b2f;
    11'b01011000011: data <= 32'hbfb22d57;
    11'b01011000100: data <= 32'hbc6cbd23;
    11'b01011000101: data <= 32'h3887c031;
    11'b01011000110: data <= 32'h3bffbc5a;
    11'b01011000111: data <= 32'hb54c38d7;
    11'b01011001000: data <= 32'hbddb3d8c;
    11'b01011001001: data <= 32'hbacb3d67;
    11'b01011001010: data <= 32'h35083d82;
    11'b01011001011: data <= 32'h248d3d06;
    11'b01011001100: data <= 32'hbd4b34c4;
    11'b01011001101: data <= 32'hbda9baa4;
    11'b01011001110: data <= 32'h36d9b941;
    11'b01011001111: data <= 32'h407c3960;
    11'b01011010000: data <= 32'h40883d09;
    11'b01011010001: data <= 32'h3c953460;
    11'b01011010010: data <= 32'h36d9b986;
    11'b01011010011: data <= 32'h32c1af64;
    11'b01011010100: data <= 32'hb4d13b2e;
    11'b01011010101: data <= 32'hbac732f9;
    11'b01011010110: data <= 32'hb73ebfa6;
    11'b01011010111: data <= 32'h388cc1f3;
    11'b01011011000: data <= 32'h39b8bed7;
    11'b01011011001: data <= 32'hb4ec33fa;
    11'b01011011010: data <= 32'hbb903b51;
    11'b01011011011: data <= 32'hb4b9382a;
    11'b01011011100: data <= 32'h33f436fe;
    11'b01011011101: data <= 32'hbabc39e8;
    11'b01011011110: data <= 32'hc0fe3793;
    11'b01011011111: data <= 32'hc08eb40d;
    11'b01011100000: data <= 32'h2796b456;
    11'b01011100001: data <= 32'h3fcc388e;
    11'b01011100010: data <= 32'h3ee73be8;
    11'b01011100011: data <= 32'h37d03759;
    11'b01011100100: data <= 32'h30e0335f;
    11'b01011100101: data <= 32'h39133c9e;
    11'b01011100110: data <= 32'h38a23f5c;
    11'b01011100111: data <= 32'haef73838;
    11'b01011101000: data <= 32'hb37fbfbf;
    11'b01011101001: data <= 32'h37a5c1be;
    11'b01011101010: data <= 32'h3b2ebdbf;
    11'b01011101011: data <= 32'h37ec342a;
    11'b01011101100: data <= 32'h328d348d;
    11'b01011101101: data <= 32'h385db8af;
    11'b01011101110: data <= 32'h35f0b851;
    11'b01011101111: data <= 32'hbcef35a2;
    11'b01011110000: data <= 32'hc1c13867;
    11'b01011110001: data <= 32'hc0d7b46e;
    11'b01011110010: data <= 32'hb1c7ba71;
    11'b01011110011: data <= 32'h3cfab4d6;
    11'b01011110100: data <= 32'h38823621;
    11'b01011110101: data <= 32'hb882389e;
    11'b01011110110: data <= 32'hb3db3b9e;
    11'b01011110111: data <= 32'h3ade3fc8;
    11'b01011111000: data <= 32'h3ae840a7;
    11'b01011111001: data <= 32'hb4403aef;
    11'b01011111010: data <= 32'hba16bd46;
    11'b01011111011: data <= 32'h308abf79;
    11'b01011111100: data <= 32'h3cf1b806;
    11'b01011111101: data <= 32'h3dcb3850;
    11'b01011111110: data <= 32'h3cffb1a7;
    11'b01011111111: data <= 32'h3ce2bd05;
    11'b01100000000: data <= 32'h39a2ba79;
    11'b01100000001: data <= 32'hbaca385d;
    11'b01100000010: data <= 32'hc06f3988;
    11'b01100000011: data <= 32'hbf1fb9c9;
    11'b01100000100: data <= 32'haf5abf60;
    11'b01100000101: data <= 32'h3858bdac;
    11'b01100000110: data <= 32'hb743b4a4;
    11'b01100000111: data <= 32'hbcdf3674;
    11'b01100001000: data <= 32'hb5033b48;
    11'b01100001001: data <= 32'h3b863ee6;
    11'b01100001010: data <= 32'h37e34025;
    11'b01100001011: data <= 32'hbcd13c33;
    11'b01100001100: data <= 32'hbf22b71d;
    11'b01100001101: data <= 32'hb61db923;
    11'b01100001110: data <= 32'h3d5a364f;
    11'b01100001111: data <= 32'h3f3c39fa;
    11'b01100010000: data <= 32'h3de3b572;
    11'b01100010001: data <= 32'h3d4ebc94;
    11'b01100010010: data <= 32'h3c55b109;
    11'b01100010011: data <= 32'h2d563d61;
    11'b01100010100: data <= 32'hbbc43c03;
    11'b01100010101: data <= 32'hbac4bc7c;
    11'b01100010110: data <= 32'h2cc1c12f;
    11'b01100010111: data <= 32'h31f0c009;
    11'b01100011000: data <= 32'hb9c4b91c;
    11'b01100011001: data <= 32'hbbdba7d3;
    11'b01100011010: data <= 32'h31c42cc9;
    11'b01100011011: data <= 32'h3c39391a;
    11'b01100011100: data <= 32'haf013d2d;
    11'b01100011101: data <= 32'hc0733c21;
    11'b01100011110: data <= 32'hc14731cd;
    11'b01100011111: data <= 32'hba9925bc;
    11'b01100100000: data <= 32'h3c1d38b6;
    11'b01100100001: data <= 32'h3cfc387c;
    11'b01100100010: data <= 32'h3988b547;
    11'b01100100011: data <= 32'h3a96b801;
    11'b01100100100: data <= 32'h3d483b86;
    11'b01100100101: data <= 32'h3bf44094;
    11'b01100100110: data <= 32'h28333d9d;
    11'b01100100111: data <= 32'hb511bc4e;
    11'b01100101000: data <= 32'h2e4ec0e4;
    11'b01100101001: data <= 32'h32a3be96;
    11'b01100101010: data <= 32'hb2a4b716;
    11'b01100101011: data <= 32'ha659b7f1;
    11'b01100101100: data <= 32'h3c1cbc35;
    11'b01100101101: data <= 32'h3d3bb8b4;
    11'b01100101110: data <= 32'hb62a38b8;
    11'b01100101111: data <= 32'hc1183bb8;
    11'b01100110000: data <= 32'hc16b34be;
    11'b01100110001: data <= 32'hbb33b2dd;
    11'b01100110010: data <= 32'h3744ac3b;
    11'b01100110011: data <= 32'h2c2fa9d2;
    11'b01100110100: data <= 32'hb8bcb5ec;
    11'b01100110101: data <= 32'h2ef72c18;
    11'b01100110110: data <= 32'h3d823ea1;
    11'b01100110111: data <= 32'h3d924179;
    11'b01100111000: data <= 32'h31a63ea6;
    11'b01100111001: data <= 32'hb8ccb867;
    11'b01100111010: data <= 32'hb316bdaf;
    11'b01100111011: data <= 32'h35f1b803;
    11'b01100111100: data <= 32'h386c3086;
    11'b01100111101: data <= 32'h3b70ba38;
    11'b01100111110: data <= 32'h3ec4bf43;
    11'b01100111111: data <= 32'h3e77bca1;
    11'b01101000000: data <= 32'haa51381c;
    11'b01101000001: data <= 32'hbf713c41;
    11'b01101000010: data <= 32'hbf892758;
    11'b01101000011: data <= 32'hb867bc1e;
    11'b01101000100: data <= 32'hac24bc4b;
    11'b01101000101: data <= 32'hbc20b9d6;
    11'b01101000110: data <= 32'hbe2fb898;
    11'b01101000111: data <= 32'hb40a2673;
    11'b01101001000: data <= 32'h3d8d3da0;
    11'b01101001001: data <= 32'h3cc740a7;
    11'b01101001010: data <= 32'hb8223e60;
    11'b01101001011: data <= 32'hbdf630cc;
    11'b01101001100: data <= 32'hba26b005;
    11'b01101001101: data <= 32'h3652398a;
    11'b01101001110: data <= 32'h3af8394d;
    11'b01101001111: data <= 32'h3c7abab7;
    11'b01101010000: data <= 32'h3eb8bf78;
    11'b01101010001: data <= 32'h3f29ba2a;
    11'b01101010010: data <= 32'h39d23c9e;
    11'b01101010011: data <= 32'hb86c3d99;
    11'b01101010100: data <= 32'hb945b414;
    11'b01101010101: data <= 32'ha842bec7;
    11'b01101010110: data <= 32'hb4b8be89;
    11'b01101010111: data <= 32'hbdccbc02;
    11'b01101011000: data <= 32'hbe5dbada;
    11'b01101011001: data <= 32'h2ae1b975;
    11'b01101011010: data <= 32'h3e123441;
    11'b01101011011: data <= 32'h39d93d18;
    11'b01101011100: data <= 32'hbdad3cfa;
    11'b01101011101: data <= 32'hc0993905;
    11'b01101011110: data <= 32'hbcb0396e;
    11'b01101011111: data <= 32'h31c53cbf;
    11'b01101100000: data <= 32'h36703994;
    11'b01101100001: data <= 32'h34acba9b;
    11'b01101100010: data <= 32'h3b6ebd81;
    11'b01101100011: data <= 32'h3ed331ab;
    11'b01101100100: data <= 32'h3de94015;
    11'b01101100101: data <= 32'h38a43f2a;
    11'b01101100110: data <= 32'h31f3b405;
    11'b01101100111: data <= 32'h33ecbe6c;
    11'b01101101000: data <= 32'hb3ddbce3;
    11'b01101101001: data <= 32'hbc65b8bc;
    11'b01101101010: data <= 32'hba83bc1b;
    11'b01101101011: data <= 32'h3aa2be96;
    11'b01101101100: data <= 32'h3f22bc51;
    11'b01101101101: data <= 32'h376533ca;
    11'b01101101110: data <= 32'hbf0d3b18;
    11'b01101101111: data <= 32'hc0ac397f;
    11'b01101110000: data <= 32'hbc4a38e1;
    11'b01101110001: data <= 32'hb05339f3;
    11'b01101110010: data <= 32'hb90231f2;
    11'b01101110011: data <= 32'hbc68bb27;
    11'b01101110100: data <= 32'haf45bae1;
    11'b01101110101: data <= 32'h3dc93b15;
    11'b01101110110: data <= 32'h3f2b40ed;
    11'b01101110111: data <= 32'h3b233fac;
    11'b01101111000: data <= 32'h30b72bbd;
    11'b01101111001: data <= 32'h2b05b9bc;
    11'b01101111010: data <= 32'haf242622;
    11'b01101111011: data <= 32'hb6bf3500;
    11'b01101111100: data <= 32'h2e72bbd3;
    11'b01101111101: data <= 32'h3de5c09b;
    11'b01101111110: data <= 32'h4002bf43;
    11'b01101111111: data <= 32'h390daef1;
    11'b01110000000: data <= 32'hbcc53a8e;
    11'b01110000001: data <= 32'hbdae3705;
    11'b01110000010: data <= 32'hb6b7ae18;
    11'b01110000011: data <= 32'hb532b21a;
    11'b01110000100: data <= 32'hbe69b7af;
    11'b01110000101: data <= 32'hc071bc35;
    11'b01110000110: data <= 32'hba3aba41;
    11'b01110000111: data <= 32'h3cff39d9;
    11'b01110001000: data <= 32'h3e613fec;
    11'b01110001001: data <= 32'h35473e4c;
    11'b01110001010: data <= 32'hb9163717;
    11'b01110001011: data <= 32'hb772373e;
    11'b01110001100: data <= 32'hacce3d89;
    11'b01110001101: data <= 32'ha86e3ca4;
    11'b01110001110: data <= 32'h35d6ba5c;
    11'b01110001111: data <= 32'h3da3c0ab;
    11'b01110010000: data <= 32'h3fc3be4c;
    11'b01110010001: data <= 32'h3c733632;
    11'b01110010010: data <= 32'ha1b13c6f;
    11'b01110010011: data <= 32'ha83a313f;
    11'b01110010100: data <= 32'h370fba46;
    11'b01110010101: data <= 32'hb46fba6d;
    11'b01110010110: data <= 32'hbfebb9c3;
    11'b01110010111: data <= 32'hc0dabc91;
    11'b01110011000: data <= 32'hb940bce7;
    11'b01110011001: data <= 32'h3d37b493;
    11'b01110011010: data <= 32'h3c993a30;
    11'b01110011011: data <= 32'hb87a3afe;
    11'b01110011100: data <= 32'hbde238f2;
    11'b01110011101: data <= 32'hbad33ccd;
    11'b01110011110: data <= 32'hb0aa401b;
    11'b01110011111: data <= 32'hb47b3dae;
    11'b01110100000: data <= 32'hb581b95f;
    11'b01110100001: data <= 32'h382abf73;
    11'b01110100010: data <= 32'h3e0cb95d;
    11'b01110100011: data <= 32'h3e303d18;
    11'b01110100100: data <= 32'h3c343dfa;
    11'b01110100101: data <= 32'h3c012c4b;
    11'b01110100110: data <= 32'h3beabb03;
    11'b01110100111: data <= 32'had0db802;
    11'b01110101000: data <= 32'hbe92b240;
    11'b01110101001: data <= 32'hbee4bbeb;
    11'b01110101010: data <= 32'h2da0bf7e;
    11'b01110101011: data <= 32'h3e43be32;
    11'b01110101100: data <= 32'h3a88b74e;
    11'b01110101101: data <= 32'hbc2d32b3;
    11'b01110101110: data <= 32'hbe6f37cc;
    11'b01110101111: data <= 32'hb94f3c8b;
    11'b01110110000: data <= 32'hb1833ed9;
    11'b01110110001: data <= 32'hbc033bd2;
    11'b01110110010: data <= 32'hbe99b9d1;
    11'b01110110011: data <= 32'hb9cbbd3e;
    11'b01110110100: data <= 32'h3b543088;
    11'b01110110101: data <= 32'h3e873f24;
    11'b01110110110: data <= 32'h3d6d3e3a;
    11'b01110110111: data <= 32'h3c623022;
    11'b01110111000: data <= 32'h3b48b458;
    11'b01110111001: data <= 32'h2d8b393b;
    11'b01110111010: data <= 32'hbb9c3b41;
    11'b01110111011: data <= 32'hb9e8b8b5;
    11'b01110111100: data <= 32'h3a7fc08a;
    11'b01110111101: data <= 32'h3effc089;
    11'b01110111110: data <= 32'h3a39bbc2;
    11'b01110111111: data <= 32'hb9dea5b8;
    11'b01111000000: data <= 32'hba4831b1;
    11'b01111000001: data <= 32'h319636dd;
    11'b01111000010: data <= 32'h9d3139f5;
    11'b01111000011: data <= 32'hbece33f2;
    11'b01111000100: data <= 32'hc17cbaf7;
    11'b01111000101: data <= 32'hbe4ebc43;
    11'b01111000110: data <= 32'h3807330a;
    11'b01111000111: data <= 32'h3d583d9a;
    11'b01111001000: data <= 32'h3a633c30;
    11'b01111001001: data <= 32'h350f313e;
    11'b01111001010: data <= 32'h35a738e1;
    11'b01111001011: data <= 32'h2ff13fec;
    11'b01111001100: data <= 32'hb7023fdb;
    11'b01111001101: data <= 32'hb44fb099;
    11'b01111001110: data <= 32'h3ad2c054;
    11'b01111001111: data <= 32'h3e2fc010;
    11'b01111010000: data <= 32'h3b72b820;
    11'b01111010001: data <= 32'h311b3446;
    11'b01111010010: data <= 32'h3884ae3a;
    11'b01111010011: data <= 32'h3d0ab5a1;
    11'b01111010100: data <= 32'h357ba97d;
    11'b01111010101: data <= 32'hbf9fae8c;
    11'b01111010110: data <= 32'hc1e8bad9;
    11'b01111010111: data <= 32'hbe23bcd8;
    11'b01111011000: data <= 32'h381db81a;
    11'b01111011001: data <= 32'h3b0633a1;
    11'b01111011010: data <= 32'hb1082f61;
    11'b01111011011: data <= 32'hb94d20a1;
    11'b01111011100: data <= 32'hb0a23c9f;
    11'b01111011101: data <= 32'h2ff04151;
    11'b01111011110: data <= 32'hb6b940af;
    11'b01111011111: data <= 32'hb9a12ca8;
    11'b01111100000: data <= 32'h253ebea2;
    11'b01111100001: data <= 32'h3b21bc53;
    11'b01111100010: data <= 32'h3c1037b6;
    11'b01111100011: data <= 32'h3bf83a0a;
    11'b01111100100: data <= 32'h3e71b395;
    11'b01111100101: data <= 32'h3fe0b95b;
    11'b01111100110: data <= 32'h397e977c;
    11'b01111100111: data <= 32'hbe09359c;
    11'b01111101000: data <= 32'hc06fb7e8;
    11'b01111101001: data <= 32'hb9b5be05;
    11'b01111101010: data <= 32'h3ae4be22;
    11'b01111101011: data <= 32'h382abc04;
    11'b01111101100: data <= 32'hbaa8b9fa;
    11'b01111101101: data <= 32'hbc2db522;
    11'b01111101110: data <= 32'ha9963c03;
    11'b01111101111: data <= 32'h347b409a;
    11'b01111110000: data <= 32'hba653f75;
    11'b01111110001: data <= 32'hbf04a967;
    11'b01111110010: data <= 32'hbcefbc5d;
    11'b01111110011: data <= 32'h2c5eaeea;
    11'b01111110100: data <= 32'h3ad43ce2;
    11'b01111110101: data <= 32'h3cbc3b5e;
    11'b01111110110: data <= 32'h3ed2b536;
    11'b01111110111: data <= 32'h3f9bb63c;
    11'b01111111000: data <= 32'h3aa23b26;
    11'b01111111001: data <= 32'hba6c3dd0;
    11'b01111111010: data <= 32'hbc6530d1;
    11'b01111111011: data <= 32'h330abe76;
    11'b01111111100: data <= 32'h3ca3c036;
    11'b01111111101: data <= 32'h35cfbe21;
    11'b01111111110: data <= 32'hba96bc2b;
    11'b01111111111: data <= 32'hb7b7b93c;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    