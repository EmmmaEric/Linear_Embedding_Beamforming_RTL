
module memory_rom_15(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h2e763e56;
    11'b00000000001: data <= 32'h2dde3ab5;
    11'b00000000010: data <= 32'h98babbea;
    11'b00000000011: data <= 32'h3a63bec9;
    11'b00000000100: data <= 32'h3ee8b159;
    11'b00000000101: data <= 32'h3e803ee2;
    11'b00000000110: data <= 32'h3aec3e4c;
    11'b00000000111: data <= 32'h3832b2f5;
    11'b00000001000: data <= 32'h369bbd2b;
    11'b00000001001: data <= 32'hb6aabaaf;
    11'b00000001010: data <= 32'hbe0eb65a;
    11'b00000001011: data <= 32'hbce7bc5f;
    11'b00000001100: data <= 32'h3897bf6b;
    11'b00000001101: data <= 32'h3ec2bd41;
    11'b00000001110: data <= 32'h384225b1;
    11'b00000001111: data <= 32'hbdf63a1a;
    11'b00000010000: data <= 32'hbfc13a7a;
    11'b00000010001: data <= 32'hba4e3c08;
    11'b00000010010: data <= 32'hb1073cd8;
    11'b00000010011: data <= 32'hbb23373c;
    11'b00000010100: data <= 32'hbd8bbb4a;
    11'b00000010101: data <= 32'hb456bc3d;
    11'b00000010110: data <= 32'h3db238c9;
    11'b00000010111: data <= 32'h3fa9403f;
    11'b00000011000: data <= 32'h3ccf3e85;
    11'b00000011001: data <= 32'h388d2048;
    11'b00000011010: data <= 32'h3587b787;
    11'b00000011011: data <= 32'hb0d6361b;
    11'b00000011100: data <= 32'hb9ee3821;
    11'b00000011101: data <= 32'hb490bc12;
    11'b00000011110: data <= 32'h3cabc0fe;
    11'b00000011111: data <= 32'h3f3ac028;
    11'b00000100000: data <= 32'h38b4b68b;
    11'b00000100001: data <= 32'hbc0538aa;
    11'b00000100010: data <= 32'hbc3c3749;
    11'b00000100011: data <= 32'hb02d33cb;
    11'b00000100100: data <= 32'hb522349c;
    11'b00000100101: data <= 32'hbf68b02b;
    11'b00000100110: data <= 32'hc10bbb84;
    11'b00000100111: data <= 32'hbbf9bacc;
    11'b00000101000: data <= 32'h3c8e384a;
    11'b00000101001: data <= 32'h3e913eb2;
    11'b00000101010: data <= 32'h38eb3d13;
    11'b00000101011: data <= 32'hb15e359b;
    11'b00000101100: data <= 32'hac203955;
    11'b00000101101: data <= 32'h27533ef5;
    11'b00000101110: data <= 32'hb3163d99;
    11'b00000101111: data <= 32'h2bffba36;
    11'b00000110000: data <= 32'h3c79c0f6;
    11'b00000110001: data <= 32'h3eccbf5a;
    11'b00000110010: data <= 32'h3c0124ad;
    11'b00000110011: data <= 32'h2fad39fc;
    11'b00000110100: data <= 32'h34e128d2;
    11'b00000110101: data <= 32'h39f3b881;
    11'b00000110110: data <= 32'hb3a8b61e;
    11'b00000110111: data <= 32'hc068b5b1;
    11'b00000111000: data <= 32'hc17dbba6;
    11'b00000111001: data <= 32'hbb97bcc8;
    11'b00000111010: data <= 32'h3c4bb663;
    11'b00000111011: data <= 32'h3c44380f;
    11'b00000111100: data <= 32'hb5da3889;
    11'b00000111101: data <= 32'hbc1a3804;
    11'b00000111110: data <= 32'hb6693d96;
    11'b00000111111: data <= 32'h2c0340da;
    11'b00001000000: data <= 32'hb5863ee6;
    11'b00001000001: data <= 32'hb862b869;
    11'b00001000010: data <= 32'h3472bf9f;
    11'b00001000011: data <= 32'h3d14bb00;
    11'b00001000100: data <= 32'h3d9f3b1f;
    11'b00001000101: data <= 32'h3ca03c30;
    11'b00001000110: data <= 32'h3d61b213;
    11'b00001000111: data <= 32'h3d5aba51;
    11'b00001001000: data <= 32'h283bb1c1;
    11'b00001001001: data <= 32'hbf2f3013;
    11'b00001001010: data <= 32'hc006ba4e;
    11'b00001001011: data <= 32'hb3f1bf2d;
    11'b00001001100: data <= 32'h3ce5be77;
    11'b00001001101: data <= 32'h38b7b9a8;
    11'b00001001110: data <= 32'hbbddafc4;
    11'b00001001111: data <= 32'hbcfc352b;
    11'b00001010000: data <= 32'hb35a3d2a;
    11'b00001010001: data <= 32'h2cf9402b;
    11'b00001010010: data <= 32'hbbf13d5e;
    11'b00001010011: data <= 32'hbf1fb7d1;
    11'b00001010100: data <= 32'hbb6bbcd9;
    11'b00001010101: data <= 32'h395b2afc;
    11'b00001010110: data <= 32'h3dd73dd4;
    11'b00001010111: data <= 32'h3dc03c5f;
    11'b00001011000: data <= 32'h3dceb280;
    11'b00001011001: data <= 32'h3d4bb49a;
    11'b00001011010: data <= 32'h34ed3b0b;
    11'b00001011011: data <= 32'hbbdb3cb1;
    11'b00001011100: data <= 32'hbb82b64f;
    11'b00001011101: data <= 32'h37f7c055;
    11'b00001011110: data <= 32'h3d69c09f;
    11'b00001011111: data <= 32'h3710bcea;
    11'b00001100000: data <= 32'hba63b688;
    11'b00001100001: data <= 32'hb83bacdc;
    11'b00001100010: data <= 32'h386537e0;
    11'b00001100011: data <= 32'h33a83c3e;
    11'b00001100100: data <= 32'hbea23900;
    11'b00001100101: data <= 32'hc1abb860;
    11'b00001100110: data <= 32'hbf15baab;
    11'b00001100111: data <= 32'h331b345a;
    11'b00001101000: data <= 32'h3c653cb4;
    11'b00001101001: data <= 32'h3a8a3907;
    11'b00001101010: data <= 32'h3932b1d2;
    11'b00001101011: data <= 32'h3a753855;
    11'b00001101100: data <= 32'h3732404b;
    11'b00001101101: data <= 32'hb53a4064;
    11'b00001101110: data <= 32'hb5562ba9;
    11'b00001101111: data <= 32'h3901c009;
    11'b00001110000: data <= 32'h3cacc011;
    11'b00001110001: data <= 32'h3864ba31;
    11'b00001110010: data <= 32'h22b8b1a3;
    11'b00001110011: data <= 32'h39e7b75f;
    11'b00001110100: data <= 32'h3e52b6bf;
    11'b00001110101: data <= 32'h389c3110;
    11'b00001110110: data <= 32'hbf5932e9;
    11'b00001110111: data <= 32'hc209b820;
    11'b00001111000: data <= 32'hbeeebb2d;
    11'b00001111001: data <= 32'h319db594;
    11'b00001111010: data <= 32'h38512f88;
    11'b00001111011: data <= 32'hb401b39a;
    11'b00001111100: data <= 32'hb699b51b;
    11'b00001111101: data <= 32'h34973c43;
    11'b00001111110: data <= 32'h38024196;
    11'b00001111111: data <= 32'hb2524124;
    11'b00010000000: data <= 32'hb9103517;
    11'b00010000001: data <= 32'hadd8bdb9;
    11'b00010000010: data <= 32'h389ebbfc;
    11'b00010000011: data <= 32'h3922345e;
    11'b00010000100: data <= 32'h3a8734c2;
    11'b00010000101: data <= 32'h3ef4b975;
    11'b00010000110: data <= 32'h4087baf5;
    11'b00010000111: data <= 32'h3b812b56;
    11'b00010001000: data <= 32'hbd8c3876;
    11'b00010001001: data <= 32'hc072b283;
    11'b00010001010: data <= 32'hbb1fbcb4;
    11'b00010001011: data <= 32'h37b7bd3c;
    11'b00010001100: data <= 32'h2d3abc38;
    11'b00010001101: data <= 32'hbc3ebc37;
    11'b00010001110: data <= 32'hbb68b926;
    11'b00010001111: data <= 32'h34c63b12;
    11'b00010010000: data <= 32'h391540cd;
    11'b00010010001: data <= 32'hb83c402b;
    11'b00010010010: data <= 32'hbe5e340d;
    11'b00010010011: data <= 32'hbcfeba15;
    11'b00010010100: data <= 32'hb1c12e86;
    11'b00010010101: data <= 32'h37fb3c7c;
    11'b00010010110: data <= 32'h3be43827;
    11'b00010010111: data <= 32'h3f38ba49;
    11'b00010011000: data <= 32'h4063b95d;
    11'b00010011001: data <= 32'h3c7f3aaa;
    11'b00010011010: data <= 32'hb8ba3e2c;
    11'b00010011011: data <= 32'hbbfc35d2;
    11'b00010011100: data <= 32'h2fd9bd3a;
    11'b00010011101: data <= 32'h3a64bf70;
    11'b00010011110: data <= 32'hb01cbe33;
    11'b00010011111: data <= 32'hbca5bd57;
    11'b00010100000: data <= 32'hb801bc04;
    11'b00010100001: data <= 32'h3c012dbc;
    11'b00010100010: data <= 32'h3bcb3cfd;
    11'b00010100011: data <= 32'hbb643c7c;
    11'b00010100100: data <= 32'hc0f3180c;
    11'b00010100101: data <= 32'hc025b587;
    11'b00010100110: data <= 32'hb96138b3;
    11'b00010100111: data <= 32'h2fa63c8e;
    11'b00010101000: data <= 32'h359a30d4;
    11'b00010101001: data <= 32'h3b27bb7b;
    11'b00010101010: data <= 32'h3dd8b027;
    11'b00010101011: data <= 32'h3c503fa0;
    11'b00010101100: data <= 32'h2d27411b;
    11'b00010101101: data <= 32'hb0943b45;
    11'b00010101110: data <= 32'h3875bc55;
    11'b00010101111: data <= 32'h39e2be2c;
    11'b00010110000: data <= 32'hb1a4bc07;
    11'b00010110001: data <= 32'hb930bb6b;
    11'b00010110010: data <= 32'h386bbce1;
    11'b00010110011: data <= 32'h400bba9f;
    11'b00010110100: data <= 32'h3dc22f38;
    11'b00010110101: data <= 32'hbbd0366a;
    11'b00010110110: data <= 32'hc12eaf6c;
    11'b00010110111: data <= 32'hbfe1b46a;
    11'b00010111000: data <= 32'hb8ba344c;
    11'b00010111001: data <= 32'hb4db3502;
    11'b00010111010: data <= 32'hb9beb99c;
    11'b00010111011: data <= 32'hb612bceb;
    11'b00010111100: data <= 32'h390d332a;
    11'b00010111101: data <= 32'h3ba640ed;
    11'b00010111110: data <= 32'h350f41c5;
    11'b00010111111: data <= 32'hb0873c5e;
    11'b00011000000: data <= 32'h2e08b8ba;
    11'b00011000001: data <= 32'h3180b801;
    11'b00011000010: data <= 32'hb4233363;
    11'b00011000011: data <= 32'haad4b103;
    11'b00011000100: data <= 32'h3dc8bd03;
    11'b00011000101: data <= 32'h4160bd6d;
    11'b00011000110: data <= 32'h3f1fb48a;
    11'b00011000111: data <= 32'hb8963776;
    11'b00011001000: data <= 32'hbf1f30ad;
    11'b00011001001: data <= 32'hbba9b5fb;
    11'b00011001010: data <= 32'ha0c4b742;
    11'b00011001011: data <= 32'hb88fb9dc;
    11'b00011001100: data <= 32'hbe5bbe14;
    11'b00011001101: data <= 32'hbcb9be59;
    11'b00011001110: data <= 32'h358a2919;
    11'b00011001111: data <= 32'h3c0a4016;
    11'b00011010000: data <= 32'h310d4083;
    11'b00011010001: data <= 32'hbab83a44;
    11'b00011010010: data <= 32'hbb4eae90;
    11'b00011010011: data <= 32'hb8cc392d;
    11'b00011010100: data <= 32'hb7bc3d6f;
    11'b00011010101: data <= 32'h2c42360b;
    11'b00011010110: data <= 32'h3de7bcfb;
    11'b00011010111: data <= 32'h4102bd43;
    11'b00011011000: data <= 32'h3f1032eb;
    11'b00011011001: data <= 32'h2ba63d1c;
    11'b00011011010: data <= 32'hb81f39d7;
    11'b00011011011: data <= 32'h3533b623;
    11'b00011011100: data <= 32'h390dbb44;
    11'b00011011101: data <= 32'hb924bcb9;
    11'b00011011110: data <= 32'hbf53bee6;
    11'b00011011111: data <= 32'hbc2bbf31;
    11'b00011100000: data <= 32'h3ac9b8f4;
    11'b00011100001: data <= 32'h3d6d3ad5;
    11'b00011100010: data <= 32'hadb23c26;
    11'b00011100011: data <= 32'hbe583292;
    11'b00011100100: data <= 32'hbeb730e8;
    11'b00011100101: data <= 32'hbc353d08;
    11'b00011100110: data <= 32'hba2a3eb0;
    11'b00011100111: data <= 32'hb78933a9;
    11'b00011101000: data <= 32'h3842bd89;
    11'b00011101001: data <= 32'h3e27bb7e;
    11'b00011101010: data <= 32'h3d9a3c7a;
    11'b00011101011: data <= 32'h3877406e;
    11'b00011101100: data <= 32'h37383d0f;
    11'b00011101101: data <= 32'h3c43b23e;
    11'b00011101110: data <= 32'h3aa0b930;
    11'b00011101111: data <= 32'hb93fb8db;
    11'b00011110000: data <= 32'hbdf0bc74;
    11'b00011110001: data <= 32'hb1f6bede;
    11'b00011110010: data <= 32'h3f1ebd70;
    11'b00011110011: data <= 32'h3f56b60f;
    11'b00011110100: data <= 32'haffd1a1a;
    11'b00011110101: data <= 32'hbedeb287;
    11'b00011110110: data <= 32'hbe2e311b;
    11'b00011110111: data <= 32'hba703c6d;
    11'b00011111000: data <= 32'hbb793c48;
    11'b00011111001: data <= 32'hbd7bb805;
    11'b00011111010: data <= 32'hbaa2bed0;
    11'b00011111011: data <= 32'h364eb924;
    11'b00011111100: data <= 32'h3bb03e9e;
    11'b00011111101: data <= 32'h399b4108;
    11'b00011111110: data <= 32'h38ef3d49;
    11'b00011111111: data <= 32'h3ad42d69;
    11'b00100000000: data <= 32'h367133d2;
    11'b00100000001: data <= 32'hba1f39ad;
    11'b00100000010: data <= 32'hbbdfa8b5;
    11'b00100000011: data <= 32'h3931bdab;
    11'b00100000100: data <= 32'h40d5bf13;
    11'b00100000101: data <= 32'h402dbb76;
    11'b00100000110: data <= 32'h2f75b2ae;
    11'b00100000111: data <= 32'hbc1faf65;
    11'b00100001000: data <= 32'hb7682d25;
    11'b00100001001: data <= 32'h2c3c380c;
    11'b00100001010: data <= 32'hbaef2f60;
    11'b00100001011: data <= 32'hc035bd29;
    11'b00100001100: data <= 32'hbf1fc007;
    11'b00100001101: data <= 32'hb226b9bb;
    11'b00100001110: data <= 32'h3a693d52;
    11'b00100001111: data <= 32'h38563f4f;
    11'b00100010000: data <= 32'h2b9639fe;
    11'b00100010001: data <= 32'ha7933404;
    11'b00100010010: data <= 32'hb54e3cfc;
    11'b00100010011: data <= 32'hbbd43fec;
    11'b00100010100: data <= 32'hba703a8a;
    11'b00100010101: data <= 32'h39febca2;
    11'b00100010110: data <= 32'h405ebecf;
    11'b00100010111: data <= 32'h3f60b8af;
    11'b00100011000: data <= 32'h37363715;
    11'b00100011001: data <= 32'h2dae369b;
    11'b00100011010: data <= 32'h3bac2d5a;
    11'b00100011011: data <= 32'h3c2928fa;
    11'b00100011100: data <= 32'hb93cb600;
    11'b00100011101: data <= 32'hc096bddb;
    11'b00100011110: data <= 32'hbf35c013;
    11'b00100011111: data <= 32'h2f54bc70;
    11'b00100100000: data <= 32'h3c42347d;
    11'b00100100001: data <= 32'h351b3799;
    11'b00100100010: data <= 32'hb944b164;
    11'b00100100011: data <= 32'hba783252;
    11'b00100100100: data <= 32'hba203f22;
    11'b00100100101: data <= 32'hbc8140ec;
    11'b00100100110: data <= 32'hbc793b48;
    11'b00100100111: data <= 32'hac21bcb7;
    11'b00100101000: data <= 32'h3c63bd62;
    11'b00100101001: data <= 32'h3c933419;
    11'b00100101010: data <= 32'h39003d74;
    11'b00100101011: data <= 32'h3bb93b81;
    11'b00100101100: data <= 32'h3f8031b3;
    11'b00100101101: data <= 32'h3e042fc8;
    11'b00100101110: data <= 32'hb8182d36;
    11'b00100101111: data <= 32'hbfd9ba00;
    11'b00100110000: data <= 32'hbc23be90;
    11'b00100110001: data <= 32'h3bfabe18;
    11'b00100110010: data <= 32'h3e21bace;
    11'b00100110011: data <= 32'h334eb9ef;
    11'b00100110100: data <= 32'hbb5cbb0b;
    11'b00100110101: data <= 32'hba351f64;
    11'b00100110110: data <= 32'hb7033e88;
    11'b00100110111: data <= 32'hbc043fe3;
    11'b00100111000: data <= 32'hbece3406;
    11'b00100111001: data <= 32'hbd44bdeb;
    11'b00100111010: data <= 32'hb365bc1b;
    11'b00100111011: data <= 32'h35f53b09;
    11'b00100111100: data <= 32'h383f3eff;
    11'b00100111101: data <= 32'h3c783b81;
    11'b00100111110: data <= 32'h3f3132d2;
    11'b00100111111: data <= 32'h3cce39c4;
    11'b00101000000: data <= 32'hb8ae3d24;
    11'b00101000001: data <= 32'hbdd2380d;
    11'b00101000010: data <= 32'hb0bdbbec;
    11'b00101000011: data <= 32'h3ecebea5;
    11'b00101000100: data <= 32'h3f03bd7f;
    11'b00101000101: data <= 32'h344dbc72;
    11'b00101000110: data <= 32'hb7efbbaf;
    11'b00101000111: data <= 32'h3241b057;
    11'b00101001000: data <= 32'h38cf3c28;
    11'b00101001001: data <= 32'hb8a73c00;
    11'b00101001010: data <= 32'hc047b8af;
    11'b00101001011: data <= 32'hc072bf1b;
    11'b00101001100: data <= 32'hbbfabb8b;
    11'b00101001101: data <= 32'h9ccf3a47;
    11'b00101001110: data <= 32'h34583cac;
    11'b00101001111: data <= 32'h389232d9;
    11'b00101010000: data <= 32'h3b772841;
    11'b00101010001: data <= 32'h37173dac;
    11'b00101010010: data <= 32'hba614101;
    11'b00101010011: data <= 32'hbca43e3b;
    11'b00101010100: data <= 32'h30bfb77a;
    11'b00101010101: data <= 32'h3e4fbdcf;
    11'b00101010110: data <= 32'h3d84bc25;
    11'b00101010111: data <= 32'h346eb81d;
    11'b00101011000: data <= 32'h351db711;
    11'b00101011001: data <= 32'h3e39b02f;
    11'b00101011010: data <= 32'h3f2337e5;
    11'b00101011011: data <= 32'hac48358e;
    11'b00101011100: data <= 32'hc04bbaef;
    11'b00101011101: data <= 32'hc07fbece;
    11'b00101011110: data <= 32'hba3abc29;
    11'b00101011111: data <= 32'h329d27c3;
    11'b00101100000: data <= 32'h292daf8b;
    11'b00101100001: data <= 32'hb24dbb5b;
    11'b00101100010: data <= 32'h26afb5a1;
    11'b00101100011: data <= 32'hae2e3ef5;
    11'b00101100100: data <= 32'hbb0641f6;
    11'b00101100101: data <= 32'hbcdb3f16;
    11'b00101100110: data <= 32'hb623b637;
    11'b00101100111: data <= 32'h3881bc43;
    11'b00101101000: data <= 32'h3774b13e;
    11'b00101101001: data <= 32'h2e7337ff;
    11'b00101101010: data <= 32'h3ba231bf;
    11'b00101101011: data <= 32'h40eeacae;
    11'b00101101100: data <= 32'h40cf35b8;
    11'b00101101101: data <= 32'h33433852;
    11'b00101101110: data <= 32'hbf05b394;
    11'b00101101111: data <= 32'hbdd8bc6a;
    11'b00101110000: data <= 32'h312fbc63;
    11'b00101110001: data <= 32'h3a04bab8;
    11'b00101110010: data <= 32'hac43bd4e;
    11'b00101110011: data <= 32'hb917bf48;
    11'b00101110100: data <= 32'hb1dcb9f4;
    11'b00101110101: data <= 32'h30523dfc;
    11'b00101110110: data <= 32'hb8a740f5;
    11'b00101110111: data <= 32'hbdcb3c5e;
    11'b00101111000: data <= 32'hbd73b9ed;
    11'b00101111001: data <= 32'hba07b9ec;
    11'b00101111010: data <= 32'hb82e38d2;
    11'b00101111011: data <= 32'hb3d23c6a;
    11'b00101111100: data <= 32'h3bd83494;
    11'b00101111101: data <= 32'h40c6b1ce;
    11'b00101111110: data <= 32'h403e3907;
    11'b00101111111: data <= 32'h30603ddf;
    11'b00110000000: data <= 32'hbcf93c01;
    11'b00110000001: data <= 32'hb75cb2fe;
    11'b00110000010: data <= 32'h3c3dbb88;
    11'b00110000011: data <= 32'h3c59bcd3;
    11'b00110000100: data <= 32'hb05bbed3;
    11'b00110000101: data <= 32'hb81abfdd;
    11'b00110000110: data <= 32'h381cbb52;
    11'b00110000111: data <= 32'h3c943b19;
    11'b00110001000: data <= 32'h2d293dab;
    11'b00110001001: data <= 32'hbe412d80;
    11'b00110001010: data <= 32'hc02bbc9e;
    11'b00110001011: data <= 32'hbe25b89e;
    11'b00110001100: data <= 32'hbc0d3a39;
    11'b00110001101: data <= 32'hb8ab3a54;
    11'b00110001110: data <= 32'h366db64c;
    11'b00110001111: data <= 32'h3dd2b8bf;
    11'b00110010000: data <= 32'h3ce53be5;
    11'b00110010001: data <= 32'hb20e40f3;
    11'b00110010010: data <= 32'hbb274026;
    11'b00110010011: data <= 32'h2cf03769;
    11'b00110010100: data <= 32'h3cccb8c6;
    11'b00110010101: data <= 32'h3a34ba7f;
    11'b00110010110: data <= 32'hb57cbc40;
    11'b00110010111: data <= 32'ha8fdbd63;
    11'b00110011000: data <= 32'h3e9bba7d;
    11'b00110011001: data <= 32'h40b534ea;
    11'b00110011010: data <= 32'h3a56386b;
    11'b00110011011: data <= 32'hbd87b73a;
    11'b00110011100: data <= 32'hc00cbca5;
    11'b00110011101: data <= 32'hbd2cb7bd;
    11'b00110011110: data <= 32'hb9fc35c0;
    11'b00110011111: data <= 32'hb9f4b432;
    11'b00110100000: data <= 32'hb63bbe36;
    11'b00110100001: data <= 32'h35d4bcd0;
    11'b00110100010: data <= 32'h37003c4c;
    11'b00110100011: data <= 32'hb5fa41b1;
    11'b00110100100: data <= 32'hba4d4091;
    11'b00110100101: data <= 32'hb02a3851;
    11'b00110100110: data <= 32'h36d6b3b4;
    11'b00110100111: data <= 32'hb1062d5d;
    11'b00110101000: data <= 32'hba182ee5;
    11'b00110101001: data <= 32'h3539b7ed;
    11'b00110101010: data <= 32'h40ddb911;
    11'b00110101011: data <= 32'h41fa2999;
    11'b00110101100: data <= 32'h3c8b36fe;
    11'b00110101101: data <= 32'hbbc9acc2;
    11'b00110101110: data <= 32'hbcd3b87c;
    11'b00110101111: data <= 32'hb322b4ab;
    11'b00110110000: data <= 32'h18c9b2e5;
    11'b00110110001: data <= 32'hb9cebd4d;
    11'b00110110010: data <= 32'hbb6bc0fa;
    11'b00110110011: data <= 32'hb045becb;
    11'b00110110100: data <= 32'h36813a1d;
    11'b00110110101: data <= 32'hae354099;
    11'b00110110110: data <= 32'hba3d3e01;
    11'b00110110111: data <= 32'hba5f2416;
    11'b00110111000: data <= 32'hb9d1a850;
    11'b00110111001: data <= 32'hbcc93b69;
    11'b00110111010: data <= 32'hbd093bd5;
    11'b00110111011: data <= 32'h3390afa3;
    11'b00110111100: data <= 32'h4098b98c;
    11'b00110111101: data <= 32'h41432dd1;
    11'b00110111110: data <= 32'h3b543c2c;
    11'b00110111111: data <= 32'hb87d3bdf;
    11'b00111000000: data <= 32'hb08d3623;
    11'b00111000001: data <= 32'h3b612b6d;
    11'b00111000010: data <= 32'h38deb6b5;
    11'b00111000011: data <= 32'hb9c3be8a;
    11'b00111000100: data <= 32'hbc02c12f;
    11'b00111000101: data <= 32'h33b6bf28;
    11'b00111000110: data <= 32'h3ce0334b;
    11'b00111000111: data <= 32'h38f83cbb;
    11'b00111001000: data <= 32'hb95e344b;
    11'b00111001001: data <= 32'hbd40b953;
    11'b00111001010: data <= 32'hbdb82837;
    11'b00111001011: data <= 32'hbeba3d19;
    11'b00111001100: data <= 32'hbe4d3be2;
    11'b00111001101: data <= 32'hb4e3b8a9;
    11'b00111001110: data <= 32'h3d40bc97;
    11'b00111001111: data <= 32'h3e2032b4;
    11'b00111010000: data <= 32'h35583f41;
    11'b00111010001: data <= 32'hb52c3fdc;
    11'b00111010010: data <= 32'h385d3c5e;
    11'b00111010011: data <= 32'h3d813709;
    11'b00111010100: data <= 32'h3842a4ca;
    11'b00111010101: data <= 32'hbb97bb88;
    11'b00111010110: data <= 32'hba2abf35;
    11'b00111010111: data <= 32'h3c78bdce;
    11'b00111011000: data <= 32'h40a4b38a;
    11'b00111011001: data <= 32'h3d8a31f5;
    11'b00111011010: data <= 32'hb659b8a2;
    11'b00111011011: data <= 32'hbccfbb6b;
    11'b00111011100: data <= 32'hbc8a2fde;
    11'b00111011101: data <= 32'hbd213c5f;
    11'b00111011110: data <= 32'hbe2732c0;
    11'b00111011111: data <= 32'hbbe2be7a;
    11'b00111100000: data <= 32'h2edbbf4e;
    11'b00111100001: data <= 32'h37163102;
    11'b00111100010: data <= 32'hafe9402d;
    11'b00111100011: data <= 32'hb3f4403e;
    11'b00111100100: data <= 32'h38843c4e;
    11'b00111100101: data <= 32'h3b2e392b;
    11'b00111100110: data <= 32'hb42a3a44;
    11'b00111100111: data <= 32'hbdc63544;
    11'b00111101000: data <= 32'hb8a8b94c;
    11'b00111101001: data <= 32'h3f11bbe9;
    11'b00111101010: data <= 32'h41cdb708;
    11'b00111101011: data <= 32'h3eb7b088;
    11'b00111101100: data <= 32'had3fb813;
    11'b00111101101: data <= 32'hb734b7d9;
    11'b00111101110: data <= 32'h26413636;
    11'b00111101111: data <= 32'hb44039c7;
    11'b00111110000: data <= 32'hbcf0b981;
    11'b00111110001: data <= 32'hbdc4c100;
    11'b00111110010: data <= 32'hb8b2c0a0;
    11'b00111110011: data <= 32'h2ddbaf63;
    11'b00111110100: data <= 32'ha9373e4f;
    11'b00111110101: data <= 32'hb1ce3d07;
    11'b00111110110: data <= 32'h2fac3509;
    11'b00111110111: data <= 32'hac2a38a9;
    11'b00111111000: data <= 32'hbcf83e20;
    11'b00111111001: data <= 32'hbfe13d86;
    11'b00111111010: data <= 32'hb9852977;
    11'b00111111011: data <= 32'h3e87ba97;
    11'b00111111100: data <= 32'h40f2b6da;
    11'b00111111101: data <= 32'h3d07337b;
    11'b00111111110: data <= 32'h2d833543;
    11'b00111111111: data <= 32'h38263631;
    11'b01000000000: data <= 32'h3d593a60;
    11'b01000000001: data <= 32'h396238b3;
    11'b01000000010: data <= 32'hbbd0bbbf;
    11'b01000000011: data <= 32'hbe19c118;
    11'b01000000100: data <= 32'hb71ac07d;
    11'b01000000101: data <= 32'h3940b71d;
    11'b01000000110: data <= 32'h38bc385f;
    11'b01000000111: data <= 32'h1d7db03a;
    11'b01000001000: data <= 32'hb485b994;
    11'b01000001001: data <= 32'hb9a73605;
    11'b01000001010: data <= 32'hbebb3f73;
    11'b01000001011: data <= 32'hc05a3e76;
    11'b01000001100: data <= 32'hbc47b0be;
    11'b01000001101: data <= 32'h39c4bcaa;
    11'b01000001110: data <= 32'h3ceab646;
    11'b01000001111: data <= 32'h35a83ad5;
    11'b01000010000: data <= 32'h29293cdf;
    11'b01000010001: data <= 32'h3cac3c40;
    11'b01000010010: data <= 32'h40083c7a;
    11'b01000010011: data <= 32'h3b263b05;
    11'b01000010100: data <= 32'hbc3fb54b;
    11'b01000010101: data <= 32'hbd79be83;
    11'b01000010110: data <= 32'h3419be6c;
    11'b01000010111: data <= 32'h3e8cb8fe;
    11'b01000011000: data <= 32'h3d4fb65f;
    11'b01000011001: data <= 32'h3443bccf;
    11'b01000011010: data <= 32'hb351bd1d;
    11'b01000011011: data <= 32'hb72e349f;
    11'b01000011100: data <= 32'hbcb63ef8;
    11'b01000011101: data <= 32'hbf7b3c24;
    11'b01000011110: data <= 32'hbde9bc23;
    11'b01000011111: data <= 32'hb6cabf41;
    11'b01000100000: data <= 32'had15b782;
    11'b01000100001: data <= 32'hb71d3c8a;
    11'b01000100010: data <= 32'hae253d8f;
    11'b01000100011: data <= 32'h3ced3bb6;
    11'b01000100100: data <= 32'h3efc3c67;
    11'b01000100101: data <= 32'h34833dbc;
    11'b01000100110: data <= 32'hbe0e3b03;
    11'b01000100111: data <= 32'hbcecb46e;
    11'b01000101000: data <= 32'h3aeeba4f;
    11'b01000101001: data <= 32'h406bb8b1;
    11'b01000101010: data <= 32'h3e3fba04;
    11'b01000101011: data <= 32'h3683bd6d;
    11'b01000101100: data <= 32'h3508bc3a;
    11'b01000101101: data <= 32'h393537e1;
    11'b01000101110: data <= 32'h28d23dc0;
    11'b01000101111: data <= 32'hbcd832cc;
    11'b01000110000: data <= 32'hbeadbf8c;
    11'b01000110001: data <= 32'hbc81c085;
    11'b01000110010: data <= 32'hb957b8f1;
    11'b01000110011: data <= 32'hb8eb3a51;
    11'b01000110100: data <= 32'hafa1389e;
    11'b01000110101: data <= 32'h3ae325d1;
    11'b01000110110: data <= 32'h3b25398e;
    11'b01000110111: data <= 32'hb9333fa1;
    11'b01000111000: data <= 32'hc0093faf;
    11'b01000111001: data <= 32'hbd0c3966;
    11'b01000111010: data <= 32'h3ad8b552;
    11'b01000111011: data <= 32'h3f4eb72f;
    11'b01000111100: data <= 32'h3bddb72f;
    11'b01000111101: data <= 32'h341db943;
    11'b01000111110: data <= 32'h3c0db41a;
    11'b01000111111: data <= 32'h3fc93b1e;
    11'b01001000000: data <= 32'h3cea3d15;
    11'b01001000001: data <= 32'hb908b0cb;
    11'b01001000010: data <= 32'hbe5abfe2;
    11'b01001000011: data <= 32'hbc30c020;
    11'b01001000100: data <= 32'hb459b94f;
    11'b01001000101: data <= 32'hadf923a0;
    11'b01001000110: data <= 32'h2b04ba53;
    11'b01001000111: data <= 32'h3767bcf8;
    11'b01001001000: data <= 32'h32b1307b;
    11'b01001001001: data <= 32'hbc7d4014;
    11'b01001001010: data <= 32'hc042406b;
    11'b01001001011: data <= 32'hbd9b396f;
    11'b01001001100: data <= 32'h31b6b82f;
    11'b01001001101: data <= 32'h38d8b62d;
    11'b01001001110: data <= 32'hb165307f;
    11'b01001001111: data <= 32'hb0ce3381;
    11'b01001010000: data <= 32'h3dc23712;
    11'b01001010001: data <= 32'h41563c99;
    11'b01001010010: data <= 32'h3ead3d79;
    11'b01001010011: data <= 32'hb825347b;
    11'b01001010100: data <= 32'hbd86bc52;
    11'b01001010101: data <= 32'hb650bcc2;
    11'b01001010110: data <= 32'h3965b7ad;
    11'b01001010111: data <= 32'h3931b986;
    11'b01001011000: data <= 32'h3481bf98;
    11'b01001011001: data <= 32'h35fcc022;
    11'b01001011010: data <= 32'h34a3b1f7;
    11'b01001011011: data <= 32'hb9363f5b;
    11'b01001011100: data <= 32'hbe723ebd;
    11'b01001011101: data <= 32'hbdd4b068;
    11'b01001011110: data <= 32'hb9c2bc9e;
    11'b01001011111: data <= 32'hb9e4b725;
    11'b01001100000: data <= 32'hbcee3824;
    11'b01001100001: data <= 32'hb88a3866;
    11'b01001100010: data <= 32'h3d8f3626;
    11'b01001100011: data <= 32'h40eb3b9f;
    11'b01001100100: data <= 32'h3ca53e63;
    11'b01001100101: data <= 32'hbb673cf7;
    11'b01001100110: data <= 32'hbcee34cb;
    11'b01001100111: data <= 32'h3463ade2;
    11'b01001101000: data <= 32'h3d70afe6;
    11'b01001101001: data <= 32'h3b6fbb34;
    11'b01001101010: data <= 32'h347fc03c;
    11'b01001101011: data <= 32'h3901bff3;
    11'b01001101100: data <= 32'h3c9cac34;
    11'b01001101101: data <= 32'h38ac3e14;
    11'b01001101110: data <= 32'hb9563aa8;
    11'b01001101111: data <= 32'hbd35bc47;
    11'b01001110000: data <= 32'hbd00be98;
    11'b01001110001: data <= 32'hbd93b7da;
    11'b01001110010: data <= 32'hbe5636c3;
    11'b01001110011: data <= 32'hb9bea917;
    11'b01001110100: data <= 32'h3befb888;
    11'b01001110101: data <= 32'h3e69344f;
    11'b01001110110: data <= 32'h31cf3ed7;
    11'b01001110111: data <= 32'hbde4402f;
    11'b01001111000: data <= 32'hbcc53d4b;
    11'b01001111001: data <= 32'h378b38b0;
    11'b01001111010: data <= 32'h3cb73219;
    11'b01001111011: data <= 32'h35a8b868;
    11'b01001111100: data <= 32'hb008bdbf;
    11'b01001111101: data <= 32'h3bb8bcb2;
    11'b01001111110: data <= 32'h407b35d3;
    11'b01001111111: data <= 32'h3f643d3a;
    11'b01010000000: data <= 32'h317c34cf;
    11'b01010000001: data <= 32'hbbf5bd5c;
    11'b01010000010: data <= 32'hbc66bde0;
    11'b01010000011: data <= 32'hbc24b4ea;
    11'b01010000100: data <= 32'hbc5e9f21;
    11'b01010000101: data <= 32'hb842bcc8;
    11'b01010000110: data <= 32'h3887bf9d;
    11'b01010000111: data <= 32'h3a48b889;
    11'b01010001000: data <= 32'hb75a3e4a;
    11'b01010001001: data <= 32'hbe784090;
    11'b01010001010: data <= 32'hbc8b3d87;
    11'b01010001011: data <= 32'h2f92378b;
    11'b01010001100: data <= 32'h3179346a;
    11'b01010001101: data <= 32'hbaed2b80;
    11'b01010001110: data <= 32'hbaa4b71f;
    11'b01010001111: data <= 32'h3c59b540;
    11'b01010010000: data <= 32'h41ae3965;
    11'b01010010001: data <= 32'h40b73cfc;
    11'b01010010010: data <= 32'h368236f0;
    11'b01010010011: data <= 32'hb9c4b949;
    11'b01010010100: data <= 32'hb6c5b84c;
    11'b01010010101: data <= 32'ha57531b1;
    11'b01010010110: data <= 32'hb34eb629;
    11'b01010010111: data <= 32'hb3dac054;
    11'b01010011000: data <= 32'h35b5c1a0;
    11'b01010011001: data <= 32'h38ccbc43;
    11'b01010011010: data <= 32'hb2603d06;
    11'b01010011011: data <= 32'hbc3d3ee3;
    11'b01010011100: data <= 32'hbb2f3835;
    11'b01010011101: data <= 32'hb70cb3eb;
    11'b01010011110: data <= 32'hbc133106;
    11'b01010011111: data <= 32'hc00e3831;
    11'b01010100000: data <= 32'hbddc2ea7;
    11'b01010100001: data <= 32'h3b00b1ab;
    11'b01010100010: data <= 32'h412a3763;
    11'b01010100011: data <= 32'h3f5b3cce;
    11'b01010100100: data <= 32'haa0d3c36;
    11'b01010100101: data <= 32'hb8ef3872;
    11'b01010100110: data <= 32'h34fb395b;
    11'b01010100111: data <= 32'h3aeb3a55;
    11'b01010101000: data <= 32'h3413b637;
    11'b01010101001: data <= 32'hb38ec0a3;
    11'b01010101010: data <= 32'h35dac180;
    11'b01010101011: data <= 32'h3c82bb8e;
    11'b01010101100: data <= 32'h3ae73ba8;
    11'b01010101101: data <= 32'h9d3a3a88;
    11'b01010101110: data <= 32'hb748b89f;
    11'b01010101111: data <= 32'hb9ccbb79;
    11'b01010110000: data <= 32'hbe662d21;
    11'b01010110001: data <= 32'hc0db3918;
    11'b01010110010: data <= 32'hbeaab152;
    11'b01010110011: data <= 32'h376bbb8d;
    11'b01010110100: data <= 32'h3eb6b52a;
    11'b01010110101: data <= 32'h39b93c0b;
    11'b01010110110: data <= 32'hba2c3e80;
    11'b01010110111: data <= 32'hb9013df8;
    11'b01010111000: data <= 32'h39773db4;
    11'b01010111001: data <= 32'h3be23cda;
    11'b01010111010: data <= 32'hb018238b;
    11'b01010111011: data <= 32'hb9cfbe60;
    11'b01010111100: data <= 32'h3666bf4c;
    11'b01010111101: data <= 32'h3faab5c4;
    11'b01010111110: data <= 32'h400d3a6a;
    11'b01010111111: data <= 32'h3b823076;
    11'b01011000000: data <= 32'h2430bc85;
    11'b01011000001: data <= 32'hb79cbba6;
    11'b01011000010: data <= 32'hbcc93529;
    11'b01011000011: data <= 32'hbf703802;
    11'b01011000100: data <= 32'hbd71bc0b;
    11'b01011000101: data <= 32'h2e0cc056;
    11'b01011000110: data <= 32'h39eabd21;
    11'b01011000111: data <= 32'hb2103948;
    11'b01011001000: data <= 32'hbc823eaf;
    11'b01011001001: data <= 32'hb84b3e03;
    11'b01011001010: data <= 32'h38d73d1a;
    11'b01011001011: data <= 32'h34ae3ce4;
    11'b01011001100: data <= 32'hbce638a4;
    11'b01011001101: data <= 32'hbe40b803;
    11'b01011001110: data <= 32'h3456b9e1;
    11'b01011001111: data <= 32'h40aa3156;
    11'b01011010000: data <= 32'h40f939e5;
    11'b01011010001: data <= 32'h3cb82504;
    11'b01011010010: data <= 32'h344bba22;
    11'b01011010011: data <= 32'h31cbb123;
    11'b01011010100: data <= 32'hae413b86;
    11'b01011010101: data <= 32'hba3b3664;
    11'b01011010110: data <= 32'hbaddbf0f;
    11'b01011010111: data <= 32'hadf7c20d;
    11'b01011011000: data <= 32'h3538bf4f;
    11'b01011011001: data <= 32'hb3d634eb;
    11'b01011011010: data <= 32'hb9cb3c64;
    11'b01011011011: data <= 32'hb1a43896;
    11'b01011011100: data <= 32'h356835f4;
    11'b01011011101: data <= 32'hb9453b39;
    11'b01011011110: data <= 32'hc0aa3c05;
    11'b01011011111: data <= 32'hc09033fc;
    11'b01011100000: data <= 32'ha861b455;
    11'b01011100001: data <= 32'h400d3032;
    11'b01011100010: data <= 32'h3f9a38b7;
    11'b01011100011: data <= 32'h38a0357c;
    11'b01011100100: data <= 32'h3258321e;
    11'b01011100101: data <= 32'h3af43be6;
    11'b01011100110: data <= 32'h3bbb3eae;
    11'b01011100111: data <= 32'h21353856;
    11'b01011101000: data <= 32'hb932bf58;
    11'b01011101001: data <= 32'hb116c1d0;
    11'b01011101010: data <= 32'h3880be67;
    11'b01011101011: data <= 32'h385230a1;
    11'b01011101100: data <= 32'h34303380;
    11'b01011101101: data <= 32'h367bb983;
    11'b01011101110: data <= 32'h33e0b8df;
    11'b01011101111: data <= 32'hbc7f38e1;
    11'b01011110000: data <= 32'hc1603ca7;
    11'b01011110001: data <= 32'hc0d93420;
    11'b01011110010: data <= 32'hb5adb9f7;
    11'b01011110011: data <= 32'h3c97b888;
    11'b01011110100: data <= 32'h39153401;
    11'b01011110101: data <= 32'hb6c8397c;
    11'b01011110110: data <= 32'ha8693bdb;
    11'b01011110111: data <= 32'h3d093ed8;
    11'b01011111000: data <= 32'h3d66402b;
    11'b01011111001: data <= 32'hac603b41;
    11'b01011111010: data <= 32'hbc1dbc7a;
    11'b01011111011: data <= 32'hb451bf6b;
    11'b01011111100: data <= 32'h3c61ba19;
    11'b01011111101: data <= 32'h3e2032c1;
    11'b01011111110: data <= 32'h3cbab713;
    11'b01011111111: data <= 32'h3b5bbdf5;
    11'b01100000000: data <= 32'h381abb90;
    11'b01100000001: data <= 32'hb9a939b8;
    11'b01100000010: data <= 32'hc0063ca1;
    11'b01100000011: data <= 32'hbf96b50d;
    11'b01100000100: data <= 32'hb81fbf18;
    11'b01100000101: data <= 32'h331abe04;
    11'b01100000110: data <= 32'hb809b1f8;
    11'b01100000111: data <= 32'hbc683943;
    11'b01100001000: data <= 32'haf113ba6;
    11'b01100001001: data <= 32'h3d2b3de9;
    11'b01100001010: data <= 32'h3b793faa;
    11'b01100001011: data <= 32'hbb8f3d27;
    11'b01100001100: data <= 32'hbf5aa9ab;
    11'b01100001101: data <= 32'hb820b85a;
    11'b01100001110: data <= 32'h3d8e2df0;
    11'b01100001111: data <= 32'h3fb63562;
    11'b01100010000: data <= 32'h3d74b933;
    11'b01100010001: data <= 32'h3c2ebda0;
    11'b01100010010: data <= 32'h3c18b646;
    11'b01100010011: data <= 32'h36013d2b;
    11'b01100010100: data <= 32'hb9d33cc5;
    11'b01100010101: data <= 32'hbc47bb40;
    11'b01100010110: data <= 32'hb7dec117;
    11'b01100010111: data <= 32'hb41dc006;
    11'b01100011000: data <= 32'hbabbb77f;
    11'b01100011001: data <= 32'hbbbb31e0;
    11'b01100011010: data <= 32'h32132858;
    11'b01100011011: data <= 32'h3cad3645;
    11'b01100011100: data <= 32'h31af3d24;
    11'b01100011101: data <= 32'hbfc83df8;
    11'b01100011110: data <= 32'hc1133a04;
    11'b01100011111: data <= 32'hba6e3271;
    11'b01100100000: data <= 32'h3c85359d;
    11'b01100100001: data <= 32'h3d5b346f;
    11'b01100100010: data <= 32'h38d5b78a;
    11'b01100100011: data <= 32'h398db959;
    11'b01100100100: data <= 32'h3df93906;
    11'b01100100101: data <= 32'h3de04009;
    11'b01100100110: data <= 32'h356d3d76;
    11'b01100100111: data <= 32'hb857bbd3;
    11'b01100101000: data <= 32'hb6fac0d1;
    11'b01100101001: data <= 32'hb0fbbe9f;
    11'b01100101010: data <= 32'hb4c7b637;
    11'b01100101011: data <= 32'hb042b7a5;
    11'b01100101100: data <= 32'h3a2fbcff;
    11'b01100101101: data <= 32'h3c99bae1;
    11'b01100101110: data <= 32'hb3d23942;
    11'b01100101111: data <= 32'hc08c3dfb;
    11'b01100110000: data <= 32'hc12a3b0b;
    11'b01100110001: data <= 32'hbb6ca290;
    11'b01100110010: data <= 32'h36dab13b;
    11'b01100110011: data <= 32'h2b19ab7d;
    11'b01100110100: data <= 32'hb944b36f;
    11'b01100110101: data <= 32'h2f8928cd;
    11'b01100110110: data <= 32'h3ed03d43;
    11'b01100110111: data <= 32'h3fd340bc;
    11'b01100111000: data <= 32'h384a3e58;
    11'b01100111001: data <= 32'hb9a2b677;
    11'b01100111010: data <= 32'hb836bd5b;
    11'b01100111011: data <= 32'h340ab894;
    11'b01100111100: data <= 32'h388f24a4;
    11'b01100111101: data <= 32'h39e7bbab;
    11'b01100111110: data <= 32'h3d05c047;
    11'b01100111111: data <= 32'h3d4fbdf0;
    11'b01101000000: data <= 32'h2c3e3813;
    11'b01101000001: data <= 32'hbe553dc6;
    11'b01101000010: data <= 32'hbf55370a;
    11'b01101000011: data <= 32'hba1abb13;
    11'b01101000100: data <= 32'hb4bcbc23;
    11'b01101000101: data <= 32'hbca8b7d2;
    11'b01101000110: data <= 32'hbe8ab333;
    11'b01101000111: data <= 32'hb3d12d06;
    11'b01101001000: data <= 32'h3ea23c47;
    11'b01101001001: data <= 32'h3eb24005;
    11'b01101001010: data <= 32'hb0f23eae;
    11'b01101001011: data <= 32'hbdb0378e;
    11'b01101001100: data <= 32'hba3d29a5;
    11'b01101001101: data <= 32'h384738b7;
    11'b01101001110: data <= 32'h3bf43758;
    11'b01101001111: data <= 32'h3b47bc3d;
    11'b01101010000: data <= 32'h3cefc060;
    11'b01101010001: data <= 32'h3e52bc94;
    11'b01101010010: data <= 32'h3bb43bbb;
    11'b01101010011: data <= 32'hb37a3df3;
    11'b01101010100: data <= 32'hb997ae8c;
    11'b01101010101: data <= 32'hb66bbe95;
    11'b01101010110: data <= 32'hb923be21;
    11'b01101010111: data <= 32'hbe86b950;
    11'b01101011000: data <= 32'hbef7b7d6;
    11'b01101011001: data <= 32'hae58b96b;
    11'b01101011010: data <= 32'h3e27ac9c;
    11'b01101011011: data <= 32'h3bf23c55;
    11'b01101011100: data <= 32'hbc723e18;
    11'b01101011101: data <= 32'hc0373c74;
    11'b01101011110: data <= 32'hbbfe3b56;
    11'b01101011111: data <= 32'h36ec3c7a;
    11'b01101100000: data <= 32'h385c38c2;
    11'b01101100001: data <= 32'h2ec2baf0;
    11'b01101100010: data <= 32'h38d8be2f;
    11'b01101100011: data <= 32'h3ecfb270;
    11'b01101100100: data <= 32'h3f8d3eae;
    11'b01101100101: data <= 32'h3ba93e7f;
    11'b01101100110: data <= 32'h3015b485;
    11'b01101100111: data <= 32'haeddbe7c;
    11'b01101101000: data <= 32'hb809bc90;
    11'b01101101001: data <= 32'hbccdb56e;
    11'b01101101010: data <= 32'hbc14ba96;
    11'b01101101011: data <= 32'h372fbf26;
    11'b01101101100: data <= 32'h3e06bdc5;
    11'b01101101101: data <= 32'h380e304e;
    11'b01101101110: data <= 32'hbe1a3cfe;
    11'b01101101111: data <= 32'hc0443cb7;
    11'b01101110000: data <= 32'hbb553aa1;
    11'b01101110001: data <= 32'h278f3a0b;
    11'b01101110010: data <= 32'hb88d351a;
    11'b01101110011: data <= 32'hbd14b90e;
    11'b01101110100: data <= 32'hb4cfba87;
    11'b01101110101: data <= 32'h3e683860;
    11'b01101110110: data <= 32'h40924007;
    11'b01101110111: data <= 32'h3d293eb8;
    11'b01101111000: data <= 32'h310f2787;
    11'b01101111001: data <= 32'hae8db9b2;
    11'b01101111010: data <= 32'hae9e29e7;
    11'b01101111011: data <= 32'hb57e365c;
    11'b01101111100: data <= 32'haf65bbca;
    11'b01101111101: data <= 32'h3b7dc122;
    11'b01101111110: data <= 32'h3e3fc06c;
    11'b01101111111: data <= 32'h38c3b3e2;
    11'b01110000000: data <= 32'hbbe03c3b;
    11'b01110000001: data <= 32'hbd2b39e8;
    11'b01110000010: data <= 32'hb6e893e3;
    11'b01110000011: data <= 32'hb5b7af69;
    11'b01110000100: data <= 32'hbeabafae;
    11'b01110000101: data <= 32'hc0cbb859;
    11'b01110000110: data <= 32'hbb78b8c2;
    11'b01110000111: data <= 32'h3d80370a;
    11'b01110001000: data <= 32'h3ff43e57;
    11'b01110001001: data <= 32'h39553ddd;
    11'b01110001010: data <= 32'hb8303893;
    11'b01110001011: data <= 32'hb5b63856;
    11'b01110001100: data <= 32'h33433d76;
    11'b01110001101: data <= 32'h33013c92;
    11'b01110001110: data <= 32'h31dabad0;
    11'b01110001111: data <= 32'h3aefc12b;
    11'b01110010000: data <= 32'h3e34bfd8;
    11'b01110010001: data <= 32'h3cb03042;
    11'b01110010010: data <= 32'h33673c56;
    11'b01110010011: data <= 32'h1a43316b;
    11'b01110010100: data <= 32'h3429bae2;
    11'b01110010101: data <= 32'hb716b9cc;
    11'b01110010110: data <= 32'hc02cb45e;
    11'b01110010111: data <= 32'hc13cb8b1;
    11'b01110011000: data <= 32'hbb4abc37;
    11'b01110011001: data <= 32'h3cd5b883;
    11'b01110011010: data <= 32'h3d2a3807;
    11'b01110011011: data <= 32'hb5a93bcc;
    11'b01110011100: data <= 32'hbd343b63;
    11'b01110011101: data <= 32'hb8973d6c;
    11'b01110011110: data <= 32'h34db4012;
    11'b01110011111: data <= 32'h28a93dcc;
    11'b01110100000: data <= 32'hb7b5b89e;
    11'b01110100001: data <= 32'h2e7dbfb9;
    11'b01110100010: data <= 32'h3d50bbe4;
    11'b01110100011: data <= 32'h3f263b3e;
    11'b01110100100: data <= 32'h3d683cec;
    11'b01110100101: data <= 32'h3bf0b0ca;
    11'b01110100110: data <= 32'h3a35bc48;
    11'b01110100111: data <= 32'hb1e1b794;
    11'b01110101000: data <= 32'hbe943153;
    11'b01110101001: data <= 32'hbf97b8b7;
    11'b01110101010: data <= 32'hb532bf63;
    11'b01110101011: data <= 32'h3cc2bf6a;
    11'b01110101100: data <= 32'h3999b900;
    11'b01110101101: data <= 32'hbbc636e3;
    11'b01110101110: data <= 32'hbddb3a99;
    11'b01110101111: data <= 32'hb6733d02;
    11'b01110110000: data <= 32'h328a3ed5;
    11'b01110110001: data <= 32'hba1e3cb2;
    11'b01110110010: data <= 32'hbf12b594;
    11'b01110110011: data <= 32'hbbf4bc7c;
    11'b01110110100: data <= 32'h3b60ac10;
    11'b01110110101: data <= 32'h3fec3d8c;
    11'b01110110110: data <= 32'h3ea73ce8;
    11'b01110110111: data <= 32'h3c64af0d;
    11'b01110111000: data <= 32'h3aa4b76c;
    11'b01110111001: data <= 32'h334c38f0;
    11'b01110111010: data <= 32'hb9d73c5f;
    11'b01110111011: data <= 32'hbaccb690;
    11'b01110111100: data <= 32'h34c0c0c8;
    11'b01110111101: data <= 32'h3cdbc131;
    11'b01110111110: data <= 32'h3867bc79;
    11'b01110111111: data <= 32'hb9c1305e;
    11'b01111000000: data <= 32'hb9d53583;
    11'b01111000001: data <= 32'h34333616;
    11'b01111000010: data <= 32'h311439d1;
    11'b01111000011: data <= 32'hbe6a38e7;
    11'b01111000100: data <= 32'hc1bbb409;
    11'b01111000101: data <= 32'hbf18b996;
    11'b01111000110: data <= 32'h384a2e9e;
    11'b01111000111: data <= 32'h3e6f3c4d;
    11'b01111001000: data <= 32'h3c083acd;
    11'b01111001001: data <= 32'h35842ddf;
    11'b01111001010: data <= 32'h37a23822;
    11'b01111001011: data <= 32'h386b3f9e;
    11'b01111001100: data <= 32'h0e784007;
    11'b01111001101: data <= 32'hb4b6acf5;
    11'b01111001110: data <= 32'h35c4c097;
    11'b01111001111: data <= 32'h3c45c0a4;
    11'b01111010000: data <= 32'h3a61b9aa;
    11'b01111010001: data <= 32'h32db333a;
    11'b01111010010: data <= 32'h383bb2ee;
    11'b01111010011: data <= 32'h3c9db8f0;
    11'b01111010100: data <= 32'h353faf85;
    11'b01111010101: data <= 32'hbf843508;
    11'b01111010110: data <= 32'hc223b228;
    11'b01111010111: data <= 32'hbf0ebac9;
    11'b01111011000: data <= 32'h3635b8e8;
    11'b01111011001: data <= 32'h3b472941;
    11'b01111011010: data <= 32'hb00e30b4;
    11'b01111011011: data <= 32'hb92930df;
    11'b01111011100: data <= 32'h2eef3ca1;
    11'b01111011101: data <= 32'h39974122;
    11'b01111011110: data <= 32'h2e7240c3;
    11'b01111011111: data <= 32'hb95d334b;
    11'b01111100000: data <= 32'hb578be7c;
    11'b01111100001: data <= 32'h3911bd01;
    11'b01111100010: data <= 32'h3c6233ed;
    11'b01111100011: data <= 32'h3c8b382b;
    11'b01111100100: data <= 32'h3e14b8a3;
    11'b01111100101: data <= 32'h3f1bbc54;
    11'b01111100110: data <= 32'h3961b0e5;
    11'b01111100111: data <= 32'hbd93395c;
    11'b01111101000: data <= 32'hc08b16b7;
    11'b01111101001: data <= 32'hbc1bbd40;
    11'b01111101010: data <= 32'h380cbebc;
    11'b01111101011: data <= 32'h34abbc60;
    11'b01111101100: data <= 32'hbbc9b864;
    11'b01111101101: data <= 32'hbc5cad94;
    11'b01111101110: data <= 32'h318d3be5;
    11'b01111101111: data <= 32'h3a31405e;
    11'b01111110000: data <= 32'hb5f63ffb;
    11'b01111110001: data <= 32'hbee2357d;
    11'b01111110010: data <= 32'hbdc5ba5f;
    11'b01111110011: data <= 32'h2936afd5;
    11'b01111110100: data <= 32'h3c643c05;
    11'b01111110101: data <= 32'h3d6c3925;
    11'b01111110110: data <= 32'h3e5fb97f;
    11'b01111110111: data <= 32'h3f16ba5c;
    11'b01111111000: data <= 32'h3c063984;
    11'b01111111001: data <= 32'hb7723e60;
    11'b01111111010: data <= 32'hbc293639;
    11'b01111111011: data <= 32'hb06dbe7c;
    11'b01111111100: data <= 32'h3964c09e;
    11'b01111111101: data <= 32'h25f0be4e;
    11'b01111111110: data <= 32'hbc1ebab6;
    11'b01111111111: data <= 32'hb8ebb846;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    