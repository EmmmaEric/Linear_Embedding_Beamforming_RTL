
module memory_rom_16(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h37133e19;
    11'b00000000001: data <= 32'h345d3a68;
    11'b00000000010: data <= 32'hb2f4bbb3;
    11'b00000000011: data <= 32'h3689bf52;
    11'b00000000100: data <= 32'h3e97b855;
    11'b00000000101: data <= 32'h3fd83d4c;
    11'b00000000110: data <= 32'h3cc13d66;
    11'b00000000111: data <= 32'h3772b52c;
    11'b00000001000: data <= 32'h2fdbbd67;
    11'b00000001001: data <= 32'hb8b1b9d0;
    11'b00000001010: data <= 32'hbe40ab7b;
    11'b00000001011: data <= 32'hbdbeba63;
    11'b00000001100: data <= 32'h30edbfbc;
    11'b00000001101: data <= 32'h3d74be9a;
    11'b00000001110: data <= 32'h3838ae2f;
    11'b00000001111: data <= 32'hbd253c45;
    11'b00000010000: data <= 32'hbede3cd9;
    11'b00000010001: data <= 32'hb86b3c9f;
    11'b00000010010: data <= 32'h2f0e3cdd;
    11'b00000010011: data <= 32'hba2a3918;
    11'b00000010100: data <= 32'hbe34b8b1;
    11'b00000010101: data <= 32'hb7f8bbcf;
    11'b00000010110: data <= 32'h3e123458;
    11'b00000010111: data <= 32'h40a93ea0;
    11'b00000011000: data <= 32'h3e1e3d53;
    11'b00000011001: data <= 32'h3877af45;
    11'b00000011010: data <= 32'h3387b848;
    11'b00000011011: data <= 32'hac143676;
    11'b00000011100: data <= 32'hb8e33954;
    11'b00000011101: data <= 32'hb801bb6d;
    11'b00000011110: data <= 32'h38c2c161;
    11'b00000011111: data <= 32'h3d3fc0d8;
    11'b00000100000: data <= 32'h37cbb83d;
    11'b00000100001: data <= 32'hbad33a4b;
    11'b00000100010: data <= 32'hbb7d3968;
    11'b00000100011: data <= 32'hacd53443;
    11'b00000100100: data <= 32'hb3f7359c;
    11'b00000100101: data <= 32'hbf55346a;
    11'b00000100110: data <= 32'hc155b5e2;
    11'b00000100111: data <= 32'hbca5b8e7;
    11'b00000101000: data <= 32'h3ce73460;
    11'b00000101001: data <= 32'h3fde3d1b;
    11'b00000101010: data <= 32'h3b063c6c;
    11'b00000101011: data <= 32'had903611;
    11'b00000101100: data <= 32'h2d32394e;
    11'b00000101101: data <= 32'h367f3ec3;
    11'b00000101110: data <= 32'h2db23dab;
    11'b00000101111: data <= 32'haeecba23;
    11'b00000110000: data <= 32'h3867c153;
    11'b00000110001: data <= 32'h3d09c055;
    11'b00000110010: data <= 32'h3bdcb27d;
    11'b00000110011: data <= 32'h347c39a2;
    11'b00000110100: data <= 32'h34e2a723;
    11'b00000110101: data <= 32'h38d4b9b0;
    11'b00000110110: data <= 32'hb506b528;
    11'b00000110111: data <= 32'hc0733036;
    11'b00000111000: data <= 32'hc1c6b55d;
    11'b00000111001: data <= 32'hbcc2bbb0;
    11'b00000111010: data <= 32'h3babb8fe;
    11'b00000111011: data <= 32'h3c9d3432;
    11'b00000111100: data <= 32'hb3693910;
    11'b00000111101: data <= 32'hbb2339b3;
    11'b00000111110: data <= 32'hadb53dcc;
    11'b00000111111: data <= 32'h38b540b5;
    11'b00001000000: data <= 32'h29093f0b;
    11'b00001000001: data <= 32'hb93cb6a5;
    11'b00001000010: data <= 32'hb0a2bfae;
    11'b00001000011: data <= 32'h3c30bc88;
    11'b00001000100: data <= 32'h3e43387e;
    11'b00001000101: data <= 32'h3d6e3a2c;
    11'b00001000110: data <= 32'h3d16b79c;
    11'b00001000111: data <= 32'h3c8abc3f;
    11'b00001001000: data <= 32'h9c43b1e8;
    11'b00001001001: data <= 32'hbee4381e;
    11'b00001001010: data <= 32'hc046b545;
    11'b00001001011: data <= 32'hb915bec9;
    11'b00001001100: data <= 32'h3abcbf61;
    11'b00001001101: data <= 32'h36c8ba8f;
    11'b00001001110: data <= 32'hbbdf2e08;
    11'b00001001111: data <= 32'hbc9638af;
    11'b00001010000: data <= 32'h2af93d3c;
    11'b00001010001: data <= 32'h383c4008;
    11'b00001010010: data <= 32'hb9663e1d;
    11'b00001010011: data <= 32'hbf5fad98;
    11'b00001010100: data <= 32'hbcafbbda;
    11'b00001010101: data <= 32'h394dae0d;
    11'b00001010110: data <= 32'h3ef73c6b;
    11'b00001010111: data <= 32'h3e913a0d;
    11'b00001011000: data <= 32'h3d7eb819;
    11'b00001011001: data <= 32'h3cebb88f;
    11'b00001011010: data <= 32'h37e63a52;
    11'b00001011011: data <= 32'hb99d3d70;
    11'b00001011100: data <= 32'hbc02b1ad;
    11'b00001011101: data <= 32'h22b9c071;
    11'b00001011110: data <= 32'h3a8cc11a;
    11'b00001011111: data <= 32'h314cbd31;
    11'b00001100000: data <= 32'hbaf0b33a;
    11'b00001100001: data <= 32'hb8462934;
    11'b00001100010: data <= 32'h392335c3;
    11'b00001100011: data <= 32'h37753bdc;
    11'b00001100100: data <= 32'hbdea3bc6;
    11'b00001100101: data <= 32'hc1c52d62;
    11'b00001100110: data <= 32'hbfa6b6dd;
    11'b00001100111: data <= 32'h345d32e7;
    11'b00001101000: data <= 32'h3d503b45;
    11'b00001101001: data <= 32'h3b7c36fe;
    11'b00001101010: data <= 32'h38c1b518;
    11'b00001101011: data <= 32'h3b3e359d;
    11'b00001101100: data <= 32'h3b413ffc;
    11'b00001101101: data <= 32'h311d406e;
    11'b00001101110: data <= 32'hb5003053;
    11'b00001101111: data <= 32'h3178c035;
    11'b00001110000: data <= 32'h3994c07b;
    11'b00001110001: data <= 32'h35e5bb04;
    11'b00001110010: data <= 32'ha68cb197;
    11'b00001110011: data <= 32'h38f2b8e0;
    11'b00001110100: data <= 32'h3dcdba0b;
    11'b00001110101: data <= 32'h38cc2713;
    11'b00001110110: data <= 32'hbef938e1;
    11'b00001110111: data <= 32'hc21d30eb;
    11'b00001111000: data <= 32'hbf8fb7fa;
    11'b00001111001: data <= 32'h2df6b611;
    11'b00001111010: data <= 32'h386d9988;
    11'b00001111011: data <= 32'hb4b7b1a9;
    11'b00001111100: data <= 32'hb791b320;
    11'b00001111101: data <= 32'h38153bce;
    11'b00001111110: data <= 32'h3c63413c;
    11'b00001111111: data <= 32'h35e2411b;
    11'b00010000000: data <= 32'hb862373c;
    11'b00010000001: data <= 32'hb66cbd81;
    11'b00010000010: data <= 32'h3588bc68;
    11'b00010000011: data <= 32'h397c3005;
    11'b00010000100: data <= 32'h3ae22f51;
    11'b00010000101: data <= 32'h3e30bc2b;
    11'b00010000110: data <= 32'h400bbd5e;
    11'b00010000111: data <= 32'h3b72b0cf;
    11'b00010001000: data <= 32'hbceb3ac3;
    11'b00010001001: data <= 32'hc06d3495;
    11'b00010001010: data <= 32'hbc82bb9f;
    11'b00010001011: data <= 32'h31ecbd87;
    11'b00010001100: data <= 32'hb0bcbc31;
    11'b00010001101: data <= 32'hbd0eba63;
    11'b00010001110: data <= 32'hbc2eb6da;
    11'b00010001111: data <= 32'h37b23a5d;
    11'b00010010000: data <= 32'h3c914068;
    11'b00010010001: data <= 32'habc5404e;
    11'b00010010010: data <= 32'hbdfd38c4;
    11'b00010010011: data <= 32'hbd8ab787;
    11'b00010010100: data <= 32'hb0f83060;
    11'b00010010101: data <= 32'h39d63be2;
    11'b00010010110: data <= 32'h3c4c34b6;
    11'b00010010111: data <= 32'h3e5cbca1;
    11'b00010011000: data <= 32'h3ffbbc88;
    11'b00010011001: data <= 32'h3d1f3886;
    11'b00010011010: data <= 32'hb3a53e8a;
    11'b00010011011: data <= 32'hbb2a3899;
    11'b00010011100: data <= 32'hb14fbd33;
    11'b00010011101: data <= 32'h3604bff5;
    11'b00010011110: data <= 32'hb75dbdf1;
    11'b00010011111: data <= 32'hbdb2bc34;
    11'b00010100000: data <= 32'hb9adbafa;
    11'b00010100001: data <= 32'h3bf6b039;
    11'b00010100010: data <= 32'h3ce53c04;
    11'b00010100011: data <= 32'hb93c3d2f;
    11'b00010100100: data <= 32'hc0d43854;
    11'b00010100101: data <= 32'hc0332f3e;
    11'b00010100110: data <= 32'hb83f39bf;
    11'b00010100111: data <= 32'h35d23c58;
    11'b00010101000: data <= 32'h35fe2cb5;
    11'b00010101001: data <= 32'h3959bc6d;
    11'b00010101010: data <= 32'h3d96b727;
    11'b00010101011: data <= 32'h3ddf3e7e;
    11'b00010101100: data <= 32'h391540f4;
    11'b00010101101: data <= 32'h2b713b60;
    11'b00010101110: data <= 32'h34edbcb4;
    11'b00010101111: data <= 32'h3621beaa;
    11'b00010110000: data <= 32'hb63bbb91;
    11'b00010110001: data <= 32'hbaaeba1b;
    11'b00010110010: data <= 32'h3457bd3d;
    11'b00010110011: data <= 32'h3f2cbcfe;
    11'b00010110100: data <= 32'h3dbbb28e;
    11'b00010110101: data <= 32'hbae638d3;
    11'b00010110110: data <= 32'hc11b3736;
    11'b00010110111: data <= 32'hbff03114;
    11'b00010111000: data <= 32'hb829363e;
    11'b00010111001: data <= 32'hb34835f5;
    11'b00010111010: data <= 32'hbad2b837;
    11'b00010111011: data <= 32'hb91dbc79;
    11'b00010111100: data <= 32'h394d2cff;
    11'b00010111101: data <= 32'h3de04063;
    11'b00010111110: data <= 32'h3b80417f;
    11'b00010111111: data <= 32'h2e673c66;
    11'b00011000000: data <= 32'ha8b2b8c4;
    11'b00011000001: data <= 32'h2b91b838;
    11'b00011000010: data <= 32'hb275347e;
    11'b00011000011: data <= 32'had94b076;
    11'b00011000100: data <= 32'h3c8bbe24;
    11'b00011000101: data <= 32'h40a8bfa3;
    11'b00011000110: data <= 32'h3eb7b955;
    11'b00011000111: data <= 32'hb74638a1;
    11'b00011001000: data <= 32'hbed2383e;
    11'b00011001001: data <= 32'hbc12b0fd;
    11'b00011001010: data <= 32'haeebb70c;
    11'b00011001011: data <= 32'hb9b6b8b9;
    11'b00011001100: data <= 32'hbf85bc8c;
    11'b00011001101: data <= 32'hbdffbd2c;
    11'b00011001110: data <= 32'h357fa908;
    11'b00011001111: data <= 32'h3db83f17;
    11'b00011010000: data <= 32'h392d4057;
    11'b00011010001: data <= 32'hb92f3b99;
    11'b00011010010: data <= 32'hbb502e4e;
    11'b00011010011: data <= 32'hb7213a15;
    11'b00011010100: data <= 32'hb1a93db9;
    11'b00011010101: data <= 32'h30ac35b7;
    11'b00011010110: data <= 32'h3cacbe23;
    11'b00011010111: data <= 32'h4051bf52;
    11'b00011011000: data <= 32'h3f16b1a0;
    11'b00011011001: data <= 32'h35693cee;
    11'b00011011010: data <= 32'hb5823a9c;
    11'b00011011011: data <= 32'h3371b718;
    11'b00011011100: data <= 32'h36b7bc18;
    11'b00011011101: data <= 32'hbb0dbc0d;
    11'b00011011110: data <= 32'hc052bd24;
    11'b00011011111: data <= 32'hbda4be1d;
    11'b00011100000: data <= 32'h3985ba54;
    11'b00011100001: data <= 32'h3e0a384c;
    11'b00011100010: data <= 32'h30893c21;
    11'b00011100011: data <= 32'hbe02385e;
    11'b00011100100: data <= 32'hbe6d381c;
    11'b00011100101: data <= 32'hba0a3dd2;
    11'b00011100110: data <= 32'hb6383f34;
    11'b00011100111: data <= 32'hb687356e;
    11'b00011101000: data <= 32'h32f2bddc;
    11'b00011101001: data <= 32'h3d2fbd00;
    11'b00011101010: data <= 32'h3e713a47;
    11'b00011101011: data <= 32'h3c1c4015;
    11'b00011101100: data <= 32'h39b93c8e;
    11'b00011101101: data <= 32'h3bfbb6ba;
    11'b00011101110: data <= 32'h395aba81;
    11'b00011101111: data <= 32'hba28b735;
    11'b00011110000: data <= 32'hbec4ba1b;
    11'b00011110001: data <= 32'hb877be8a;
    11'b00011110010: data <= 32'h3dc1bedc;
    11'b00011110011: data <= 32'h3ed6ba29;
    11'b00011110100: data <= 32'haf892787;
    11'b00011110101: data <= 32'hbee03192;
    11'b00011110110: data <= 32'hbde637da;
    11'b00011110111: data <= 32'hb85e3d04;
    11'b00011111000: data <= 32'hb96d3cff;
    11'b00011111001: data <= 32'hbdc9b213;
    11'b00011111010: data <= 32'hbcb9bded;
    11'b00011111011: data <= 32'h33c3b9ba;
    11'b00011111100: data <= 32'h3d303d9c;
    11'b00011111101: data <= 32'h3ced409c;
    11'b00011111110: data <= 32'h3b1e3ca2;
    11'b00011111111: data <= 32'h3ad0ae8a;
    11'b00100000000: data <= 32'h372930ca;
    11'b00100000001: data <= 32'hb8ba3ade;
    11'b00100000010: data <= 32'hbbc131c5;
    11'b00100000011: data <= 32'h3527be17;
    11'b00100000100: data <= 32'h3fe3c081;
    11'b00100000101: data <= 32'h3f5abd77;
    11'b00100000110: data <= 32'h2c8fb35f;
    11'b00100000111: data <= 32'hbc1f2f1d;
    11'b00100001000: data <= 32'hb6f931b8;
    11'b00100001001: data <= 32'h319737aa;
    11'b00100001010: data <= 32'hba8c34d5;
    11'b00100001011: data <= 32'hc0aaba67;
    11'b00100001100: data <= 32'hc05bbe51;
    11'b00100001101: data <= 32'hb58bb948;
    11'b00100001110: data <= 32'h3c483c7d;
    11'b00100001111: data <= 32'h3b6b3eaa;
    11'b00100010000: data <= 32'h331739c3;
    11'b00100010001: data <= 32'h26913403;
    11'b00100010010: data <= 32'haab23d25;
    11'b00100010011: data <= 32'hb831404b;
    11'b00100010100: data <= 32'hb8de3bd0;
    11'b00100010101: data <= 32'h37a2bd29;
    11'b00100010110: data <= 32'h3f0bc046;
    11'b00100010111: data <= 32'h3eb2bbcd;
    11'b00100011000: data <= 32'h384d3553;
    11'b00100011001: data <= 32'h31a03627;
    11'b00100011010: data <= 32'h3ba0b00b;
    11'b00100011011: data <= 32'h3c1ab207;
    11'b00100011100: data <= 32'hb9bcb325;
    11'b00100011101: data <= 32'hc11cbb6f;
    11'b00100011110: data <= 32'hc069be63;
    11'b00100011111: data <= 32'hb040bc70;
    11'b00100100000: data <= 32'h3c66293e;
    11'b00100100001: data <= 32'h36ab3650;
    11'b00100100010: data <= 32'hb96da55c;
    11'b00100100011: data <= 32'hb9f935de;
    11'b00100100100: data <= 32'hb5c33f9e;
    11'b00100100101: data <= 32'hb880414c;
    11'b00100100110: data <= 32'hbb263c8a;
    11'b00100100111: data <= 32'hb523bc89;
    11'b00100101000: data <= 32'h3a36be37;
    11'b00100101001: data <= 32'h3cb095bf;
    11'b00100101010: data <= 32'h3b413cc7;
    11'b00100101011: data <= 32'h3c9439a8;
    11'b00100101100: data <= 32'h3f79b374;
    11'b00100101101: data <= 32'h3dfdb2b1;
    11'b00100101110: data <= 32'hb7a73219;
    11'b00100101111: data <= 32'hc027b4de;
    11'b00100110000: data <= 32'hbd7abd80;
    11'b00100110001: data <= 32'h391dbed1;
    11'b00100110010: data <= 32'h3d3fbca8;
    11'b00100110011: data <= 32'h2c1aba31;
    11'b00100110100: data <= 32'hbc5ab947;
    11'b00100110101: data <= 32'hba0f318e;
    11'b00100110110: data <= 32'hacae3ec0;
    11'b00100110111: data <= 32'hb8664049;
    11'b00100111000: data <= 32'hbe6b38f3;
    11'b00100111001: data <= 32'hbe6ebca0;
    11'b00100111010: data <= 32'hb736bba2;
    11'b00100111011: data <= 32'h386e3a32;
    11'b00100111100: data <= 32'h3b2f3e5e;
    11'b00100111101: data <= 32'h3d2c3966;
    11'b00100111110: data <= 32'h3f34b1d7;
    11'b00100111111: data <= 32'h3d54370d;
    11'b00101000000: data <= 32'hb49f3d87;
    11'b00101000001: data <= 32'hbd3e3a81;
    11'b00101000010: data <= 32'hb5cdbb74;
    11'b00101000011: data <= 32'h3d30bff7;
    11'b00101000100: data <= 32'h3da7bee5;
    11'b00101000101: data <= 32'h25e0bc94;
    11'b00101000110: data <= 32'hb98bbaa5;
    11'b00101000111: data <= 32'h3119b1a6;
    11'b00101001000: data <= 32'h3a823b10;
    11'b00101001001: data <= 32'hb58e3c6a;
    11'b00101001010: data <= 32'hc06daea7;
    11'b00101001011: data <= 32'hc11dbd00;
    11'b00101001100: data <= 32'hbcb9b9a6;
    11'b00101001101: data <= 32'h31453a1f;
    11'b00101001110: data <= 32'h38273c54;
    11'b00101001111: data <= 32'h38d42d85;
    11'b00101010000: data <= 32'h3b58b17d;
    11'b00101010001: data <= 32'h39ef3d23;
    11'b00101010010: data <= 32'hb373413b;
    11'b00101010011: data <= 32'hba5a3f1a;
    11'b00101010100: data <= 32'h2942b7c3;
    11'b00101010101: data <= 32'h3ce4bf0a;
    11'b00101010110: data <= 32'h3c7dbd40;
    11'b00101010111: data <= 32'h311bb880;
    11'b00101011000: data <= 32'h32dfb800;
    11'b00101011001: data <= 32'h3df4b776;
    11'b00101011010: data <= 32'h3f672ded;
    11'b00101011011: data <= 32'h234c35a9;
    11'b00101011100: data <= 32'hc090b60b;
    11'b00101011101: data <= 32'hc121bcaf;
    11'b00101011110: data <= 32'hbbe9bac7;
    11'b00101011111: data <= 32'h32a4a422;
    11'b00101100000: data <= 32'h238fafdb;
    11'b00101100001: data <= 32'hb646bad5;
    11'b00101100010: data <= 32'haaa5b5a0;
    11'b00101100011: data <= 32'h348a3edc;
    11'b00101100100: data <= 32'hb2a74233;
    11'b00101100101: data <= 32'hba653ffd;
    11'b00101100110: data <= 32'hb75cb4af;
    11'b00101100111: data <= 32'h3513bca7;
    11'b00101101000: data <= 32'h36b6b435;
    11'b00101101001: data <= 32'h329e3773;
    11'b00101101010: data <= 32'h3bbfa7e8;
    11'b00101101011: data <= 32'h40c7b8db;
    11'b00101101100: data <= 32'h40dab199;
    11'b00101101101: data <= 32'h357d37a3;
    11'b00101101110: data <= 32'hbf0d30db;
    11'b00101101111: data <= 32'hbeacba11;
    11'b00101110000: data <= 32'had4abc6c;
    11'b00101110001: data <= 32'h386abbde;
    11'b00101110010: data <= 32'hb5a0bd1e;
    11'b00101110011: data <= 32'hbc11be8d;
    11'b00101110100: data <= 32'hb57ab984;
    11'b00101110101: data <= 32'h374f3db6;
    11'b00101110110: data <= 32'ha6dd4118;
    11'b00101110111: data <= 32'hbcb33d89;
    11'b00101111000: data <= 32'hbdf7b6cd;
    11'b00101111001: data <= 32'hbb2eb87b;
    11'b00101111010: data <= 32'hb6123999;
    11'b00101111011: data <= 32'h0dd53c86;
    11'b00101111100: data <= 32'h3c112c60;
    11'b00101111101: data <= 32'h4094b992;
    11'b00101111110: data <= 32'h406b30cc;
    11'b00101111111: data <= 32'h374b3d9b;
    11'b00110000000: data <= 32'hbbf53cff;
    11'b00110000001: data <= 32'hb7faaf1b;
    11'b00110000010: data <= 32'h3aa1bc98;
    11'b00110000011: data <= 32'h3a67bda7;
    11'b00110000100: data <= 32'hb803be8a;
    11'b00110000101: data <= 32'hbb6ebf3b;
    11'b00110000110: data <= 32'h34cebc07;
    11'b00110000111: data <= 32'h3d3d38eb;
    11'b00110001000: data <= 32'h363c3d77;
    11'b00110001001: data <= 32'hbe0536d1;
    11'b00110001010: data <= 32'hc092b963;
    11'b00110001011: data <= 32'hbe82b366;
    11'b00110001100: data <= 32'hba913bd3;
    11'b00110001101: data <= 32'hb6603b34;
    11'b00110001110: data <= 32'h34e1b782;
    11'b00110001111: data <= 32'h3d29bb2c;
    11'b00110010000: data <= 32'h3da4398c;
    11'b00110010001: data <= 32'h35b040e9;
    11'b00110010010: data <= 32'hb6be4071;
    11'b00110010011: data <= 32'h31943703;
    11'b00110010100: data <= 32'h3c29babd;
    11'b00110010101: data <= 32'h38a9bbb1;
    11'b00110010110: data <= 32'hb884bbb2;
    11'b00110010111: data <= 32'hb553bd39;
    11'b00110011000: data <= 32'h3dbbbc9b;
    11'b00110011001: data <= 32'h40bbb2d5;
    11'b00110011010: data <= 32'h3b2d35e0;
    11'b00110011011: data <= 32'hbdc7b073;
    11'b00110011100: data <= 32'hc075b98c;
    11'b00110011101: data <= 32'hbd7ab229;
    11'b00110011110: data <= 32'hb938381b;
    11'b00110011111: data <= 32'hba43ade5;
    11'b00110100000: data <= 32'hb9bfbdb7;
    11'b00110100001: data <= 32'h2dedbd06;
    11'b00110100010: data <= 32'h39493b98;
    11'b00110100011: data <= 32'h341541b7;
    11'b00110100100: data <= 32'hb45a40ce;
    11'b00110100101: data <= 32'ha16a3876;
    11'b00110100110: data <= 32'h35d6b53e;
    11'b00110100111: data <= 32'hb0472f5c;
    11'b00110101000: data <= 32'hb9c23457;
    11'b00110101001: data <= 32'h32a9b86c;
    11'b00110101010: data <= 32'h4077bc96;
    11'b00110101011: data <= 32'h41dbb8de;
    11'b00110101100: data <= 32'h3cd531b9;
    11'b00110101101: data <= 32'hbbb63078;
    11'b00110101110: data <= 32'hbd33b48f;
    11'b00110101111: data <= 32'hb485b393;
    11'b00110110000: data <= 32'ha998b2ba;
    11'b00110110001: data <= 32'hbbf5bc88;
    11'b00110110010: data <= 32'hbdc9c073;
    11'b00110110011: data <= 32'hb803be87;
    11'b00110110100: data <= 32'h387f393b;
    11'b00110110101: data <= 32'h36814088;
    11'b00110110110: data <= 32'hb6f13e8c;
    11'b00110110111: data <= 32'hba313217;
    11'b00110111000: data <= 32'hb9bd2fef;
    11'b00110111001: data <= 32'hbbba3ca7;
    11'b00110111010: data <= 32'hbc113cec;
    11'b00110111011: data <= 32'h3275b14a;
    11'b00110111100: data <= 32'h402dbcb4;
    11'b00110111101: data <= 32'h412db7c4;
    11'b00110111110: data <= 32'h3c7f3a8a;
    11'b00110111111: data <= 32'hb5533c55;
    11'b00111000000: data <= 32'hab4c3681;
    11'b00111000001: data <= 32'h3b4cb096;
    11'b00111000010: data <= 32'h380ab853;
    11'b00111000011: data <= 32'hbc39bdc0;
    11'b00111000100: data <= 32'hbe2cc0a0;
    11'b00111000101: data <= 32'hb103bf34;
    11'b00111000110: data <= 32'h3cf3a9ca;
    11'b00111000111: data <= 32'h3aec3c13;
    11'b00111001000: data <= 32'hb8c1368d;
    11'b00111001001: data <= 32'hbdb4b5d3;
    11'b00111001010: data <= 32'hbd8e3574;
    11'b00111001011: data <= 32'hbd753e6f;
    11'b00111001100: data <= 32'hbd4c3d3a;
    11'b00111001101: data <= 32'hb6d5b7fe;
    11'b00111001110: data <= 32'h3c1ebda0;
    11'b00111001111: data <= 32'h3e2ab036;
    11'b00111010000: data <= 32'h39c63ec9;
    11'b00111010001: data <= 32'h2f253ff5;
    11'b00111010010: data <= 32'h3a253b98;
    11'b00111010011: data <= 32'h3dc1302f;
    11'b00111010100: data <= 32'h3825b046;
    11'b00111010101: data <= 32'hbc84b9b0;
    11'b00111010110: data <= 32'hbc95be5c;
    11'b00111010111: data <= 32'h3a2cbea4;
    11'b00111011000: data <= 32'h406db9e3;
    11'b00111011001: data <= 32'h3d94afa3;
    11'b00111011010: data <= 32'hb815b7a6;
    11'b00111011011: data <= 32'hbd80b928;
    11'b00111011100: data <= 32'hbc5435d6;
    11'b00111011101: data <= 32'hbc0e3d62;
    11'b00111011110: data <= 32'hbdd23858;
    11'b00111011111: data <= 32'hbd42bd75;
    11'b00111100000: data <= 32'hb4b5bf3b;
    11'b00111100001: data <= 32'h37742abb;
    11'b00111100010: data <= 32'h35584020;
    11'b00111100011: data <= 32'h32fc4040;
    11'b00111100100: data <= 32'h3a453b70;
    11'b00111100101: data <= 32'h3c1136f8;
    11'b00111100110: data <= 32'had333a90;
    11'b00111100111: data <= 32'hbd593917;
    11'b00111101000: data <= 32'hb9b9b824;
    11'b00111101001: data <= 32'h3e06bd65;
    11'b00111101010: data <= 32'h4179bc3e;
    11'b00111101011: data <= 32'h3e72b807;
    11'b00111101100: data <= 32'hb20ab7ab;
    11'b00111101101: data <= 32'hb860b61b;
    11'b00111101110: data <= 32'h2ee135f5;
    11'b00111101111: data <= 32'hae723a1b;
    11'b00111110000: data <= 32'hbd69b668;
    11'b00111110001: data <= 32'hbfcdc040;
    11'b00111110010: data <= 32'hbc4fc043;
    11'b00111110011: data <= 32'h2c09b05c;
    11'b00111110100: data <= 32'h34da3e30;
    11'b00111110101: data <= 32'h2e2a3d12;
    11'b00111110110: data <= 32'h31ed3483;
    11'b00111110111: data <= 32'h2c1938a6;
    11'b00111111000: data <= 32'hbb053f0e;
    11'b00111111001: data <= 32'hbe7d3f1c;
    11'b00111111010: data <= 32'hb956323a;
    11'b00111111011: data <= 32'h3da4bca2;
    11'b00111111100: data <= 32'h40a4bba8;
    11'b00111111101: data <= 32'h3d1ea9e9;
    11'b00111111110: data <= 32'h310034d6;
    11'b00111111111: data <= 32'h38b5343c;
    11'b01000000000: data <= 32'h3de937c9;
    11'b01000000001: data <= 32'h3a4c36da;
    11'b01000000010: data <= 32'hbca5b9d8;
    11'b01000000011: data <= 32'hc015c04e;
    11'b01000000100: data <= 32'hbb64c031;
    11'b01000000101: data <= 32'h3857b8a2;
    11'b01000000110: data <= 32'h39943678;
    11'b01000000111: data <= 32'ha5bcb01e;
    11'b01000001000: data <= 32'hb6d5b8f4;
    11'b01000001001: data <= 32'hb8dc3825;
    11'b01000001010: data <= 32'hbcf2405d;
    11'b01000001011: data <= 32'hbf17401a;
    11'b01000001100: data <= 32'hbc502dd6;
    11'b01000001101: data <= 32'h372abd2d;
    11'b01000001110: data <= 32'h3c75b937;
    11'b01000001111: data <= 32'h38413a0b;
    11'b01000010000: data <= 32'h34da3cb8;
    11'b01000010001: data <= 32'h3d7a3a45;
    11'b01000010010: data <= 32'h406b393b;
    11'b01000010011: data <= 32'h3c43394d;
    11'b01000010100: data <= 32'hbc6cadc6;
    11'b01000010101: data <= 32'hbec3bd29;
    11'b01000010110: data <= 32'hae8abe7e;
    11'b01000010111: data <= 32'h3dd8bbbb;
    11'b01000011000: data <= 32'h3cd7b96a;
    11'b01000011001: data <= 32'h0f8cbcec;
    11'b01000011010: data <= 32'hb802bccc;
    11'b01000011011: data <= 32'hb6013606;
    11'b01000011100: data <= 32'hba283fd3;
    11'b01000011101: data <= 32'hbe653dae;
    11'b01000011110: data <= 32'hbeacb97b;
    11'b01000011111: data <= 32'hba7bbeb6;
    11'b01000100000: data <= 32'hb1c2b71a;
    11'b01000100001: data <= 32'hb1fe3ccf;
    11'b01000100010: data <= 32'h329f3d83;
    11'b01000100011: data <= 32'h3da43964;
    11'b01000100100: data <= 32'h3fc7398e;
    11'b01000100101: data <= 32'h38b83d59;
    11'b01000100110: data <= 32'hbd243cbe;
    11'b01000100111: data <= 32'hbd0d9279;
    11'b01000101000: data <= 32'h395ebba9;
    11'b01000101001: data <= 32'h400fbc36;
    11'b01000101010: data <= 32'h3d74bc4b;
    11'b01000101011: data <= 32'h2ea0bda6;
    11'b01000101100: data <= 32'h2ce2bc68;
    11'b01000101101: data <= 32'h39ef3562;
    11'b01000101110: data <= 32'h359e3d94;
    11'b01000101111: data <= 32'hbc893793;
    11'b01000110000: data <= 32'hc014bde8;
    11'b01000110001: data <= 32'hbe5ebfda;
    11'b01000110010: data <= 32'hba4cb75f;
    11'b01000110011: data <= 32'hb6dd3b3b;
    11'b01000110100: data <= 32'h201d38ba;
    11'b01000110101: data <= 32'h3ac0b144;
    11'b01000110110: data <= 32'h3c1837b5;
    11'b01000110111: data <= 32'hb2f44000;
    11'b01000111000: data <= 32'hbe3540a1;
    11'b01000111001: data <= 32'hbc5a3b7c;
    11'b01000111010: data <= 32'h3a14b812;
    11'b01000111011: data <= 32'h3ebdbaaf;
    11'b01000111100: data <= 32'h3ae9b937;
    11'b01000111101: data <= 32'h2ee8b995;
    11'b01000111110: data <= 32'h3b72b78a;
    11'b01000111111: data <= 32'h402f3718;
    11'b01001000000: data <= 32'h3de93bca;
    11'b01001000001: data <= 32'hb9259f2e;
    11'b01001000010: data <= 32'hbfeabe4f;
    11'b01001000011: data <= 32'hbde4bf26;
    11'b01001000100: data <= 32'hb692b8ba;
    11'b01001000101: data <= 32'had9f287f;
    11'b01001000110: data <= 32'haf96ba41;
    11'b01001000111: data <= 32'h31cbbd41;
    11'b01001001000: data <= 32'h33872d9e;
    11'b01001001001: data <= 32'hb9334077;
    11'b01001001010: data <= 32'hbe63413d;
    11'b01001001011: data <= 32'hbce33bc4;
    11'b01001001100: data <= 32'h2b85b862;
    11'b01001001101: data <= 32'h380fb813;
    11'b01001001110: data <= 32'hb041318a;
    11'b01001001111: data <= 32'hae363430;
    11'b01001010000: data <= 32'h3dfe2f90;
    11'b01001010001: data <= 32'h41b53853;
    11'b01001010010: data <= 32'h3fb83bc8;
    11'b01001010011: data <= 32'hb7113634;
    11'b01001010100: data <= 32'hbe54ba05;
    11'b01001010101: data <= 32'hb92bbc4d;
    11'b01001010110: data <= 32'h386db8ec;
    11'b01001010111: data <= 32'h37c0ba83;
    11'b01001011000: data <= 32'hb063bfa6;
    11'b01001011001: data <= 32'had72c034;
    11'b01001011010: data <= 32'h33c2b3f8;
    11'b01001011011: data <= 32'hb3833fbc;
    11'b01001011100: data <= 32'hbcd23ffc;
    11'b01001011101: data <= 32'hbdcf31ee;
    11'b01001011110: data <= 32'hbba2bbc3;
    11'b01001011111: data <= 32'hba86b472;
    11'b01001100000: data <= 32'hbc5c3a2d;
    11'b01001100001: data <= 32'hb6fd394a;
    11'b01001100010: data <= 32'h3dbf2cb3;
    11'b01001100011: data <= 32'h4137364d;
    11'b01001100100: data <= 32'h3df03d38;
    11'b01001100101: data <= 32'hb90b3da7;
    11'b01001100110: data <= 32'hbc8e387e;
    11'b01001100111: data <= 32'h33d7b0c2;
    11'b01001101000: data <= 32'h3d33b6a6;
    11'b01001101001: data <= 32'h39b4bc51;
    11'b01001101010: data <= 32'hb1eec041;
    11'b01001101011: data <= 32'h31aac028;
    11'b01001101100: data <= 32'h3c70b516;
    11'b01001101101: data <= 32'h3b373d6b;
    11'b01001101110: data <= 32'hb77d3bad;
    11'b01001101111: data <= 32'hbe03ba12;
    11'b01001110000: data <= 32'hbe51bd5a;
    11'b01001110001: data <= 32'hbddeb1b3;
    11'b01001110010: data <= 32'hbdd23a0e;
    11'b01001110011: data <= 32'hb9b12f9f;
    11'b01001110100: data <= 32'h3abdba25;
    11'b01001110101: data <= 32'h3e7dada0;
    11'b01001110110: data <= 32'h386a3e82;
    11'b01001110111: data <= 32'hbbda40b9;
    11'b01001111000: data <= 32'hbb053e36;
    11'b01001111001: data <= 32'h38af3788;
    11'b01001111010: data <= 32'h3cc5ac75;
    11'b01001111011: data <= 32'h3347b8e8;
    11'b01001111100: data <= 32'hb6f8bd7e;
    11'b01001111101: data <= 32'h3978bd6d;
    11'b01001111110: data <= 32'h4087b04b;
    11'b01001111111: data <= 32'h402e3afd;
    11'b01010000000: data <= 32'h338d3422;
    11'b01010000001: data <= 32'hbd0bbc5c;
    11'b01010000010: data <= 32'hbd92bcc9;
    11'b01010000011: data <= 32'hbc4face7;
    11'b01010000100: data <= 32'hbc453369;
    11'b01010000101: data <= 32'hba3fbc31;
    11'b01010000110: data <= 32'h3064bfec;
    11'b01010000111: data <= 32'h3926b9d2;
    11'b01010001000: data <= 32'haeb43e87;
    11'b01010001001: data <= 32'hbc544128;
    11'b01010001010: data <= 32'hba7a3e64;
    11'b01010001011: data <= 32'h32ef36f8;
    11'b01010001100: data <= 32'h334d336c;
    11'b01010001101: data <= 32'hbaa533de;
    11'b01010001110: data <= 32'hbb45b40d;
    11'b01010001111: data <= 32'h3be3b874;
    11'b01010010000: data <= 32'h41d6290e;
    11'b01010010001: data <= 32'h412639a0;
    11'b01010010010: data <= 32'h37ea3561;
    11'b01010010011: data <= 32'hbac6b7cd;
    11'b01010010100: data <= 32'hb83fb6ee;
    11'b01010010101: data <= 32'h248531b0;
    11'b01010010110: data <= 32'hb4e4b530;
    11'b01010010111: data <= 32'hb9aec01c;
    11'b01010011000: data <= 32'hb43cc1a6;
    11'b01010011001: data <= 32'h35a7bcb3;
    11'b01010011010: data <= 32'h2d1b3d11;
    11'b01010011011: data <= 32'hb9463fa5;
    11'b01010011100: data <= 32'hba1939b0;
    11'b01010011101: data <= 32'hb7beb0a8;
    11'b01010011110: data <= 32'hbbac35f9;
    11'b01010011111: data <= 32'hbf763b9e;
    11'b01010100000: data <= 32'hbda436bf;
    11'b01010100001: data <= 32'h3a7eb5cd;
    11'b01010100010: data <= 32'h413daf2a;
    11'b01010100011: data <= 32'h401e3a2c;
    11'b01010100100: data <= 32'h31ee3c27;
    11'b01010100101: data <= 32'hb7b5396b;
    11'b01010100110: data <= 32'h372a38af;
    11'b01010100111: data <= 32'h3c1138af;
    11'b01010101000: data <= 32'h3150b6e9;
    11'b01010101001: data <= 32'hb9dfc06b;
    11'b01010101010: data <= 32'hb3c3c187;
    11'b01010101011: data <= 32'h3b27bcae;
    11'b01010101100: data <= 32'h3c3439f5;
    11'b01010101101: data <= 32'h31923a66;
    11'b01010101110: data <= 32'hb88db76a;
    11'b01010101111: data <= 32'hbb47ba0a;
    11'b01010110000: data <= 32'hbe2c36c8;
    11'b01010110001: data <= 32'hc0763c99;
    11'b01010110010: data <= 32'hbea9327a;
    11'b01010110011: data <= 32'h33cfbc15;
    11'b01010110100: data <= 32'h3e44b974;
    11'b01010110101: data <= 32'h3b5c3aa2;
    11'b01010110110: data <= 32'hb6603f04;
    11'b01010110111: data <= 32'hb49b3e5f;
    11'b01010111000: data <= 32'h3bcd3cf9;
    11'b01010111001: data <= 32'h3ce83bc4;
    11'b01010111010: data <= 32'hafa129ae;
    11'b01010111011: data <= 32'hbc38bd95;
    11'b01010111100: data <= 32'ha0a5bf79;
    11'b01010111101: data <= 32'h3f29ba2a;
    11'b01010111110: data <= 32'h404e3576;
    11'b01010111111: data <= 32'h3b97ac3e;
    11'b01011000000: data <= 32'hb350bc6c;
    11'b01011000001: data <= 32'hb95fbaa7;
    11'b01011000010: data <= 32'hbc633896;
    11'b01011000011: data <= 32'hbed23b28;
    11'b01011000100: data <= 32'hbe32b980;
    11'b01011000101: data <= 32'hb61ac046;
    11'b01011000110: data <= 32'h3715bda9;
    11'b01011000111: data <= 32'ha91e3975;
    11'b01011001000: data <= 32'hb9e43f81;
    11'b01011001001: data <= 32'hb25e3e57;
    11'b01011001010: data <= 32'h3af03c74;
    11'b01011001011: data <= 32'h386d3c85;
    11'b01011001100: data <= 32'hbc443aab;
    11'b01011001101: data <= 32'hbe8bb0bc;
    11'b01011001110: data <= 32'h2e74ba35;
    11'b01011001111: data <= 32'h409fb588;
    11'b01011010000: data <= 32'h412d31b8;
    11'b01011010001: data <= 32'h3ca2b38e;
    11'b01011010010: data <= 32'h2e24ba74;
    11'b01011010011: data <= 32'h3086b255;
    11'b01011010100: data <= 32'h2f073b82;
    11'b01011010101: data <= 32'hb960387e;
    11'b01011010110: data <= 32'hbce2be21;
    11'b01011010111: data <= 32'hba00c1de;
    11'b01011011000: data <= 32'had15bf6f;
    11'b01011011001: data <= 32'hb17d359b;
    11'b01011011010: data <= 32'hb77d3ceb;
    11'b01011011011: data <= 32'haa3538cb;
    11'b01011011100: data <= 32'h369234a1;
    11'b01011011101: data <= 32'hb71b3c17;
    11'b01011011110: data <= 32'hc01c3df4;
    11'b01011011111: data <= 32'hc05939ee;
    11'b01011100000: data <= 32'hae2bb418;
    11'b01011100001: data <= 32'h4001b501;
    11'b01011100010: data <= 32'h3ff1312a;
    11'b01011100011: data <= 32'h392032b1;
    11'b01011100100: data <= 32'h33803094;
    11'b01011100101: data <= 32'h3c3f3a30;
    11'b01011100110: data <= 32'h3d3a3dae;
    11'b01011100111: data <= 32'h302a383d;
    11'b01011101000: data <= 32'hbc21be97;
    11'b01011101001: data <= 32'hba4ec19b;
    11'b01011101010: data <= 32'h3267bec0;
    11'b01011101011: data <= 32'h3879259d;
    11'b01011101100: data <= 32'h34e9318a;
    11'b01011101101: data <= 32'h33daba14;
    11'b01011101110: data <= 32'h2ef5b932;
    11'b01011101111: data <= 32'hbbb33ab3;
    11'b01011110000: data <= 32'hc0bd3ee1;
    11'b01011110001: data <= 32'hc0a03a40;
    11'b01011110010: data <= 32'hb818b932;
    11'b01011110011: data <= 32'h3bf8ba6e;
    11'b01011110100: data <= 32'h39682eb2;
    11'b01011110101: data <= 32'hb4393a16;
    11'b01011110110: data <= 32'h31b13bba;
    11'b01011110111: data <= 32'h3e663d95;
    11'b01011111000: data <= 32'h3f173ef7;
    11'b01011111001: data <= 32'h30453b38;
    11'b01011111010: data <= 32'hbcfcbaed;
    11'b01011111011: data <= 32'hb95abf02;
    11'b01011111100: data <= 32'h3b36bbdf;
    11'b01011111101: data <= 32'h3e2ab012;
    11'b01011111110: data <= 32'h3c3cb97e;
    11'b01011111111: data <= 32'h3898be9d;
    11'b01100000000: data <= 32'h34bcbc25;
    11'b01100000001: data <= 32'hb8443aca;
    11'b01100000010: data <= 32'hbed83e46;
    11'b01100000011: data <= 32'hbfaf2edf;
    11'b01100000100: data <= 32'hbb1fbe78;
    11'b01100000101: data <= 32'haf14be13;
    11'b01100000110: data <= 32'hb841acc9;
    11'b01100000111: data <= 32'hbb763b0c;
    11'b01100001000: data <= 32'h2e3c3ba8;
    11'b01100001001: data <= 32'h3e533ca5;
    11'b01100001010: data <= 32'h3d523eaa;
    11'b01100001011: data <= 32'hb91c3ddb;
    11'b01100001100: data <= 32'hbf3735bb;
    11'b01100001101: data <= 32'hb900b6b3;
    11'b01100001110: data <= 32'h3d7fb2ca;
    11'b01100001111: data <= 32'h3fd3adc4;
    11'b01100010000: data <= 32'h3cc3bb6f;
    11'b01100010001: data <= 32'h39b8be66;
    11'b01100010010: data <= 32'h3b4fb8dd;
    11'b01100010011: data <= 32'h39303cb6;
    11'b01100010100: data <= 32'hb7313d4c;
    11'b01100010101: data <= 32'hbcf6b930;
    11'b01100010110: data <= 32'hbc23c0c0;
    11'b01100010111: data <= 32'hb982bfa4;
    11'b01100011000: data <= 32'hbb62b46d;
    11'b01100011001: data <= 32'hbb3b363b;
    11'b01100011010: data <= 32'h32189fb0;
    11'b01100011011: data <= 32'h3ce73011;
    11'b01100011100: data <= 32'h374a3cdb;
    11'b01100011101: data <= 32'hbe493f84;
    11'b01100011110: data <= 32'hc0a13d26;
    11'b01100011111: data <= 32'hb9f435f5;
    11'b01100100000: data <= 32'h3cb52e34;
    11'b01100100001: data <= 32'h3d79a51e;
    11'b01100100010: data <= 32'h37d0b8b9;
    11'b01100100011: data <= 32'h383fba6e;
    11'b01100100100: data <= 32'h3e5e3492;
    11'b01100100101: data <= 32'h3f7e3e98;
    11'b01100100110: data <= 32'h390b3d0c;
    11'b01100100111: data <= 32'hb9edbaab;
    11'b01100101000: data <= 32'hbb99c082;
    11'b01100101001: data <= 32'hb819be56;
    11'b01100101010: data <= 32'hb603b50c;
    11'b01100101011: data <= 32'hb380b6fa;
    11'b01100101100: data <= 32'h37b4bd8c;
    11'b01100101101: data <= 32'h3b7bbc5d;
    11'b01100101110: data <= 32'hadf23988;
    11'b01100101111: data <= 32'hbf913fd0;
    11'b01100110000: data <= 32'hc0a93db1;
    11'b01100110001: data <= 32'hbb4a321b;
    11'b01100110010: data <= 32'h361bb40b;
    11'b01100110011: data <= 32'h297dac71;
    11'b01100110100: data <= 32'hb98aad57;
    11'b01100110101: data <= 32'h2fb52145;
    11'b01100110110: data <= 32'h3fc83b4c;
    11'b01100110111: data <= 32'h40d93f8a;
    11'b01100111000: data <= 32'h3af93dbc;
    11'b01100111001: data <= 32'hba30b3a4;
    11'b01100111010: data <= 32'hba72bcc5;
    11'b01100111011: data <= 32'h2fbbb8eb;
    11'b01100111100: data <= 32'h387baec7;
    11'b01100111101: data <= 32'h3818bc60;
    11'b01100111110: data <= 32'h3a14c0b8;
    11'b01100111111: data <= 32'h3bc9bef6;
    11'b01101000000: data <= 32'h31ae37ab;
    11'b01101000001: data <= 32'hbceb3f03;
    11'b01101000010: data <= 32'hbec73aa5;
    11'b01101000011: data <= 32'hbb81b991;
    11'b01101000100: data <= 32'hb81bbb91;
    11'b01101000101: data <= 32'hbcf6b334;
    11'b01101000110: data <= 32'hbe943058;
    11'b01101000111: data <= 32'hb3323024;
    11'b01101001000: data <= 32'h3f653975;
    11'b01101001001: data <= 32'h40253e64;
    11'b01101001010: data <= 32'h32e63ea8;
    11'b01101001011: data <= 32'hbd233a2c;
    11'b01101001100: data <= 32'hba0732ce;
    11'b01101001101: data <= 32'h392f3756;
    11'b01101001110: data <= 32'h3c483378;
    11'b01101001111: data <= 32'h3944bceb;
    11'b01101010000: data <= 32'h39d1c0ce;
    11'b01101010001: data <= 32'h3d2bbddb;
    11'b01101010010: data <= 32'h3c9b39d9;
    11'b01101010011: data <= 32'h2e383e04;
    11'b01101010100: data <= 32'hb9a12b10;
    11'b01101010101: data <= 32'hb9ffbe12;
    11'b01101010110: data <= 32'hbbabbd6e;
    11'b01101010111: data <= 32'hbef0b4b7;
    11'b01101011000: data <= 32'hbf3aae55;
    11'b01101011001: data <= 32'hb3eab91d;
    11'b01101011010: data <= 32'h3defb67f;
    11'b01101011011: data <= 32'h3cd43ab6;
    11'b01101011100: data <= 32'hba013eea;
    11'b01101011101: data <= 32'hbf443e2f;
    11'b01101011110: data <= 32'hba3a3c73;
    11'b01101011111: data <= 32'h39503bfd;
    11'b01101100000: data <= 32'h394c376c;
    11'b01101100001: data <= 32'had6ebaf0;
    11'b01101100010: data <= 32'h340ebe90;
    11'b01101100011: data <= 32'h3e77b88e;
    11'b01101100100: data <= 32'h40693cdf;
    11'b01101100101: data <= 32'h3d293d84;
    11'b01101100110: data <= 32'h2c22b4ce;
    11'b01101100111: data <= 32'hb74ebe3b;
    11'b01101101000: data <= 32'hb9ebbc06;
    11'b01101101001: data <= 32'hbcfaac8a;
    11'b01101101010: data <= 32'hbcb3b8a3;
    11'b01101101011: data <= 32'h2a0dbf5d;
    11'b01101101100: data <= 32'h3c9fbef3;
    11'b01101101101: data <= 32'h38362492;
    11'b01101101110: data <= 32'hbcdc3e32;
    11'b01101101111: data <= 32'hbf4d3e76;
    11'b01101110000: data <= 32'hb9bc3c09;
    11'b01101110001: data <= 32'h322c39d9;
    11'b01101110010: data <= 32'hb7c036f9;
    11'b01101110011: data <= 32'hbd81b56e;
    11'b01101110100: data <= 32'hb795b9da;
    11'b01101110101: data <= 32'h3eb731dd;
    11'b01101110110: data <= 32'h41563dde;
    11'b01101110111: data <= 32'h3e823d71;
    11'b01101111000: data <= 32'h31329b38;
    11'b01101111001: data <= 32'hb414b962;
    11'b01101111010: data <= 32'hadd32c39;
    11'b01101111011: data <= 32'hb3f1376a;
    11'b01101111100: data <= 32'hb533bb60;
    11'b01101111101: data <= 32'h35aac16a;
    11'b01101111110: data <= 32'h3c2dc100;
    11'b01101111111: data <= 32'h383cb5fa;
    11'b01110000000: data <= 32'hb9d53cfc;
    11'b01110000001: data <= 32'hbc673c03;
    11'b01110000010: data <= 32'hb6c32e02;
    11'b01110000011: data <= 32'hb5f6a894;
    11'b01110000100: data <= 32'hbe9a33d8;
    11'b01110000101: data <= 32'hc0eba051;
    11'b01110000110: data <= 32'hbc2db60a;
    11'b01110000111: data <= 32'h3dbd3020;
    11'b01110001000: data <= 32'h40923c74;
    11'b01110001001: data <= 32'h3bc73d25;
    11'b01110001010: data <= 32'hb62b3962;
    11'b01110001011: data <= 32'hb36b38d9;
    11'b01110001100: data <= 32'h38243d21;
    11'b01110001101: data <= 32'h37673c47;
    11'b01110001110: data <= 32'h9e64baf0;
    11'b01110001111: data <= 32'h3487c16b;
    11'b01110010000: data <= 32'h3c58c082;
    11'b01110010001: data <= 32'h3cb2b019;
    11'b01110010010: data <= 32'h37673c08;
    11'b01110010011: data <= 32'h291c3156;
    11'b01110010100: data <= 32'h2c4abb2a;
    11'b01110010101: data <= 32'hb8b4b8e6;
    11'b01110010110: data <= 32'hc03031f8;
    11'b01110010111: data <= 32'hc15e97e9;
    11'b01110011000: data <= 32'hbc7dbaa3;
    11'b01110011001: data <= 32'h3c37ba84;
    11'b01110011010: data <= 32'h3d7c32af;
    11'b01110011011: data <= 32'hb0303c1c;
    11'b01110011100: data <= 32'hbc473cbc;
    11'b01110011101: data <= 32'hb4473dca;
    11'b01110011110: data <= 32'h39e73fae;
    11'b01110011111: data <= 32'h35a33da3;
    11'b01110100000: data <= 32'hb8c2b74a;
    11'b01110100001: data <= 32'hb528bf9f;
    11'b01110100010: data <= 32'h3c52bd04;
    11'b01110100011: data <= 32'h3fc337e2;
    11'b01110100100: data <= 32'h3e5a3b45;
    11'b01110100101: data <= 32'h3b7eb5c0;
    11'b01110100110: data <= 32'h3834bcdb;
    11'b01110100111: data <= 32'hb47cb6ca;
    11'b01110101000: data <= 32'hbe443828;
    11'b01110101001: data <= 32'hbfedb124;
    11'b01110101010: data <= 32'hb9c5beeb;
    11'b01110101011: data <= 32'h3a0ec023;
    11'b01110101100: data <= 32'h3864ba1f;
    11'b01110101101: data <= 32'hbad2390a;
    11'b01110101110: data <= 32'hbd013c7e;
    11'b01110101111: data <= 32'hafe63d3c;
    11'b01110110000: data <= 32'h38923e7e;
    11'b01110110001: data <= 32'hb7d13d41;
    11'b01110110010: data <= 32'hbf3329e4;
    11'b01110110011: data <= 32'hbcdebb07;
    11'b01110110100: data <= 32'h3b10b43b;
    11'b01110110101: data <= 32'h40783b5f;
    11'b01110110110: data <= 32'h3f913ab3;
    11'b01110110111: data <= 32'h3c32b583;
    11'b01110111000: data <= 32'h39adb913;
    11'b01110111001: data <= 32'h35ba3868;
    11'b01110111010: data <= 32'hb7943ce7;
    11'b01110111011: data <= 32'hbb59b2c9;
    11'b01110111100: data <= 32'hb369c0ca;
    11'b01110111101: data <= 32'h38f6c199;
    11'b01110111110: data <= 32'h34bbbcdb;
    11'b01110111111: data <= 32'hb95f349d;
    11'b01111000000: data <= 32'hb91a37ec;
    11'b01111000001: data <= 32'h35673507;
    11'b01111000010: data <= 32'h35083965;
    11'b01111000011: data <= 32'hbdb63b94;
    11'b01111000100: data <= 32'hc1b4360c;
    11'b01111000101: data <= 32'hbf8bb4bb;
    11'b01111000110: data <= 32'h3856a44c;
    11'b01111000111: data <= 32'h3f373999;
    11'b01111001000: data <= 32'h3caf38e4;
    11'b01111001001: data <= 32'h35b623b9;
    11'b01111001010: data <= 32'h389e3662;
    11'b01111001011: data <= 32'h3ba03ef3;
    11'b01111001100: data <= 32'h37083fde;
    11'b01111001101: data <= 32'hb4db9f95;
    11'b01111001110: data <= 32'hb0bec0a2;
    11'b01111001111: data <= 32'h384ac100;
    11'b01111010000: data <= 32'h38ffbaf0;
    11'b01111010001: data <= 32'h3423318e;
    11'b01111010010: data <= 32'h377eb533;
    11'b01111010011: data <= 32'h3beebad4;
    11'b01111010100: data <= 32'h34c1b201;
    11'b01111010101: data <= 32'hbf0c39b7;
    11'b01111010110: data <= 32'hc21337b0;
    11'b01111010111: data <= 32'hbfa3b717;
    11'b01111011000: data <= 32'h33c4b978;
    11'b01111011001: data <= 32'h3b2eb113;
    11'b01111011010: data <= 32'hadc13177;
    11'b01111011011: data <= 32'hb8c7349d;
    11'b01111011100: data <= 32'h35af3c6a;
    11'b01111011101: data <= 32'h3cf540b4;
    11'b01111011110: data <= 32'h38f1409b;
    11'b01111011111: data <= 32'hb8d435f3;
    11'b01111100000: data <= 32'hb97fbe07;
    11'b01111100001: data <= 32'h3584bd71;
    11'b01111100010: data <= 32'h3c7e16d3;
    11'b01111100011: data <= 32'h3ce43434;
    11'b01111100100: data <= 32'h3d6dbb27;
    11'b01111100101: data <= 32'h3dffbdc5;
    11'b01111100110: data <= 32'h3901b4c5;
    11'b01111100111: data <= 32'hbcd93ba6;
    11'b01111101000: data <= 32'hc06f37f6;
    11'b01111101001: data <= 32'hbd29bc39;
    11'b01111101010: data <= 32'h300cbf04;
    11'b01111101011: data <= 32'h2a36bc88;
    11'b01111101100: data <= 32'hbc45b534;
    11'b01111101101: data <= 32'hbc5630d6;
    11'b01111101110: data <= 32'h361a3b64;
    11'b01111101111: data <= 32'h3cec3fd9;
    11'b01111110000: data <= 32'h2cad400f;
    11'b01111110001: data <= 32'hbe6939b1;
    11'b01111110010: data <= 32'hbe55b768;
    11'b01111110011: data <= 32'h2151b027;
    11'b01111110100: data <= 32'h3d2839f0;
    11'b01111110101: data <= 32'h3dda355b;
    11'b01111110110: data <= 32'h3d9fbc0f;
    11'b01111110111: data <= 32'h3e39bca6;
    11'b01111111000: data <= 32'h3c883738;
    11'b01111111001: data <= 32'haec53ea0;
    11'b01111111010: data <= 32'hbb7238df;
    11'b01111111011: data <= 32'hb7d3be33;
    11'b01111111100: data <= 32'h30fcc0cd;
    11'b01111111101: data <= 32'hb518be2f;
    11'b01111111110: data <= 32'hbcbfb8c5;
    11'b01111111111: data <= 32'hb9bfb635;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    