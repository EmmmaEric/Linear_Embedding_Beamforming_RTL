
module memory_rom_8(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbe523145;
    11'b00000000001: data <= 32'hba892f92;
    11'b00000000010: data <= 32'h3c07a890;
    11'b00000000011: data <= 32'h3ee139fc;
    11'b00000000100: data <= 32'h32993ee8;
    11'b00000000101: data <= 32'hbeb03eb9;
    11'b00000000110: data <= 32'hbe1b3b52;
    11'b00000000111: data <= 32'h341a381e;
    11'b00000001000: data <= 32'h3d3c35c6;
    11'b00000001001: data <= 32'h3a7bb75d;
    11'b00000001010: data <= 32'h357abe23;
    11'b00000001011: data <= 32'h3c3dbd01;
    11'b00000001100: data <= 32'h3f823835;
    11'b00000001101: data <= 32'h3d723e90;
    11'b00000001110: data <= 32'ha4513816;
    11'b00000001111: data <= 32'hba90bde9;
    11'b00000010000: data <= 32'hbb0abf9a;
    11'b00000010001: data <= 32'hbc29b9e4;
    11'b00000010010: data <= 32'hbcdbaf52;
    11'b00000010011: data <= 32'hb787bb17;
    11'b00000010100: data <= 32'h3af9bda9;
    11'b00000010101: data <= 32'h3c28b4a4;
    11'b00000010110: data <= 32'hb88a3dd7;
    11'b00000010111: data <= 32'hc01e3ff4;
    11'b00000011000: data <= 32'hbe463d01;
    11'b00000011001: data <= 32'h26fd3884;
    11'b00000011010: data <= 32'h37a63534;
    11'b00000011011: data <= 32'hb659b0a0;
    11'b00000011100: data <= 32'hb846b9cc;
    11'b00000011101: data <= 32'h3c1db4f7;
    11'b00000011110: data <= 32'h41173c5c;
    11'b00000011111: data <= 32'h40413ee7;
    11'b00000100000: data <= 32'h3697386c;
    11'b00000100001: data <= 32'hb8fdbbf3;
    11'b00000100010: data <= 32'hb7d6bc22;
    11'b00000100011: data <= 32'hb3eeaf50;
    11'b00000100100: data <= 32'hb4cab528;
    11'b00000100101: data <= 32'h2c7cbf7d;
    11'b00000100110: data <= 32'h3ad2c11a;
    11'b00000100111: data <= 32'h3a6ebc01;
    11'b00000101000: data <= 32'hb8163cb4;
    11'b00000101001: data <= 32'hbe783ec9;
    11'b00000101010: data <= 32'hbcf0392d;
    11'b00000101011: data <= 32'hb59fb10d;
    11'b00000101100: data <= 32'hb970a8aa;
    11'b00000101101: data <= 32'hbefb2dd3;
    11'b00000101110: data <= 32'hbd90b181;
    11'b00000101111: data <= 32'h3a712954;
    11'b00000110000: data <= 32'h410e3c26;
    11'b00000110001: data <= 32'h3f853e85;
    11'b00000110010: data <= 32'h10b23bec;
    11'b00000110011: data <= 32'hb9ee3091;
    11'b00000110100: data <= 32'ha4113501;
    11'b00000110101: data <= 32'h38bb39c5;
    11'b00000110110: data <= 32'h35e8b45e;
    11'b00000110111: data <= 32'h3472c077;
    11'b00000111000: data <= 32'h3ae5c189;
    11'b00000111001: data <= 32'h3ca1bbb8;
    11'b00000111010: data <= 32'h36d43c49;
    11'b00000111011: data <= 32'hb7963c4b;
    11'b00000111100: data <= 32'hb89fb5c2;
    11'b00000111101: data <= 32'hb858bc04;
    11'b00000111110: data <= 32'hbdb3b56e;
    11'b00000111111: data <= 32'hc0da30da;
    11'b00001000000: data <= 32'hbeddb49e;
    11'b00001000001: data <= 32'h3873b885;
    11'b00001000010: data <= 32'h3faa330d;
    11'b00001000011: data <= 32'h3b353cfa;
    11'b00001000100: data <= 32'hbacf3dbd;
    11'b00001000101: data <= 32'hbbf53cc6;
    11'b00001000110: data <= 32'h340c3d5c;
    11'b00001000111: data <= 32'h3ab03d35;
    11'b00001001000: data <= 32'h317e1dbb;
    11'b00001001001: data <= 32'hb214bf38;
    11'b00001001010: data <= 32'h39d3c00f;
    11'b00001001011: data <= 32'h3f29b4a7;
    11'b00001001100: data <= 32'h3e9b3cad;
    11'b00001001101: data <= 32'h39be385f;
    11'b00001001110: data <= 32'h2d27bbff;
    11'b00001001111: data <= 32'hb604bce7;
    11'b00001010000: data <= 32'hbd3eb177;
    11'b00001010001: data <= 32'hc02a30c1;
    11'b00001010010: data <= 32'hbd71bbaa;
    11'b00001010011: data <= 32'h370fbf31;
    11'b00001010100: data <= 32'h3cb1bba2;
    11'b00001010101: data <= 32'haa4c397e;
    11'b00001010110: data <= 32'hbda33e10;
    11'b00001010111: data <= 32'hbc1b3de7;
    11'b00001011000: data <= 32'h34453dc6;
    11'b00001011001: data <= 32'h353b3d3a;
    11'b00001011010: data <= 32'hbb0d3532;
    11'b00001011011: data <= 32'hbccdbb95;
    11'b00001011100: data <= 32'h3621bb8a;
    11'b00001011101: data <= 32'h406436f3;
    11'b00001011110: data <= 32'h40b33d11;
    11'b00001011111: data <= 32'h3ced3614;
    11'b00001100000: data <= 32'h35f8ba8e;
    11'b00001100001: data <= 32'h2ac3b828;
    11'b00001100010: data <= 32'hb7ac389a;
    11'b00001100011: data <= 32'hbc373435;
    11'b00001100100: data <= 32'hb967bea0;
    11'b00001100101: data <= 32'h3740c1b5;
    11'b00001100110: data <= 32'h3a1abf1c;
    11'b00001100111: data <= 32'hb4733403;
    11'b00001101000: data <= 32'hbc8c3c92;
    11'b00001101001: data <= 32'hb8b13aae;
    11'b00001101010: data <= 32'h32a73926;
    11'b00001101011: data <= 32'hb83a3a9e;
    11'b00001101100: data <= 32'hc049382a;
    11'b00001101101: data <= 32'hc063b40b;
    11'b00001101110: data <= 32'ha97eb534;
    11'b00001101111: data <= 32'h401b387f;
    11'b00001110000: data <= 32'h40213c5e;
    11'b00001110001: data <= 32'h3a3e3815;
    11'b00001110010: data <= 32'h31a71fa8;
    11'b00001110011: data <= 32'h37dd39dd;
    11'b00001110100: data <= 32'h37983e42;
    11'b00001110101: data <= 32'hb0963878;
    11'b00001110110: data <= 32'hb477bf6a;
    11'b00001110111: data <= 32'h369cc211;
    11'b00001111000: data <= 32'h3aa8bef7;
    11'b00001111001: data <= 32'h358e31ad;
    11'b00001111010: data <= 32'hae49384e;
    11'b00001111011: data <= 32'h337ab446;
    11'b00001111100: data <= 32'h34c1b6b3;
    11'b00001111101: data <= 32'hbc4e3559;
    11'b00001111110: data <= 32'hc19238cd;
    11'b00001111111: data <= 32'hc11eaf34;
    11'b00010000000: data <= 32'hb504b8f7;
    11'b00010000001: data <= 32'h3dbdb052;
    11'b00010000010: data <= 32'h3c04385c;
    11'b00010000011: data <= 32'hb4233935;
    11'b00010000100: data <= 32'hb4233aa9;
    11'b00010000101: data <= 32'h3a0b3ee4;
    11'b00010000110: data <= 32'h3b924075;
    11'b00010000111: data <= 32'ha8773b52;
    11'b00010001000: data <= 32'hb8dbbd8c;
    11'b00010001001: data <= 32'h304dc072;
    11'b00010001010: data <= 32'h3c99bb4d;
    11'b00010001011: data <= 32'h3d4b370a;
    11'b00010001100: data <= 32'h3c3927ad;
    11'b00010001101: data <= 32'h3c0ebc6d;
    11'b00010001110: data <= 32'h38cabb81;
    11'b00010001111: data <= 32'hbb24357f;
    11'b00010010000: data <= 32'hc0c439bd;
    11'b00010010001: data <= 32'hc02db782;
    11'b00010010010: data <= 32'hb4aabe58;
    11'b00010010011: data <= 32'h39b6bd0f;
    11'b00010010100: data <= 32'hafe4b145;
    11'b00010010101: data <= 32'hbc6b385b;
    11'b00010010110: data <= 32'hb77a3c0b;
    11'b00010010111: data <= 32'h3ae43f22;
    11'b00010011000: data <= 32'h39e84054;
    11'b00010011001: data <= 32'hba773c8b;
    11'b00010011010: data <= 32'hbe3eb863;
    11'b00010011011: data <= 32'hb615bbd4;
    11'b00010011100: data <= 32'h3d4c2da5;
    11'b00010011101: data <= 32'h3f8c39d3;
    11'b00010011110: data <= 32'h3e28b26b;
    11'b00010011111: data <= 32'h3d29bcda;
    11'b00010100000: data <= 32'h3bd3b82a;
    11'b00010100001: data <= 32'hac533c11;
    11'b00010100010: data <= 32'hbcdf3c06;
    11'b00010100011: data <= 32'hbc95bb40;
    11'b00010100100: data <= 32'had3ec0f6;
    11'b00010100101: data <= 32'h343cc024;
    11'b00010100110: data <= 32'hb8fdb916;
    11'b00010100111: data <= 32'hbc853148;
    11'b00010101000: data <= 32'hafca35bb;
    11'b00010101001: data <= 32'h3bc43af0;
    11'b00010101010: data <= 32'h313a3dd5;
    11'b00010101011: data <= 32'hbf8a3c8d;
    11'b00010101100: data <= 32'hc1163148;
    11'b00010101101: data <= 32'hbb1baec8;
    11'b00010101110: data <= 32'h3c793832;
    11'b00010101111: data <= 32'h3e433962;
    11'b00010110000: data <= 32'h3bf5b32f;
    11'b00010110001: data <= 32'h3b3fb96d;
    11'b00010110010: data <= 32'h3cf73837;
    11'b00010110011: data <= 32'h3b233ffe;
    11'b00010110100: data <= 32'hac6f3db1;
    11'b00010110101: data <= 32'hb6f5bbe9;
    11'b00010110110: data <= 32'h26c8c132;
    11'b00010110111: data <= 32'h326bbfd9;
    11'b00010111000: data <= 32'hb4bbb88e;
    11'b00010111001: data <= 32'hb515b4bb;
    11'b00010111010: data <= 32'h397fb9f8;
    11'b00010111011: data <= 32'h3cd8b6a1;
    11'b00010111100: data <= 32'hb3383933;
    11'b00010111101: data <= 32'hc0e43c2d;
    11'b00010111110: data <= 32'hc1b9369c;
    11'b00010111111: data <= 32'hbc49ae92;
    11'b00011000000: data <= 32'h38d32cdb;
    11'b00011000001: data <= 32'h37f730d3;
    11'b00011000010: data <= 32'hb3ceb40f;
    11'b00011000011: data <= 32'h3152aa4a;
    11'b00011000100: data <= 32'h3d423dab;
    11'b00011000101: data <= 32'h3dca4147;
    11'b00011000110: data <= 32'h355c3efc;
    11'b00011000111: data <= 32'hb7d6b8a3;
    11'b00011001000: data <= 32'hb28cbf19;
    11'b00011001001: data <= 32'h3579bba7;
    11'b00011001010: data <= 32'h3740a5f5;
    11'b00011001011: data <= 32'h39bdb8e1;
    11'b00011001100: data <= 32'h3ddebe99;
    11'b00011001101: data <= 32'h3e23bce5;
    11'b00011001110: data <= 32'haa8d35d2;
    11'b00011001111: data <= 32'hc00a3c55;
    11'b00011010000: data <= 32'hc07b3342;
    11'b00011010001: data <= 32'hba5fba8a;
    11'b00011010010: data <= 32'h2c66bb4e;
    11'b00011010011: data <= 32'hb973b895;
    11'b00011010100: data <= 32'hbd7fb6e7;
    11'b00011010101: data <= 32'hb5b12dd8;
    11'b00011010110: data <= 32'h3d3f3dc8;
    11'b00011010111: data <= 32'h3d9540ea;
    11'b00011011000: data <= 32'hb1733f05;
    11'b00011011001: data <= 32'hbd1c2dd2;
    11'b00011011010: data <= 32'hb9e3b7c1;
    11'b00011011011: data <= 32'h367d3522;
    11'b00011011100: data <= 32'h3b7838ba;
    11'b00011011101: data <= 32'h3ca4b9a2;
    11'b00011011110: data <= 32'h3ea6bf96;
    11'b00011011111: data <= 32'h3f03bc5a;
    11'b00011100000: data <= 32'h390f3abd;
    11'b00011100001: data <= 32'hba853d85;
    11'b00011100010: data <= 32'hbc23ac98;
    11'b00011100011: data <= 32'hb418be59;
    11'b00011100100: data <= 32'hb320beaa;
    11'b00011100101: data <= 32'hbd3bbbfe;
    11'b00011100110: data <= 32'hbec6b9a9;
    11'b00011100111: data <= 32'hb37eb74b;
    11'b00011101000: data <= 32'h3da637ea;
    11'b00011101001: data <= 32'h3bcc3e09;
    11'b00011101010: data <= 32'hbc5c3dbb;
    11'b00011101011: data <= 32'hc063390e;
    11'b00011101100: data <= 32'hbceb3804;
    11'b00011101101: data <= 32'h33de3c40;
    11'b00011101110: data <= 32'h396c3a57;
    11'b00011101111: data <= 32'h38acb98f;
    11'b00011110000: data <= 32'h3c44be17;
    11'b00011110001: data <= 32'h3ed9b33c;
    11'b00011110010: data <= 32'h3da93ef9;
    11'b00011110011: data <= 32'h36fa3f38;
    11'b00011110100: data <= 32'h9fcdb0c7;
    11'b00011110101: data <= 32'h3086beed;
    11'b00011110110: data <= 32'hb335be1e;
    11'b00011110111: data <= 32'hbc92ba12;
    11'b00011111000: data <= 32'hbc60bb34;
    11'b00011111001: data <= 32'h378fbd8f;
    11'b00011111010: data <= 32'h3eb2bb08;
    11'b00011111011: data <= 32'h39113621;
    11'b00011111100: data <= 32'hbe8f3c17;
    11'b00011111101: data <= 32'hc0f83a4f;
    11'b00011111110: data <= 32'hbd1e3955;
    11'b00011111111: data <= 32'haa033ada;
    11'b00100000000: data <= 32'hb3963669;
    11'b00100000001: data <= 32'hb9e6ba00;
    11'b00100000010: data <= 32'h2411bbd0;
    11'b00100000011: data <= 32'h3dd038f5;
    11'b00100000100: data <= 32'h3f6840b8;
    11'b00100000101: data <= 32'h3bfa4012;
    11'b00100000110: data <= 32'h32aa2d95;
    11'b00100000111: data <= 32'h2cf5bc24;
    11'b00100001000: data <= 32'hae82b72f;
    11'b00100001001: data <= 32'hb80b2d4c;
    11'b00100001010: data <= 32'hb059bb08;
    11'b00100001011: data <= 32'h3ce9c050;
    11'b00100001100: data <= 32'h3fc8bf5c;
    11'b00100001101: data <= 32'h397db266;
    11'b00100001110: data <= 32'hbd453ad4;
    11'b00100001111: data <= 32'hbf3338d1;
    11'b00100010000: data <= 32'hb9de2d57;
    11'b00100010001: data <= 32'hb418a558;
    11'b00100010010: data <= 32'hbd16b4aa;
    11'b00100010011: data <= 32'hc007bb49;
    11'b00100010100: data <= 32'hba98ba1d;
    11'b00100010101: data <= 32'h3ccf39cf;
    11'b00100010110: data <= 32'h3f1a4041;
    11'b00100010111: data <= 32'h39183f3b;
    11'b00100011000: data <= 32'hb6e73744;
    11'b00100011001: data <= 32'hb67b2efc;
    11'b00100011010: data <= 32'ha9e83bc4;
    11'b00100011011: data <= 32'h8a173c1f;
    11'b00100011100: data <= 32'h35bfb989;
    11'b00100011101: data <= 32'h3d90c0b5;
    11'b00100011110: data <= 32'h3fe0bf6f;
    11'b00100011111: data <= 32'h3c642e04;
    11'b00100100000: data <= 32'hb4073c4c;
    11'b00100100001: data <= 32'hb752352b;
    11'b00100100010: data <= 32'h30c0b95d;
    11'b00100100011: data <= 32'hb3b2ba64;
    11'b00100100100: data <= 32'hbf4fb99c;
    11'b00100100101: data <= 32'hc0febc28;
    11'b00100100110: data <= 32'hbb66bc50;
    11'b00100100111: data <= 32'h3cc4adf5;
    11'b00100101000: data <= 32'h3d7f3c38;
    11'b00100101001: data <= 32'hb3783c97;
    11'b00100101010: data <= 32'hbd5f3960;
    11'b00100101011: data <= 32'hbb223c09;
    11'b00100101100: data <= 32'haeaa3f8c;
    11'b00100101101: data <= 32'hac643df8;
    11'b00100101110: data <= 32'hae2bb843;
    11'b00100101111: data <= 32'h3984bff7;
    11'b00100110000: data <= 32'h3e6ebc4a;
    11'b00100110001: data <= 32'h3e363bab;
    11'b00100110010: data <= 32'h3b343df9;
    11'b00100110011: data <= 32'h3a0331db;
    11'b00100110100: data <= 32'h3abfbba7;
    11'b00100110101: data <= 32'haab6ba26;
    11'b00100110110: data <= 32'hbea7b60e;
    11'b00100110111: data <= 32'hbffebb88;
    11'b00100111000: data <= 32'hb4a0bec7;
    11'b00100111001: data <= 32'h3dc2bd70;
    11'b00100111010: data <= 32'h3c00b41d;
    11'b00100111011: data <= 32'hbb133686;
    11'b00100111100: data <= 32'hbee838c8;
    11'b00100111101: data <= 32'hbb113ca3;
    11'b00100111110: data <= 32'hb0ab3f3a;
    11'b00100111111: data <= 32'hb97e3cd9;
    11'b00101000000: data <= 32'hbd3ab874;
    11'b00101000001: data <= 32'hb85abdbc;
    11'b00101000010: data <= 32'h3bfeb130;
    11'b00101000011: data <= 32'h3ee53e9b;
    11'b00101000100: data <= 32'h3dbb3ec2;
    11'b00101000101: data <= 32'h3c7a32c3;
    11'b00101000110: data <= 32'h3b80b83c;
    11'b00101000111: data <= 32'h3026326f;
    11'b00101001000: data <= 32'hbc1a3915;
    11'b00101001001: data <= 32'hbc0bb883;
    11'b00101001010: data <= 32'h3835c058;
    11'b00101001011: data <= 32'h3ec9c08e;
    11'b00101001100: data <= 32'h3b1abc0f;
    11'b00101001101: data <= 32'hba6427e6;
    11'b00101001110: data <= 32'hbc9a350e;
    11'b00101001111: data <= 32'hb1d638aa;
    11'b00101010000: data <= 32'h9f433b7b;
    11'b00101010001: data <= 32'hbdad37be;
    11'b00101010010: data <= 32'hc110b9bc;
    11'b00101010011: data <= 32'hbe50bc63;
    11'b00101010100: data <= 32'h37e330cd;
    11'b00101010101: data <= 32'h3e0b3e20;
    11'b00101010110: data <= 32'h3c503d51;
    11'b00101010111: data <= 32'h382b33f9;
    11'b00101011000: data <= 32'h373e3503;
    11'b00101011001: data <= 32'h31d13e40;
    11'b00101011010: data <= 32'hb6ec3f2a;
    11'b00101011011: data <= 32'hb576ad38;
    11'b00101011100: data <= 32'h3a6ac062;
    11'b00101011101: data <= 32'h3e79c098;
    11'b00101011110: data <= 32'h3bfcba63;
    11'b00101011111: data <= 32'ha77a32c3;
    11'b00101100000: data <= 32'h301827f7;
    11'b00101100001: data <= 32'h3b54b35e;
    11'b00101100010: data <= 32'h355c2427;
    11'b00101100011: data <= 32'hbf10a8d6;
    11'b00101100100: data <= 32'hc205ba37;
    11'b00101100101: data <= 32'hbf2abc95;
    11'b00101100110: data <= 32'h364bb62a;
    11'b00101100111: data <= 32'h3c54383b;
    11'b00101101000: data <= 32'h31653744;
    11'b00101101001: data <= 32'hb7f22fb3;
    11'b00101101010: data <= 32'hb06a3bd0;
    11'b00101101011: data <= 32'h313440f2;
    11'b00101101100: data <= 32'hb46740cd;
    11'b00101101101: data <= 32'hb83b32f8;
    11'b00101101110: data <= 32'h31e0bf18;
    11'b00101101111: data <= 32'h3c38bdf1;
    11'b00101110000: data <= 32'h3c653065;
    11'b00101110001: data <= 32'h3af139bd;
    11'b00101110010: data <= 32'h3d53b00e;
    11'b00101110011: data <= 32'h3f2db99f;
    11'b00101110100: data <= 32'h39b9b279;
    11'b00101110101: data <= 32'hbe0d3208;
    11'b00101110110: data <= 32'hc0feb803;
    11'b00101110111: data <= 32'hbc7cbda7;
    11'b00101111000: data <= 32'h399fbd89;
    11'b00101111001: data <= 32'h399bba32;
    11'b00101111010: data <= 32'hb914b7fa;
    11'b00101111011: data <= 32'hbc6eb246;
    11'b00101111100: data <= 32'hb3a33c08;
    11'b00101111101: data <= 32'h344540c7;
    11'b00101111110: data <= 32'hb8814041;
    11'b00101111111: data <= 32'hbddd3158;
    11'b00110000000: data <= 32'hbc23bcd6;
    11'b00110000001: data <= 32'h32dcb734;
    11'b00110000010: data <= 32'h3be03c24;
    11'b00110000011: data <= 32'h3cfe3c20;
    11'b00110000100: data <= 32'h3ed2b2c4;
    11'b00110000101: data <= 32'h3fc5b8a2;
    11'b00110000110: data <= 32'h3b5137e8;
    11'b00110000111: data <= 32'hbae33cb3;
    11'b00110001000: data <= 32'hbda22f45;
    11'b00110001001: data <= 32'haffbbe4b;
    11'b00110001010: data <= 32'h3c54c03f;
    11'b00110001011: data <= 32'h380bbe32;
    11'b00110001100: data <= 32'hba99bbd6;
    11'b00110001101: data <= 32'hba6ab861;
    11'b00110001110: data <= 32'h36b93668;
    11'b00110001111: data <= 32'h39193dc2;
    11'b00110010000: data <= 32'hbbb53cfe;
    11'b00110010001: data <= 32'hc0faaf42;
    11'b00110010010: data <= 32'hc02fba86;
    11'b00110010011: data <= 32'hb7132f03;
    11'b00110010100: data <= 32'h392b3cb9;
    11'b00110010101: data <= 32'h3ab939dc;
    11'b00110010110: data <= 32'h3c36b63a;
    11'b00110010111: data <= 32'h3d61acbf;
    11'b00110011000: data <= 32'h3ae23e8e;
    11'b00110011001: data <= 32'hb36340b7;
    11'b00110011010: data <= 32'hb8253a49;
    11'b00110011011: data <= 32'h369cbdaa;
    11'b00110011100: data <= 32'h3c58c020;
    11'b00110011101: data <= 32'h36c8bd33;
    11'b00110011110: data <= 32'hb63ab9dc;
    11'b00110011111: data <= 32'h33fcba07;
    11'b00110100000: data <= 32'h3e2fb706;
    11'b00110100001: data <= 32'h3ccb353b;
    11'b00110100010: data <= 32'hbc57378e;
    11'b00110100011: data <= 32'hc1bbb472;
    11'b00110100100: data <= 32'hc097b99d;
    11'b00110100101: data <= 32'hb837ae75;
    11'b00110100110: data <= 32'h341b36b0;
    11'b00110100111: data <= 32'hae08b140;
    11'b00110101000: data <= 32'hb031ba0d;
    11'b00110101001: data <= 32'h381d3547;
    11'b00110101010: data <= 32'h39c040da;
    11'b00110101011: data <= 32'h2b5941f5;
    11'b00110101100: data <= 32'hb6513c7f;
    11'b00110101101: data <= 32'h29e4bbec;
    11'b00110101110: data <= 32'h3823bcdf;
    11'b00110101111: data <= 32'h3476b32a;
    11'b00110110000: data <= 32'h3311a17a;
    11'b00110110001: data <= 32'h3d41ba42;
    11'b00110110010: data <= 32'h40eabc0e;
    11'b00110110011: data <= 32'h3eafb1e9;
    11'b00110110100: data <= 32'hba3636f7;
    11'b00110110101: data <= 32'hc09ca578;
    11'b00110110110: data <= 32'hbe0bb9d5;
    11'b00110110111: data <= 32'ha86fba59;
    11'b00110111000: data <= 32'h96d3b9d7;
    11'b00110111001: data <= 32'hbbd4bcab;
    11'b00110111010: data <= 32'hbc11bcdc;
    11'b00110111011: data <= 32'h30873415;
    11'b00110111100: data <= 32'h3a364093;
    11'b00110111101: data <= 32'h9f97413f;
    11'b00110111110: data <= 32'hbc0f3b73;
    11'b00110111111: data <= 32'hbbfdb83f;
    11'b00111000000: data <= 32'hb61faf63;
    11'b00111000001: data <= 32'ha56c3b71;
    11'b00111000010: data <= 32'h373538a3;
    11'b00111000011: data <= 32'h3e7eba57;
    11'b00111000100: data <= 32'h411dbc5c;
    11'b00111000101: data <= 32'h3f1c3226;
    11'b00111000110: data <= 32'hb2823cea;
    11'b00111000111: data <= 32'hbca23934;
    11'b00111001000: data <= 32'hb473b962;
    11'b00111001001: data <= 32'h38f3bd5b;
    11'b00111001010: data <= 32'hae72bdb7;
    11'b00111001011: data <= 32'hbd60be8b;
    11'b00111001100: data <= 32'hbc1dbe20;
    11'b00111001101: data <= 32'h38b4b4ed;
    11'b00111001110: data <= 32'h3cc33d21;
    11'b00111001111: data <= 32'hb1933e20;
    11'b00111010000: data <= 32'hbf3f362f;
    11'b00111010001: data <= 32'hbfe0b3f7;
    11'b00111010010: data <= 32'hbc3e38ca;
    11'b00111010011: data <= 32'hb6253d91;
    11'b00111010100: data <= 32'h29bc381c;
    11'b00111010101: data <= 32'h3b57bbf3;
    11'b00111010110: data <= 32'h3f1cba93;
    11'b00111010111: data <= 32'h3dec3c58;
    11'b00111011000: data <= 32'h34f1409f;
    11'b00111011001: data <= 32'hb03c3d7c;
    11'b00111011010: data <= 32'h3896b6f3;
    11'b00111011011: data <= 32'h3b06bcf3;
    11'b00111011100: data <= 32'hb1c4bc83;
    11'b00111011101: data <= 32'hbc91bcfb;
    11'b00111011110: data <= 32'hb3edbe1e;
    11'b00111011111: data <= 32'h3e64bc22;
    11'b00111100000: data <= 32'h3f452a72;
    11'b00111100001: data <= 32'hb15a3724;
    11'b00111100010: data <= 32'hc035aac2;
    11'b00111100011: data <= 32'hc03db14d;
    11'b00111100100: data <= 32'hbc2d38e7;
    11'b00111100101: data <= 32'hb8e83b53;
    11'b00111100110: data <= 32'hba58b3f7;
    11'b00111100111: data <= 32'hb5f5bdbd;
    11'b00111101000: data <= 32'h3934b8ad;
    11'b00111101001: data <= 32'h3c343f03;
    11'b00111101010: data <= 32'h384f41c3;
    11'b00111101011: data <= 32'h32863e9a;
    11'b00111101100: data <= 32'h3814af4d;
    11'b00111101101: data <= 32'h377cb76c;
    11'b00111101110: data <= 32'hb65b2963;
    11'b00111101111: data <= 32'hb9cfb3f3;
    11'b00111110000: data <= 32'h3951bd14;
    11'b00111110001: data <= 32'h40eabe1c;
    11'b00111110010: data <= 32'h408cb947;
    11'b00111110011: data <= 32'h2de42dce;
    11'b00111110100: data <= 32'hbe572328;
    11'b00111110101: data <= 32'hbd01b049;
    11'b00111110110: data <= 32'hb4e0304a;
    11'b00111110111: data <= 32'hb8c3aa9f;
    11'b00111111000: data <= 32'hbe56bccc;
    11'b00111111001: data <= 32'hbdc4bfaa;
    11'b00111111010: data <= 32'haa9cb94f;
    11'b00111111011: data <= 32'h3b173e7d;
    11'b00111111100: data <= 32'h381540e7;
    11'b00111111101: data <= 32'hb2283cfc;
    11'b00111111110: data <= 32'hb5322e01;
    11'b00111111111: data <= 32'hb5ed385a;
    11'b01000000000: data <= 32'hba013d79;
    11'b01000000001: data <= 32'hb86c396b;
    11'b01000000010: data <= 32'h3b9fbc1d;
    11'b01000000011: data <= 32'h40ffbe74;
    11'b01000000100: data <= 32'h406cb814;
    11'b01000000101: data <= 32'h372f392b;
    11'b01000000110: data <= 32'hb83238d8;
    11'b01000000111: data <= 32'h30989d41;
    11'b01000001000: data <= 32'h3978b4f6;
    11'b01000001001: data <= 32'hb6bdb99a;
    11'b01000001010: data <= 32'hbfbcbe7f;
    11'b01000001011: data <= 32'hbeb8c039;
    11'b01000001100: data <= 32'h3022bc38;
    11'b01000001101: data <= 32'h3cc5398b;
    11'b01000001110: data <= 32'h36c03cd6;
    11'b01000001111: data <= 32'hbacf35fe;
    11'b01000010000: data <= 32'hbcdc2dcf;
    11'b01000010001: data <= 32'hbc123ce3;
    11'b01000010010: data <= 32'hbc2e401c;
    11'b01000010011: data <= 32'hbab23b39;
    11'b01000010100: data <= 32'h34edbc5c;
    11'b01000010101: data <= 32'h3e58bdac;
    11'b01000010110: data <= 32'h3e6c32ff;
    11'b01000010111: data <= 32'h39653e7a;
    11'b01000011000: data <= 32'h37393d34;
    11'b01000011001: data <= 32'h3ce032c9;
    11'b01000011010: data <= 32'h3d0ab46f;
    11'b01000011011: data <= 32'hb53cb712;
    11'b01000011100: data <= 32'hbf2abc7e;
    11'b01000011101: data <= 32'hbc56bf56;
    11'b01000011110: data <= 32'h3c00be05;
    11'b01000011111: data <= 32'h3f2bb7b1;
    11'b01000100000: data <= 32'h371eae46;
    11'b01000100001: data <= 32'hbca5b67a;
    11'b01000100010: data <= 32'hbd8da851;
    11'b01000100011: data <= 32'hbb523d1f;
    11'b01000100100: data <= 32'hbc2a3f1f;
    11'b01000100101: data <= 32'hbdb134fa;
    11'b01000100110: data <= 32'hbb5cbdf8;
    11'b01000100111: data <= 32'h33c9bce4;
    11'b01000101000: data <= 32'h3a913ae3;
    11'b01000101001: data <= 32'h39524061;
    11'b01000101010: data <= 32'h3a843e13;
    11'b01000101011: data <= 32'h3d7f3594;
    11'b01000101100: data <= 32'h3c39347c;
    11'b01000101101: data <= 32'hb7c9395a;
    11'b01000101110: data <= 32'hbdbd2cf7;
    11'b01000101111: data <= 32'hb37abcdc;
    11'b01000110000: data <= 32'h3f5ebef2;
    11'b01000110001: data <= 32'h406bbccd;
    11'b01000110010: data <= 32'h3891b980;
    11'b01000110011: data <= 32'hba8bb8ab;
    11'b01000110100: data <= 32'hb895ada6;
    11'b01000110101: data <= 32'h20f43af5;
    11'b01000110110: data <= 32'hb9673b45;
    11'b01000110111: data <= 32'hbfc2b8cd;
    11'b01000111000: data <= 32'hbff1bfcf;
    11'b01000111001: data <= 32'hb9a3bcde;
    11'b01000111010: data <= 32'h35ec3ae8;
    11'b01000111011: data <= 32'h381e3f3a;
    11'b01000111100: data <= 32'h37c73b9f;
    11'b01000111101: data <= 32'h39573374;
    11'b01000111110: data <= 32'h348a3c11;
    11'b01000111111: data <= 32'hbaa23fed;
    11'b01001000000: data <= 32'hbce13d06;
    11'b01001000001: data <= 32'h30c1b93a;
    11'b01001000010: data <= 32'h3fb3bea5;
    11'b01001000011: data <= 32'h4007bc73;
    11'b01001000100: data <= 32'h391ab4a4;
    11'b01001000101: data <= 32'ha418adee;
    11'b01001000110: data <= 32'h3a6e277a;
    11'b01001000111: data <= 32'h3d0336b8;
    11'b01001001000: data <= 32'hb0fb3290;
    11'b01001001001: data <= 32'hc030bc40;
    11'b01001001010: data <= 32'hc08dc019;
    11'b01001001011: data <= 32'hb9afbd70;
    11'b01001001100: data <= 32'h38483188;
    11'b01001001101: data <= 32'h366c38b1;
    11'b01001001110: data <= 32'hb0d1b17a;
    11'b01001001111: data <= 32'hb3a9b031;
    11'b01001010000: data <= 32'hb64c3de7;
    11'b01001010001: data <= 32'hbc3b416c;
    11'b01001010010: data <= 32'hbd353ec8;
    11'b01001010011: data <= 32'hb485b83b;
    11'b01001010100: data <= 32'h3c27bdab;
    11'b01001010101: data <= 32'h3cacb6c2;
    11'b01001010110: data <= 32'h37fc394d;
    11'b01001010111: data <= 32'h39cb38f2;
    11'b01001011000: data <= 32'h3fad32b5;
    11'b01001011001: data <= 32'h402334ce;
    11'b01001011010: data <= 32'h316d3473;
    11'b01001011011: data <= 32'hbf7fb8c5;
    11'b01001011100: data <= 32'hbee9be38;
    11'b01001011101: data <= 32'h2eaebdd1;
    11'b01001011110: data <= 32'h3c83ba0c;
    11'b01001011111: data <= 32'h367fba0f;
    11'b01001100000: data <= 32'hb88cbcdb;
    11'b01001100001: data <= 32'hb888b83d;
    11'b01001100010: data <= 32'hb5583db2;
    11'b01001100011: data <= 32'hbaf840fc;
    11'b01001100100: data <= 32'hbe393cc8;
    11'b01001100101: data <= 32'hbd0fbb2a;
    11'b01001100110: data <= 32'hb55ebcd8;
    11'b01001100111: data <= 32'h2e9734a1;
    11'b01001101000: data <= 32'h31a53d6d;
    11'b01001101001: data <= 32'h3b943b15;
    11'b01001101010: data <= 32'h4045326c;
    11'b01001101011: data <= 32'h3ffc387c;
    11'b01001101100: data <= 32'h2d543c9a;
    11'b01001101101: data <= 32'hbe043904;
    11'b01001101110: data <= 32'hbab3b931;
    11'b01001101111: data <= 32'h3c28bd5f;
    11'b01001110000: data <= 32'h3e62bd3c;
    11'b01001110001: data <= 32'h36c5bda8;
    11'b01001110010: data <= 32'hb7b8be43;
    11'b01001110011: data <= 32'h25f9b99e;
    11'b01001110100: data <= 32'h38d13be5;
    11'b01001110101: data <= 32'hb33f3e6c;
    11'b01001110110: data <= 32'hbedd331e;
    11'b01001110111: data <= 32'hc048bd9e;
    11'b01001111000: data <= 32'hbd6cbc83;
    11'b01001111001: data <= 32'hb87f3813;
    11'b01001111010: data <= 32'hb08b3cbb;
    11'b01001111011: data <= 32'h38973524;
    11'b01001111100: data <= 32'h3dbfb19b;
    11'b01001111101: data <= 32'h3cca3b83;
    11'b01001111110: data <= 32'hb4c94085;
    11'b01001111111: data <= 32'hbcf43f85;
    11'b01010000000: data <= 32'hb4683137;
    11'b01010000001: data <= 32'h3d42bc33;
    11'b01010000010: data <= 32'h3dadbc9a;
    11'b01010000011: data <= 32'h341dbc2f;
    11'b01010000100: data <= 32'ha6bcbc5c;
    11'b01010000101: data <= 32'h3cc3b886;
    11'b01010000110: data <= 32'h3fae380c;
    11'b01010000111: data <= 32'h38923a10;
    11'b01010001000: data <= 32'hbe6eb6b1;
    11'b01010001001: data <= 32'hc0acbe26;
    11'b01010001010: data <= 32'hbda3bc48;
    11'b01010001011: data <= 32'hb75f30a5;
    11'b01010001100: data <= 32'hb44f3185;
    11'b01010001101: data <= 32'had7dbafb;
    11'b01010001110: data <= 32'h36b4baab;
    11'b01010001111: data <= 32'h35c83c66;
    11'b01010010000: data <= 32'hb8a641bf;
    11'b01010010001: data <= 32'hbca140c5;
    11'b01010010010: data <= 32'hb67a366b;
    11'b01010010011: data <= 32'h391fb9fc;
    11'b01010010100: data <= 32'h381bb6f7;
    11'b01010010101: data <= 32'hb1d2a330;
    11'b01010010110: data <= 32'h3648b3e0;
    11'b01010010111: data <= 32'h4058b524;
    11'b01010011000: data <= 32'h41a3342b;
    11'b01010011001: data <= 32'h3c3c3876;
    11'b01010011010: data <= 32'hbd20b143;
    11'b01010011011: data <= 32'hbf02bc00;
    11'b01010011100: data <= 32'hb85abafa;
    11'b01010011101: data <= 32'h336db72e;
    11'b01010011110: data <= 32'hb276bc19;
    11'b01010011111: data <= 32'hb8c7c007;
    11'b01010100000: data <= 32'hb0d2bdc4;
    11'b01010100001: data <= 32'h32a83b2b;
    11'b01010100010: data <= 32'hb6064135;
    11'b01010100011: data <= 32'hbc8c3f72;
    11'b01010100100: data <= 32'hbc31a68d;
    11'b01010100101: data <= 32'hb89ab8bb;
    11'b01010100110: data <= 32'hb94a3590;
    11'b01010100111: data <= 32'hba0a3b22;
    11'b01010101000: data <= 32'h36b0335c;
    11'b01010101001: data <= 32'h40a7b523;
    11'b01010101010: data <= 32'h41813468;
    11'b01010101011: data <= 32'h3bac3c63;
    11'b01010101100: data <= 32'hbb7d3b1d;
    11'b01010101101: data <= 32'hba6e241e;
    11'b01010101110: data <= 32'h3897b7a9;
    11'b01010101111: data <= 32'h3b34ba1c;
    11'b01010110000: data <= 32'hb0dcbe6f;
    11'b01010110001: data <= 32'hb9c9c0cf;
    11'b01010110010: data <= 32'h2f90be9c;
    11'b01010110011: data <= 32'h3bb4373a;
    11'b01010110100: data <= 32'h35ed3eaa;
    11'b01010110101: data <= 32'hbbfa39de;
    11'b01010110110: data <= 32'hbe9eb9c4;
    11'b01010110111: data <= 32'hbe0cb878;
    11'b01010111000: data <= 32'hbd9939fa;
    11'b01010111001: data <= 32'hbcad3c17;
    11'b01010111010: data <= 32'h957db089;
    11'b01010111011: data <= 32'h3e51ba40;
    11'b01010111100: data <= 32'h3f5135a1;
    11'b01010111101: data <= 32'h36973fa7;
    11'b01010111110: data <= 32'hb9d74018;
    11'b01010111111: data <= 32'hadc33b6f;
    11'b01011000000: data <= 32'h3c8da822;
    11'b01011000001: data <= 32'h3b69b820;
    11'b01011000010: data <= 32'hb60fbcc6;
    11'b01011000011: data <= 32'hb87abf5e;
    11'b01011000100: data <= 32'h3bd7bd89;
    11'b01011000101: data <= 32'h40592799;
    11'b01011000110: data <= 32'h3d283985;
    11'b01011000111: data <= 32'hb97db1ba;
    11'b01011001000: data <= 32'hbedcbc45;
    11'b01011001001: data <= 32'hbe12b77c;
    11'b01011001010: data <= 32'hbd023945;
    11'b01011001011: data <= 32'hbcd6352c;
    11'b01011001100: data <= 32'hb8e9bcdf;
    11'b01011001101: data <= 32'h3742be49;
    11'b01011001110: data <= 32'h39ec3456;
    11'b01011001111: data <= 32'hade140b4;
    11'b01011010000: data <= 32'hb9274101;
    11'b01011010001: data <= 32'h28863ca8;
    11'b01011010010: data <= 32'h3a39338b;
    11'b01011010011: data <= 32'h30e9319c;
    11'b01011010100: data <= 32'hbb99ac72;
    11'b01011010101: data <= 32'hb68eba2a;
    11'b01011010110: data <= 32'h3f06bb58;
    11'b01011010111: data <= 32'h420bb23f;
    11'b01011011000: data <= 32'h3f423421;
    11'b01011011001: data <= 32'hb55eb3ba;
    11'b01011011010: data <= 32'hbc7eb976;
    11'b01011011011: data <= 32'hb894b0aa;
    11'b01011011100: data <= 32'hb5ce3599;
    11'b01011011101: data <= 32'hbb76b926;
    11'b01011011110: data <= 32'hbc58c09d;
    11'b01011011111: data <= 32'hb52bc083;
    11'b01011100000: data <= 32'h3455a378;
    11'b01011100001: data <= 32'hac0e4014;
    11'b01011100010: data <= 32'hb82a3fa3;
    11'b01011100011: data <= 32'hb51238a0;
    11'b01011100100: data <= 32'hb1fd32b3;
    11'b01011100101: data <= 32'hbbbb3b4d;
    11'b01011100110: data <= 32'hbe883c15;
    11'b01011100111: data <= 32'hb8252466;
    11'b01011101000: data <= 32'h3f56b9bf;
    11'b01011101001: data <= 32'h41cbb419;
    11'b01011101010: data <= 32'h3e643812;
    11'b01011101011: data <= 32'hb05f3856;
    11'b01011101100: data <= 32'hb2eb344e;
    11'b01011101101: data <= 32'h39b1361b;
    11'b01011101110: data <= 32'h38dc32e7;
    11'b01011101111: data <= 32'hb952bc7c;
    11'b01011110000: data <= 32'hbd08c14e;
    11'b01011110001: data <= 32'hb550c0cc;
    11'b01011110010: data <= 32'h39e8b5b8;
    11'b01011110011: data <= 32'h38ce3c87;
    11'b01011110100: data <= 32'hb386390c;
    11'b01011110101: data <= 32'hb9a0b676;
    11'b01011110110: data <= 32'hbbe723ac;
    11'b01011110111: data <= 32'hbeb03d54;
    11'b01011111000: data <= 32'hc00f3da9;
    11'b01011111001: data <= 32'hbb1aaad1;
    11'b01011111010: data <= 32'h3c65bc48;
    11'b01011111011: data <= 32'h3f5cb528;
    11'b01011111100: data <= 32'h3a4a3c50;
    11'b01011111101: data <= 32'hb1043e26;
    11'b01011111110: data <= 32'h37fc3ca3;
    11'b01011111111: data <= 32'h3e1b3ae5;
    11'b01100000000: data <= 32'h3b933784;
    11'b01100000001: data <= 32'hba0eb994;
    11'b01100000010: data <= 32'hbce5bfe9;
    11'b01100000011: data <= 32'h3446bf96;
    11'b01100000100: data <= 32'h3f0cb885;
    11'b01100000101: data <= 32'h3dff314f;
    11'b01100000110: data <= 32'h30eab82d;
    11'b01100000111: data <= 32'hb99fbc4d;
    11'b01100001000: data <= 32'hbbb3ab53;
    11'b01100001001: data <= 32'hbdbf3d6a;
    11'b01100001010: data <= 32'hbf863be7;
    11'b01100001011: data <= 32'hbd3dbb57;
    11'b01100001100: data <= 32'ha15bbf58;
    11'b01100001101: data <= 32'h382fb81a;
    11'b01100001110: data <= 32'haa513da1;
    11'b01100001111: data <= 32'hb42b3fbf;
    11'b01100010000: data <= 32'h39b53d53;
    11'b01100010001: data <= 32'h3dc53bf2;
    11'b01100010010: data <= 32'h368e3c07;
    11'b01100010011: data <= 32'hbd293695;
    11'b01100010100: data <= 32'hbcd0b98d;
    11'b01100010101: data <= 32'h3b24bc66;
    11'b01100010110: data <= 32'h4110b8a0;
    11'b01100010111: data <= 32'h3ff1b555;
    11'b01100011000: data <= 32'h36c4baeb;
    11'b01100011001: data <= 32'hb303bb9e;
    11'b01100011010: data <= 32'ha68f32a1;
    11'b01100011011: data <= 32'hb5b73cbd;
    11'b01100011100: data <= 32'hbd263281;
    11'b01100011101: data <= 32'hbe3cbfa3;
    11'b01100011110: data <= 32'hbaaec100;
    11'b01100011111: data <= 32'hb34fba29;
    11'b01100100000: data <= 32'hb4fb3c9f;
    11'b01100100001: data <= 32'hb31f3d5e;
    11'b01100100010: data <= 32'h380238a5;
    11'b01100100011: data <= 32'h39803969;
    11'b01100100100: data <= 32'hb8bc3e17;
    11'b01100100101: data <= 32'hbfe03e23;
    11'b01100100110: data <= 32'hbd5435fd;
    11'b01100100111: data <= 32'h3bdeb8aa;
    11'b01100101000: data <= 32'h40c9b829;
    11'b01100101001: data <= 32'h3e87b2e4;
    11'b01100101010: data <= 32'h35e8b507;
    11'b01100101011: data <= 32'h37b3b09c;
    11'b01100101100: data <= 32'h3d2139e5;
    11'b01100101101: data <= 32'h3b1b3c73;
    11'b01100101110: data <= 32'hb977b3c6;
    11'b01100101111: data <= 32'hbe51c077;
    11'b01100110000: data <= 32'hbbb4c113;
    11'b01100110001: data <= 32'ha35bbb40;
    11'b01100110010: data <= 32'h31b036d6;
    11'b01100110011: data <= 32'h2bc52977;
    11'b01100110100: data <= 32'h32b4b957;
    11'b01100110101: data <= 32'ha956305d;
    11'b01100110110: data <= 32'hbd133f0e;
    11'b01100110111: data <= 32'hc0984011;
    11'b01100111000: data <= 32'hbe303899;
    11'b01100111001: data <= 32'h365db9cd;
    11'b01100111010: data <= 32'h3d45b889;
    11'b01100111011: data <= 32'h388e33a3;
    11'b01100111100: data <= 32'h1d2b3892;
    11'b01100111101: data <= 32'h3c0239a5;
    11'b01100111110: data <= 32'h40603cba;
    11'b01100111111: data <= 32'h3e0d3d10;
    11'b01101000000: data <= 32'hb8382c39;
    11'b01101000001: data <= 32'hbdffbe2b;
    11'b01101000010: data <= 32'hb7d6bf3c;
    11'b01101000011: data <= 32'h3aecba43;
    11'b01101000100: data <= 32'h3c12b565;
    11'b01101000101: data <= 32'h370abcc5;
    11'b01101000110: data <= 32'h313bbe8c;
    11'b01101000111: data <= 32'hadfdb2f7;
    11'b01101001000: data <= 32'hbc153ed8;
    11'b01101001001: data <= 32'hbfcf3eef;
    11'b01101001010: data <= 32'hbea8af64;
    11'b01101001011: data <= 32'hb81abda1;
    11'b01101001100: data <= 32'haccbba1a;
    11'b01101001101: data <= 32'hb8983889;
    11'b01101001110: data <= 32'hb6963c0a;
    11'b01101001111: data <= 32'h3c733af5;
    11'b01101010000: data <= 32'h40773ca1;
    11'b01101010001: data <= 32'h3cb73e26;
    11'b01101010010: data <= 32'hbb993be3;
    11'b01101010011: data <= 32'hbdf3b216;
    11'b01101010100: data <= 32'h2e54b99d;
    11'b01101010101: data <= 32'h3e8db758;
    11'b01101010110: data <= 32'h3dfeb9a6;
    11'b01101010111: data <= 32'h38c5bea7;
    11'b01101011000: data <= 32'h36dabefe;
    11'b01101011001: data <= 32'h3963ae70;
    11'b01101011010: data <= 32'h2f7a3e2b;
    11'b01101011011: data <= 32'hbc3a3c0e;
    11'b01101011100: data <= 32'hbe40bc4e;
    11'b01101011101: data <= 32'hbcbdc021;
    11'b01101011110: data <= 32'hbba2bb91;
    11'b01101011111: data <= 32'hbc6937ba;
    11'b01101100000: data <= 32'hb87e387c;
    11'b01101100001: data <= 32'h3b182c99;
    11'b01101100010: data <= 32'h3e41387b;
    11'b01101100011: data <= 32'h33b63ed1;
    11'b01101100100: data <= 32'hbe743fc5;
    11'b01101100101: data <= 32'hbe4c3c04;
    11'b01101100110: data <= 32'h34f42f1c;
    11'b01101100111: data <= 32'h3e7ab167;
    11'b01101101000: data <= 32'h3c71b86c;
    11'b01101101001: data <= 32'h34adbcde;
    11'b01101101010: data <= 32'h3a60bc27;
    11'b01101101011: data <= 32'h3f3c366b;
    11'b01101101100: data <= 32'h3def3dd1;
    11'b01101101101: data <= 32'hb04f37db;
    11'b01101101110: data <= 32'hbd3cbdfc;
    11'b01101101111: data <= 32'hbd02c02a;
    11'b01101110000: data <= 32'hbae0baf3;
    11'b01101110001: data <= 32'hba052b85;
    11'b01101110010: data <= 32'hb54bb88d;
    11'b01101110011: data <= 32'h38c0bd2b;
    11'b01101110100: data <= 32'h3a62b4f7;
    11'b01101110101: data <= 32'hb80e3e8e;
    11'b01101110110: data <= 32'hbfbf40b5;
    11'b01101110111: data <= 32'hbe783d57;
    11'b01101111000: data <= 32'h9eff30d2;
    11'b01101111001: data <= 32'h39a5b018;
    11'b01101111010: data <= 32'habc1ae97;
    11'b01101111011: data <= 32'hb676b54a;
    11'b01101111100: data <= 32'h3becb09b;
    11'b01101111101: data <= 32'h41383ad3;
    11'b01101111110: data <= 32'h40803dea;
    11'b01101111111: data <= 32'h33d9388d;
    11'b01110000000: data <= 32'hbc65bba9;
    11'b01110000001: data <= 32'hba35bd08;
    11'b01110000010: data <= 32'ha0dfb6c4;
    11'b01110000011: data <= 32'h2e77b5eb;
    11'b01110000100: data <= 32'h2bc5bebf;
    11'b01110000101: data <= 32'h375cc0d3;
    11'b01110000110: data <= 32'h3871bb6d;
    11'b01110000111: data <= 32'hb6763da4;
    11'b01110001000: data <= 32'hbe124014;
    11'b01110001001: data <= 32'hbdbb399d;
    11'b01110001010: data <= 32'hb8aab810;
    11'b01110001011: data <= 32'hb87eb545;
    11'b01110001100: data <= 32'hbd74347e;
    11'b01110001101: data <= 32'hbc7a3420;
    11'b01110001110: data <= 32'h3b1230ed;
    11'b01110001111: data <= 32'h413e3a3f;
    11'b01110010000: data <= 32'h3ffd3dec;
    11'b01110010001: data <= 32'haf203cab;
    11'b01110010010: data <= 32'hbc4c3435;
    11'b01110010011: data <= 32'hb0ee21cb;
    11'b01110010100: data <= 32'h3aff334b;
    11'b01110010101: data <= 32'h399bb7c1;
    11'b01110010110: data <= 32'h3236c039;
    11'b01110010111: data <= 32'h37f3c143;
    11'b01110011000: data <= 32'h3c16bb61;
    11'b01110011001: data <= 32'h38c83ccf;
    11'b01110011010: data <= 32'hb7753d30;
    11'b01110011011: data <= 32'hbbe8b562;
    11'b01110011100: data <= 32'hbbc5bd11;
    11'b01110011101: data <= 32'hbd89b815;
    11'b01110011110: data <= 32'hc00d361c;
    11'b01110011111: data <= 32'hbdb92d36;
    11'b01110100000: data <= 32'h38a9b808;
    11'b01110100001: data <= 32'h3fbe2981;
    11'b01110100010: data <= 32'h3c0e3d37;
    11'b01110100011: data <= 32'hbad63f46;
    11'b01110100100: data <= 32'hbcb03d8f;
    11'b01110100101: data <= 32'h32803bde;
    11'b01110100110: data <= 32'h3c6539d9;
    11'b01110100111: data <= 32'h3747b2ed;
    11'b01110101000: data <= 32'hb345be99;
    11'b01110101001: data <= 32'h3847bfa3;
    11'b01110101010: data <= 32'h3f5fb5ee;
    11'b01110101011: data <= 32'h3f8d3c83;
    11'b01110101100: data <= 32'h39143949;
    11'b01110101101: data <= 32'hb794bbc3;
    11'b01110101110: data <= 32'hbb0cbdb6;
    11'b01110101111: data <= 32'hbd16b57d;
    11'b01110110000: data <= 32'hbece343b;
    11'b01110110001: data <= 32'hbcc1b9e5;
    11'b01110110010: data <= 32'h34cdbf21;
    11'b01110110011: data <= 32'h3c55bc10;
    11'b01110110100: data <= 32'h2d173b84;
    11'b01110110101: data <= 32'hbd494011;
    11'b01110110110: data <= 32'hbc9d3ecc;
    11'b01110110111: data <= 32'h31393c5b;
    11'b01110111000: data <= 32'h37ce3a79;
    11'b01110111001: data <= 32'hb8fa33b6;
    11'b01110111010: data <= 32'hbc74b995;
    11'b01110111011: data <= 32'h3674badd;
    11'b01110111100: data <= 32'h40d43327;
    11'b01110111101: data <= 32'h41423c7b;
    11'b01110111110: data <= 32'h3c7937eb;
    11'b01110111111: data <= 32'hb176b9c8;
    11'b01111000000: data <= 32'hb5ebb9a8;
    11'b01111000001: data <= 32'hb5f7348f;
    11'b01111000010: data <= 32'hb9cc3189;
    11'b01111000011: data <= 32'hb954be68;
    11'b01111000100: data <= 32'h3105c1c0;
    11'b01111000101: data <= 32'h390dbf19;
    11'b01111000110: data <= 32'hae26387f;
    11'b01111000111: data <= 32'hbc153e97;
    11'b01111001000: data <= 32'hba6f3c1d;
    11'b01111001001: data <= 32'haccd3586;
    11'b01111001010: data <= 32'hb81937fe;
    11'b01111001011: data <= 32'hbf9538f4;
    11'b01111001100: data <= 32'hc0002c47;
    11'b01111001101: data <= 32'h2e2ab4bc;
    11'b01111001110: data <= 32'h40a53492;
    11'b01111001111: data <= 32'h40b13be1;
    11'b01111010000: data <= 32'h39c03a1c;
    11'b01111010001: data <= 32'hb3043309;
    11'b01111010010: data <= 32'h33d0383b;
    11'b01111010011: data <= 32'h39443c86;
    11'b01111010100: data <= 32'h2fbb34dc;
    11'b01111010101: data <= 32'hb624bf8f;
    11'b01111010110: data <= 32'h2dadc225;
    11'b01111010111: data <= 32'h3a4bbf14;
    11'b01111011000: data <= 32'h38f73621;
    11'b01111011001: data <= 32'ha2953b3d;
    11'b01111011010: data <= 32'hb0cfb046;
    11'b01111011011: data <= 32'hb1c5b917;
    11'b01111011100: data <= 32'hbcad3132;
    11'b01111011101: data <= 32'hc1193a58;
    11'b01111011110: data <= 32'hc0b831a8;
    11'b01111011111: data <= 32'hb332b954;
    11'b01111100000: data <= 32'h3e78b645;
    11'b01111100001: data <= 32'h3d0938c7;
    11'b01111100010: data <= 32'hb30c3c6d;
    11'b01111100011: data <= 32'hb78c3ca0;
    11'b01111100100: data <= 32'h392f3e03;
    11'b01111100101: data <= 32'h3c923eee;
    11'b01111100110: data <= 32'h3138392b;
    11'b01111100111: data <= 32'hb9c8bd8e;
    11'b01111101000: data <= 32'hac85c089;
    11'b01111101001: data <= 32'h3d25bc37;
    11'b01111101010: data <= 32'h3ecc373f;
    11'b01111101011: data <= 32'h3c6233aa;
    11'b01111101100: data <= 32'h3811bc03;
    11'b01111101101: data <= 32'h2911bc55;
    11'b01111101110: data <= 32'hbbf43331;
    11'b01111101111: data <= 32'hc0533ace;
    11'b01111110000: data <= 32'hbffcb515;
    11'b01111110001: data <= 32'hb62fbedc;
    11'b01111110010: data <= 32'h39f7bdd5;
    11'b01111110011: data <= 32'h2f082ad3;
    11'b01111110100: data <= 32'hbbc33c8f;
    11'b01111110101: data <= 32'hb8a33d84;
    11'b01111110110: data <= 32'h3a0e3e47;
    11'b01111110111: data <= 32'h3acc3ef5;
    11'b01111111000: data <= 32'hb95d3c10;
    11'b01111111001: data <= 32'hbe6fb6bc;
    11'b01111111010: data <= 32'hb678bc17;
    11'b01111111011: data <= 32'h3e89b1eb;
    11'b01111111100: data <= 32'h40a838b8;
    11'b01111111101: data <= 32'h3e42aa22;
    11'b01111111110: data <= 32'h3a5dbc42;
    11'b01111111111: data <= 32'h3810b8f6;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    