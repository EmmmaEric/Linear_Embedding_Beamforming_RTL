
module memory_rom_49(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3deb386b;
    11'b00000000001: data <= 32'h3b1c342d;
    11'b00000000010: data <= 32'hbaa9b55c;
    11'b00000000011: data <= 32'hbd2bbd6a;
    11'b00000000100: data <= 32'h3673beb2;
    11'b00000000101: data <= 32'h405abaff;
    11'b00000000110: data <= 32'h3f75b1f3;
    11'b00000000111: data <= 32'h2e44b842;
    11'b00000001000: data <= 32'hbc08bb31;
    11'b00000001001: data <= 32'hbb91a546;
    11'b00000001010: data <= 32'hbb843cd1;
    11'b00000001011: data <= 32'hbdd83a40;
    11'b00000001100: data <= 32'hbe09bc9e;
    11'b00000001101: data <= 32'hb8d6c02e;
    11'b00000001110: data <= 32'h32c1b8dc;
    11'b00000001111: data <= 32'h305a3e58;
    11'b00000010000: data <= 32'ha7314042;
    11'b00000010001: data <= 32'h38983cb4;
    11'b00000010010: data <= 32'h3c3e38ef;
    11'b00000010011: data <= 32'h30d23bcf;
    11'b00000010100: data <= 32'hbd543b9d;
    11'b00000010101: data <= 32'hbca3ae46;
    11'b00000010110: data <= 32'h3bd5bc36;
    11'b00000010111: data <= 32'h415abba5;
    11'b00000011000: data <= 32'h401eb7ae;
    11'b00000011001: data <= 32'h34eab812;
    11'b00000011010: data <= 32'hb4f9b82f;
    11'b00000011011: data <= 32'h34333386;
    11'b00000011100: data <= 32'h333f3b18;
    11'b00000011101: data <= 32'hbbcea926;
    11'b00000011110: data <= 32'hbf55bfdf;
    11'b00000011111: data <= 32'hbd0dc109;
    11'b00000100000: data <= 32'hb201ba99;
    11'b00000100001: data <= 32'h30b13c60;
    11'b00000100010: data <= 32'h1d843cca;
    11'b00000100011: data <= 32'h31163403;
    11'b00000100100: data <= 32'h313f35b7;
    11'b00000100101: data <= 32'hba343e5d;
    11'b00000100110: data <= 32'hbf533ff0;
    11'b00000100111: data <= 32'hbd0b396e;
    11'b00000101000: data <= 32'h3a9bba57;
    11'b00000101001: data <= 32'h4057bb17;
    11'b00000101010: data <= 32'h3deeaecb;
    11'b00000101011: data <= 32'h349c349b;
    11'b00000101100: data <= 32'h38433504;
    11'b00000101101: data <= 32'h3e4f3910;
    11'b00000101110: data <= 32'h3d193a31;
    11'b00000101111: data <= 32'hb8acb45d;
    11'b00000110000: data <= 32'hbf55bfbb;
    11'b00000110001: data <= 32'hbc6ac0a4;
    11'b00000110010: data <= 32'h35a1bc02;
    11'b00000110011: data <= 32'h3a02313b;
    11'b00000110100: data <= 32'h3201b2e5;
    11'b00000110101: data <= 32'hb2eebb3b;
    11'b00000110110: data <= 32'hb6c6a628;
    11'b00000110111: data <= 32'hbc8e3f3d;
    11'b00000111000: data <= 32'hbfc04065;
    11'b00000111001: data <= 32'hbe253824;
    11'b00000111010: data <= 32'ha6f3bc6b;
    11'b00000111011: data <= 32'h3b0abac2;
    11'b00000111100: data <= 32'h36b637ed;
    11'b00000111101: data <= 32'h29603c8d;
    11'b00000111110: data <= 32'h3c303b71;
    11'b00000111111: data <= 32'h40783b12;
    11'b00001000000: data <= 32'h3e323c02;
    11'b00001000001: data <= 32'hb8e8359d;
    11'b00001000010: data <= 32'hbea2bb88;
    11'b00001000011: data <= 32'hb69bbe12;
    11'b00001000100: data <= 32'h3d41bbdb;
    11'b00001000101: data <= 32'h3dd5b921;
    11'b00001000110: data <= 32'h3688bd13;
    11'b00001000111: data <= 32'hb23ebe47;
    11'b00001001000: data <= 32'hb0d7b2be;
    11'b00001001001: data <= 32'hb8583e8f;
    11'b00001001010: data <= 32'hbde23e75;
    11'b00001001011: data <= 32'hbf10b5c0;
    11'b00001001100: data <= 32'hbc38befd;
    11'b00001001101: data <= 32'hb6e2bb4b;
    11'b00001001110: data <= 32'hb7d73a4e;
    11'b00001001111: data <= 32'hb3923d27;
    11'b00001010000: data <= 32'h3c1439f4;
    11'b00001010001: data <= 32'h3fc939bf;
    11'b00001010010: data <= 32'h3b993da1;
    11'b00001010011: data <= 32'hbc403dea;
    11'b00001010100: data <= 32'hbe1b3722;
    11'b00001010101: data <= 32'h323db881;
    11'b00001010110: data <= 32'h3f7eba30;
    11'b00001010111: data <= 32'h3e85bafe;
    11'b00001011000: data <= 32'h36e2bd8f;
    11'b00001011001: data <= 32'h3345bd7b;
    11'b00001011010: data <= 32'h3b3ba80b;
    11'b00001011011: data <= 32'h39f73d55;
    11'b00001011100: data <= 32'hb92d3a61;
    11'b00001011101: data <= 32'hbf17bcd3;
    11'b00001011110: data <= 32'hbe84c054;
    11'b00001011111: data <= 32'hbbdfbbe2;
    11'b00001100000: data <= 32'hb996383e;
    11'b00001100001: data <= 32'hb50e37fc;
    11'b00001100010: data <= 32'h38efb4ab;
    11'b00001100011: data <= 32'h3c58300e;
    11'b00001100100: data <= 32'h24533ec4;
    11'b00001100101: data <= 32'hbe3e40d1;
    11'b00001100110: data <= 32'hbe1a3d8b;
    11'b00001100111: data <= 32'h337ba974;
    11'b00001101000: data <= 32'h3dfeb862;
    11'b00001101001: data <= 32'h3bacb808;
    11'b00001101010: data <= 32'h2e44b945;
    11'b00001101011: data <= 32'h39ebb87a;
    11'b00001101100: data <= 32'h403635df;
    11'b00001101101: data <= 32'h3fda3ca0;
    11'b00001101110: data <= 32'h294336a1;
    11'b00001101111: data <= 32'hbe49bd28;
    11'b00001110000: data <= 32'hbdd5bf94;
    11'b00001110001: data <= 32'hb84cbb06;
    11'b00001110010: data <= 32'hb114ad25;
    11'b00001110011: data <= 32'hb092ba5d;
    11'b00001110100: data <= 32'h32a4be79;
    11'b00001110101: data <= 32'h3637b8a2;
    11'b00001110110: data <= 32'hb73e3eae;
    11'b00001110111: data <= 32'hbe7a412f;
    11'b00001111000: data <= 32'hbe373d5d;
    11'b00001111001: data <= 32'hb517b3de;
    11'b00001111010: data <= 32'h353cb798;
    11'b00001111011: data <= 32'hb4672f24;
    11'b00001111100: data <= 32'hb7de3432;
    11'b00001111101: data <= 32'h3bdb30bc;
    11'b00001111110: data <= 32'h417038c4;
    11'b00001111111: data <= 32'h40c13cb8;
    11'b00010000000: data <= 32'h31603a1a;
    11'b00010000001: data <= 32'hbd54b6bc;
    11'b00010000010: data <= 32'hba18bb70;
    11'b00010000011: data <= 32'h375db80d;
    11'b00010000100: data <= 32'h38f0b8bb;
    11'b00010000101: data <= 32'h2ccdbf2f;
    11'b00010000110: data <= 32'h2c65c0e5;
    11'b00010000111: data <= 32'h36a7bbc2;
    11'b00010001000: data <= 32'h249a3d97;
    11'b00010001001: data <= 32'hbc0a4003;
    11'b00010001010: data <= 32'hbdc03762;
    11'b00010001011: data <= 32'hbc27bb71;
    11'b00010001100: data <= 32'hbb60b862;
    11'b00010001101: data <= 32'hbd7a3832;
    11'b00010001110: data <= 32'hbc163900;
    11'b00010001111: data <= 32'h3a822daa;
    11'b00010010000: data <= 32'h40d93507;
    11'b00010010001: data <= 32'h3f3b3d0a;
    11'b00010010010: data <= 32'hb4a23e52;
    11'b00010010011: data <= 32'hbcd33b2d;
    11'b00010010100: data <= 32'hac2d3335;
    11'b00010010101: data <= 32'h3ccc9c6b;
    11'b00010010110: data <= 32'h3b53b927;
    11'b00010010111: data <= 32'h21fcbfa1;
    11'b00010011000: data <= 32'h324fc0a1;
    11'b00010011001: data <= 32'h3cabba97;
    11'b00010011010: data <= 32'h3cea3c57;
    11'b00010011011: data <= 32'h25333c7f;
    11'b00010011100: data <= 32'hbc79b845;
    11'b00010011101: data <= 32'hbd96bde2;
    11'b00010011110: data <= 32'hbddbb887;
    11'b00010011111: data <= 32'hbebb3831;
    11'b00010100000: data <= 32'hbcbc2ff5;
    11'b00010100001: data <= 32'h3623bae1;
    11'b00010100010: data <= 32'h3e12b7a6;
    11'b00010100011: data <= 32'h3a0e3ccc;
    11'b00010100100: data <= 32'hbb384088;
    11'b00010100101: data <= 32'hbcb33f4a;
    11'b00010100110: data <= 32'h32393b1c;
    11'b00010100111: data <= 32'h3c6235bf;
    11'b00010101000: data <= 32'h3579b2f9;
    11'b00010101001: data <= 32'hb80cbc95;
    11'b00010101010: data <= 32'h35c7bdaf;
    11'b00010101011: data <= 32'h4036b537;
    11'b00010101100: data <= 32'h40da3b2f;
    11'b00010101101: data <= 32'h3b13386f;
    11'b00010101110: data <= 32'hb9cabafa;
    11'b00010101111: data <= 32'hbc8abd3c;
    11'b00010110000: data <= 32'hbbfab4ba;
    11'b00010110001: data <= 32'hbc67340f;
    11'b00010110010: data <= 32'hbb80bb2d;
    11'b00010110011: data <= 32'ha671c054;
    11'b00010110100: data <= 32'h3953bd8b;
    11'b00010110101: data <= 32'h2a643b7c;
    11'b00010110110: data <= 32'hbc5540a5;
    11'b00010110111: data <= 32'hbc473f11;
    11'b00010111000: data <= 32'ha8533981;
    11'b00010111001: data <= 32'h32783662;
    11'b00010111010: data <= 32'hbaea365f;
    11'b00010111011: data <= 32'hbd42ae4e;
    11'b00010111100: data <= 32'h3529b7f1;
    11'b00010111101: data <= 32'h411f28cf;
    11'b00010111110: data <= 32'h41ac3a90;
    11'b00010111111: data <= 32'h3c3d38d0;
    11'b00011000000: data <= 32'hb783b485;
    11'b00011000001: data <= 32'hb6d0b620;
    11'b00011000010: data <= 32'h2e7334d4;
    11'b00011000011: data <= 32'hb04d2ab5;
    11'b00011000100: data <= 32'hb8a5bedb;
    11'b00011000101: data <= 32'hb373c1ff;
    11'b00011000110: data <= 32'h36b6bf7c;
    11'b00011000111: data <= 32'h33b638c3;
    11'b00011001000: data <= 32'hb83e3ecf;
    11'b00011001001: data <= 32'hb9dc3a73;
    11'b00011001010: data <= 32'hb6d3b0ed;
    11'b00011001011: data <= 32'hbabf322e;
    11'b00011001100: data <= 32'hbfe43ad6;
    11'b00011001101: data <= 32'hbff03811;
    11'b00011001110: data <= 32'h282ab474;
    11'b00011001111: data <= 32'h406bb14c;
    11'b00011010000: data <= 32'h406a3995;
    11'b00011010001: data <= 32'h37bc3c56;
    11'b00011010010: data <= 32'hb74e3a84;
    11'b00011010011: data <= 32'h34c73a56;
    11'b00011010100: data <= 32'h3c3a3be1;
    11'b00011010101: data <= 32'h36f73187;
    11'b00011010110: data <= 32'hb856befb;
    11'b00011010111: data <= 32'hb47bc1a6;
    11'b00011011000: data <= 32'h3ab8be9a;
    11'b00011011001: data <= 32'h3cdc35e0;
    11'b00011011010: data <= 32'h38243a62;
    11'b00011011011: data <= 32'hb26db61d;
    11'b00011011100: data <= 32'hb884bba6;
    11'b00011011101: data <= 32'hbd212ae8;
    11'b00011011110: data <= 32'hc08a3bff;
    11'b00011011111: data <= 32'hc03f353d;
    11'b00011100000: data <= 32'hb59fbbd3;
    11'b00011100001: data <= 32'h3d1dbbb5;
    11'b00011100010: data <= 32'h3be43686;
    11'b00011100011: data <= 32'hb6093e0b;
    11'b00011100100: data <= 32'hb87c3e76;
    11'b00011100101: data <= 32'h39673dda;
    11'b00011100110: data <= 32'h3d083d86;
    11'b00011100111: data <= 32'h2fc238cb;
    11'b00011101000: data <= 32'hbc31bb9f;
    11'b00011101001: data <= 32'hb591bf25;
    11'b00011101010: data <= 32'h3df9bb6a;
    11'b00011101011: data <= 32'h4089351f;
    11'b00011101100: data <= 32'h3da33053;
    11'b00011101101: data <= 32'h3483bc0a;
    11'b00011101110: data <= 32'hb404bc42;
    11'b00011101111: data <= 32'hba3434a0;
    11'b00011110000: data <= 32'hbe4a3b9e;
    11'b00011110001: data <= 32'hbebcb64b;
    11'b00011110010: data <= 32'hb8ffc03d;
    11'b00011110011: data <= 32'h35a5bfa5;
    11'b00011110100: data <= 32'h1b4e1eaf;
    11'b00011110101: data <= 32'hbab73ddb;
    11'b00011110110: data <= 32'hb8213e05;
    11'b00011110111: data <= 32'h393d3cb7;
    11'b00011111000: data <= 32'h39633d16;
    11'b00011111001: data <= 32'hbb403c64;
    11'b00011111010: data <= 32'hbf9c30e8;
    11'b00011111011: data <= 32'hb880b8d4;
    11'b00011111100: data <= 32'h3f31b466;
    11'b00011111101: data <= 32'h4139354f;
    11'b00011111110: data <= 32'h3e239d64;
    11'b00011111111: data <= 32'h370db9e1;
    11'b00100000000: data <= 32'h35f1b55f;
    11'b00100000001: data <= 32'h35fd3b70;
    11'b00100000010: data <= 32'hb5e83ba3;
    11'b00100000011: data <= 32'hbc28bc16;
    11'b00100000100: data <= 32'hb9c0c1bf;
    11'b00100000101: data <= 32'hab6fc0c3;
    11'b00100000110: data <= 32'hafdbb4b9;
    11'b00100000111: data <= 32'hb80b3b22;
    11'b00100001000: data <= 32'hb0bd37ee;
    11'b00100001001: data <= 32'h37b8300a;
    11'b00100001010: data <= 32'hb0e53a57;
    11'b00100001011: data <= 32'hbfb43db3;
    11'b00100001100: data <= 32'hc12c3b38;
    11'b00100001101: data <= 32'hbaf7ac61;
    11'b00100001110: data <= 32'h3dcfb375;
    11'b00100001111: data <= 32'h3fb93266;
    11'b00100010000: data <= 32'h3a373403;
    11'b00100010001: data <= 32'h32912f75;
    11'b00100010010: data <= 32'h3bb639e7;
    11'b00100010011: data <= 32'h3dd03e9e;
    11'b00100010100: data <= 32'h381c3c96;
    11'b00100010101: data <= 32'hb9dcbc11;
    11'b00100010110: data <= 32'hb9f8c14d;
    11'b00100010111: data <= 32'h307bc007;
    11'b00100011000: data <= 32'h38abb4fb;
    11'b00100011001: data <= 32'h36c62f06;
    11'b00100011010: data <= 32'h3717ba6b;
    11'b00100011011: data <= 32'h376fbbdb;
    11'b00100011100: data <= 32'hb82135dc;
    11'b00100011101: data <= 32'hc0593e14;
    11'b00100011110: data <= 32'hc13d3b75;
    11'b00100011111: data <= 32'hbc5ab7b4;
    11'b00100100000: data <= 32'h3901bb1c;
    11'b00100100001: data <= 32'h38e1b0f8;
    11'b00100100010: data <= 32'hb60e3826;
    11'b00100100011: data <= 32'hb2403a6d;
    11'b00100100100: data <= 32'h3d0f3d73;
    11'b00100100101: data <= 32'h3f683ff6;
    11'b00100100110: data <= 32'h38033dd6;
    11'b00100100111: data <= 32'hbc45b4de;
    11'b00100101000: data <= 32'hbaf9be16;
    11'b00100101001: data <= 32'h38dbbc0c;
    11'b00100101010: data <= 32'h3df4abd4;
    11'b00100101011: data <= 32'h3d11b758;
    11'b00100101100: data <= 32'h3b46be76;
    11'b00100101101: data <= 32'h39c6bda0;
    11'b00100101110: data <= 32'hab933668;
    11'b00100101111: data <= 32'hbd963e0d;
    11'b00100110000: data <= 32'hbfb9369a;
    11'b00100110001: data <= 32'hbc4cbdc7;
    11'b00100110010: data <= 32'hb245bf20;
    11'b00100110011: data <= 32'hb862b89c;
    11'b00100110100: data <= 32'hbcad378a;
    11'b00100110101: data <= 32'hb62039b0;
    11'b00100110110: data <= 32'h3d0e3c0c;
    11'b00100110111: data <= 32'h3de73ead;
    11'b00100111000: data <= 32'hb51d3ec9;
    11'b00100111001: data <= 32'hbf6a398f;
    11'b00100111010: data <= 32'hbc87b186;
    11'b00100111011: data <= 32'h3ae3a5dd;
    11'b00100111100: data <= 32'h3f4332c8;
    11'b00100111101: data <= 32'h3d5bb8c1;
    11'b00100111110: data <= 32'h3b37be37;
    11'b00100111111: data <= 32'h3c7cbb48;
    11'b00101000000: data <= 32'h3bea3ba3;
    11'b00101000001: data <= 32'ha91a3e4e;
    11'b00101000010: data <= 32'hbb94afed;
    11'b00101000011: data <= 32'hbb11c04e;
    11'b00101000100: data <= 32'hb89ec06b;
    11'b00101000101: data <= 32'hbb1fba15;
    11'b00101000110: data <= 32'hbc642cbf;
    11'b00101000111: data <= 32'hb016b2c7;
    11'b00101001000: data <= 32'h3ca0b1c2;
    11'b00101001001: data <= 32'h3a333ae3;
    11'b00101001010: data <= 32'hbd0f3ee6;
    11'b00101001011: data <= 32'hc1033d92;
    11'b00101001100: data <= 32'hbd7a38a2;
    11'b00101001101: data <= 32'h391e34fe;
    11'b00101001110: data <= 32'h3cd03343;
    11'b00101001111: data <= 32'h3757b663;
    11'b00101010000: data <= 32'h35c5bad7;
    11'b00101010001: data <= 32'h3daa2bed;
    11'b00101010010: data <= 32'h40013e9d;
    11'b00101010011: data <= 32'h3c3b3ef7;
    11'b00101010100: data <= 32'hb51bb235;
    11'b00101010101: data <= 32'hb9cdbfe9;
    11'b00101010110: data <= 32'hb6d3bef4;
    11'b00101010111: data <= 32'hb5c1b806;
    11'b00101011000: data <= 32'hb4d3b6d0;
    11'b00101011001: data <= 32'h36fcbdbf;
    11'b00101011010: data <= 32'h3c98bdff;
    11'b00101011011: data <= 32'h36202df4;
    11'b00101011100: data <= 32'hbe2d3e63;
    11'b00101011101: data <= 32'hc0eb3dcd;
    11'b00101011110: data <= 32'hbd6a35c2;
    11'b00101011111: data <= 32'h2c72b193;
    11'b00101100000: data <= 32'ha9d4ad9f;
    11'b00101100001: data <= 32'hbb37b164;
    11'b00101100010: data <= 32'hb64fb1da;
    11'b00101100011: data <= 32'h3ddc3998;
    11'b00101100100: data <= 32'h40d13fbc;
    11'b00101100101: data <= 32'h3d043f79;
    11'b00101100110: data <= 32'hb72234b9;
    11'b00101100111: data <= 32'hba48bb56;
    11'b00101101000: data <= 32'ha1ffb854;
    11'b00101101001: data <= 32'h37dc2ea1;
    11'b00101101010: data <= 32'h3845b9c8;
    11'b00101101011: data <= 32'h3af7c07d;
    11'b00101101100: data <= 32'h3d16c04a;
    11'b00101101101: data <= 32'h393dafad;
    11'b00101101110: data <= 32'hbaa73df9;
    11'b00101101111: data <= 32'hbe5d3be5;
    11'b00101110000: data <= 32'hbbf2b81d;
    11'b00101110001: data <= 32'hb788bc22;
    11'b00101110010: data <= 32'hbcbfb7e2;
    11'b00101110011: data <= 32'hbfb5b030;
    11'b00101110100: data <= 32'hbaefb037;
    11'b00101110101: data <= 32'h3d523691;
    11'b00101110110: data <= 32'h402c3dd7;
    11'b00101110111: data <= 32'h38683f1f;
    11'b00101111000: data <= 32'hbcad3c0e;
    11'b00101111001: data <= 32'hbc243684;
    11'b00101111010: data <= 32'h3490398b;
    11'b00101111011: data <= 32'h3b5b3992;
    11'b00101111100: data <= 32'h394cb982;
    11'b00101111101: data <= 32'h39f0c074;
    11'b00101111110: data <= 32'h3d86bf2e;
    11'b00101111111: data <= 32'h3dbc3561;
    11'b00110000000: data <= 32'h37e73e28;
    11'b00110000001: data <= 32'hb5bd3706;
    11'b00110000010: data <= 32'hb743bd23;
    11'b00110000011: data <= 32'hb932be09;
    11'b00110000100: data <= 32'hbe46b8b5;
    11'b00110000101: data <= 32'hc010b486;
    11'b00110000110: data <= 32'hb9ffba74;
    11'b00110000111: data <= 32'h3cc5b9f5;
    11'b00110001000: data <= 32'h3d95368a;
    11'b00110001001: data <= 32'hb6bc3dc7;
    11'b00110001010: data <= 32'hbf703ded;
    11'b00110001011: data <= 32'hbcdb3cc5;
    11'b00110001100: data <= 32'h34323cf0;
    11'b00110001101: data <= 32'h38363b2b;
    11'b00110001110: data <= 32'hb1a6b708;
    11'b00110001111: data <= 32'ha6b3be39;
    11'b00110010000: data <= 32'h3d3ebaa5;
    11'b00110010001: data <= 32'h40653c3c;
    11'b00110010010: data <= 32'h3e793eae;
    11'b00110010011: data <= 32'h380932e6;
    11'b00110010100: data <= 32'habf4bd33;
    11'b00110010101: data <= 32'hb6a0bc57;
    11'b00110010110: data <= 32'hbc4fb01d;
    11'b00110010111: data <= 32'hbd1eb6e4;
    11'b00110011000: data <= 32'hb1dcbf1b;
    11'b00110011001: data <= 32'h3cabc02b;
    11'b00110011010: data <= 32'h3b21b8ed;
    11'b00110011011: data <= 32'hbae73c26;
    11'b00110011100: data <= 32'hbf763dae;
    11'b00110011101: data <= 32'hbc1a3c14;
    11'b00110011110: data <= 32'h24f73aa9;
    11'b00110011111: data <= 32'hb78138e2;
    11'b00110100000: data <= 32'hbe36b260;
    11'b00110100001: data <= 32'hbc34ba77;
    11'b00110100010: data <= 32'h3c2cab73;
    11'b00110100011: data <= 32'h40e83d9a;
    11'b00110100100: data <= 32'h3f763ea4;
    11'b00110100101: data <= 32'h3806368b;
    11'b00110100110: data <= 32'haa87b7bf;
    11'b00110100111: data <= 32'h23e32fcd;
    11'b00110101000: data <= 32'hb1cd3a06;
    11'b00110101001: data <= 32'hb56fb62e;
    11'b00110101010: data <= 32'h3511c0cf;
    11'b00110101011: data <= 32'h3cc2c191;
    11'b00110101100: data <= 32'h3b3bbbf6;
    11'b00110101101: data <= 32'hb6283a81;
    11'b00110101110: data <= 32'hbbfb3b67;
    11'b00110101111: data <= 32'hb6573001;
    11'b00110110000: data <= 32'hb14fae35;
    11'b00110110001: data <= 32'hbda73096;
    11'b00110110010: data <= 32'hc146ae0a;
    11'b00110110011: data <= 32'hbeeab84c;
    11'b00110110100: data <= 32'h39e7b005;
    11'b00110110101: data <= 32'h40263b8a;
    11'b00110110110: data <= 32'h3ca53d47;
    11'b00110110111: data <= 32'hb40a3a2a;
    11'b00110111000: data <= 32'hb592390b;
    11'b00110111001: data <= 32'h35ad3dae;
    11'b00110111010: data <= 32'h36d63e59;
    11'b00110111011: data <= 32'h9c9db047;
    11'b00110111100: data <= 32'h3328c09e;
    11'b00110111101: data <= 32'h3c4ec0e7;
    11'b00110111110: data <= 32'h3d58b862;
    11'b00110111111: data <= 32'h39c93b0e;
    11'b00111000000: data <= 32'h34c93593;
    11'b00111000001: data <= 32'h369eba52;
    11'b00111000010: data <= 32'had48ba16;
    11'b00111000011: data <= 32'hbec69e8d;
    11'b00111000100: data <= 32'hc18eab9a;
    11'b00111000101: data <= 32'hbeabbb15;
    11'b00111000110: data <= 32'h38b4bc3b;
    11'b00111000111: data <= 32'h3d70b155;
    11'b00111001000: data <= 32'h2cc23991;
    11'b00111001001: data <= 32'hbc703b84;
    11'b00111001010: data <= 32'hb8c13d2c;
    11'b00111001011: data <= 32'h37b54009;
    11'b00111001100: data <= 32'h355b3f91;
    11'b00111001101: data <= 32'hb8f4316e;
    11'b00111001110: data <= 32'hb8b4be6e;
    11'b00111001111: data <= 32'h39b7bd99;
    11'b00111010000: data <= 32'h3f1a3513;
    11'b00111010001: data <= 32'h3ed33c58;
    11'b00111010010: data <= 32'h3cf31ffe;
    11'b00111010011: data <= 32'h3bb4bc4f;
    11'b00111010100: data <= 32'h3416b87b;
    11'b00111010101: data <= 32'hbca637a5;
    11'b00111010110: data <= 32'hbfdd2cb3;
    11'b00111010111: data <= 32'hbbe9be12;
    11'b00111011000: data <= 32'h3913c07b;
    11'b00111011001: data <= 32'h3a1dbd1e;
    11'b00111011010: data <= 32'hb8e52d45;
    11'b00111011011: data <= 32'hbd5a39cc;
    11'b00111011100: data <= 32'hb6783c45;
    11'b00111011101: data <= 32'h37fb3e59;
    11'b00111011110: data <= 32'hb52e3e24;
    11'b00111011111: data <= 32'hbf4e359f;
    11'b00111100000: data <= 32'hbed5ba53;
    11'b00111100001: data <= 32'h3274b68d;
    11'b00111100010: data <= 32'h3f513b08;
    11'b00111100011: data <= 32'h3f8a3c64;
    11'b00111100100: data <= 32'h3cf5a820;
    11'b00111100101: data <= 32'h3ba1b8bc;
    11'b00111100110: data <= 32'h3936377b;
    11'b00111100111: data <= 32'hb2c33dd1;
    11'b00111101000: data <= 32'hbaaf363e;
    11'b00111101001: data <= 32'hb463bfa0;
    11'b00111101010: data <= 32'h39a0c1b7;
    11'b00111101011: data <= 32'h3897bec6;
    11'b00111101100: data <= 32'hb744b1b1;
    11'b00111101101: data <= 32'hb9473341;
    11'b00111101110: data <= 32'h35022ffb;
    11'b00111101111: data <= 32'h38ce37f5;
    11'b00111110000: data <= 32'hbbfe3af1;
    11'b00111110001: data <= 32'hc1a23640;
    11'b00111110010: data <= 32'hc0e6b58f;
    11'b00111110011: data <= 32'hb249b161;
    11'b00111110100: data <= 32'h3d9e38ff;
    11'b00111110101: data <= 32'h3c88397f;
    11'b00111110110: data <= 32'h35b428e7;
    11'b00111110111: data <= 32'h37b63379;
    11'b00111111000: data <= 32'h3b563ea7;
    11'b00111111001: data <= 32'h385240c2;
    11'b00111111010: data <= 32'hb2a03a4f;
    11'b00111111011: data <= 32'hb0c4bee2;
    11'b00111111100: data <= 32'h385bc0f3;
    11'b00111111101: data <= 32'h39c7bc9e;
    11'b00111111110: data <= 32'h35982772;
    11'b00111111111: data <= 32'h3832b481;
    11'b01000000000: data <= 32'h3cefbb48;
    11'b01000000001: data <= 32'h3b07b711;
    11'b01000000010: data <= 32'hbc9637d0;
    11'b01000000011: data <= 32'hc1cf370c;
    11'b01000000100: data <= 32'hc0abb6dc;
    11'b01000000101: data <= 32'hb40eba4c;
    11'b01000000110: data <= 32'h39eeb5b9;
    11'b01000000111: data <= 32'hab64ab87;
    11'b01000001000: data <= 32'hba0ca6ed;
    11'b01000001001: data <= 32'h14a539cf;
    11'b01000001010: data <= 32'h3c1e406b;
    11'b01000001011: data <= 32'h39874158;
    11'b01000001100: data <= 32'hb8083c34;
    11'b01000001101: data <= 32'hba84bc2f;
    11'b01000001110: data <= 32'h2c08bd52;
    11'b01000001111: data <= 32'h3b32ab5f;
    11'b01000010000: data <= 32'h3c84376e;
    11'b01000010001: data <= 32'h3da4b8b0;
    11'b01000010010: data <= 32'h3f43bdab;
    11'b01000010011: data <= 32'h3ceeb879;
    11'b01000010100: data <= 32'hb8e73a70;
    11'b01000010101: data <= 32'hc006396f;
    11'b01000010110: data <= 32'hbdd0ba47;
    11'b01000010111: data <= 32'h219cbef4;
    11'b01000011000: data <= 32'h3246bda9;
    11'b01000011001: data <= 32'hbb89b9f4;
    11'b01000011010: data <= 32'hbd33b513;
    11'b01000011011: data <= 32'h12dc376d;
    11'b01000011100: data <= 32'h3c863ed6;
    11'b01000011101: data <= 32'h34fe404c;
    11'b01000011110: data <= 32'hbdd53c28;
    11'b01000011111: data <= 32'hbf7cb48a;
    11'b01000100000: data <= 32'hb86cb118;
    11'b01000100001: data <= 32'h3a953a8c;
    11'b01000100010: data <= 32'h3cf23982;
    11'b01000100011: data <= 32'h3d6cb979;
    11'b01000100100: data <= 32'h3ebebcd3;
    11'b01000100101: data <= 32'h3de33259;
    11'b01000100110: data <= 32'h34953ed2;
    11'b01000100111: data <= 32'hb9be3c78;
    11'b01000101000: data <= 32'hb6e2bbfa;
    11'b01000101001: data <= 32'h34f6c080;
    11'b01000101010: data <= 32'ha6bebf22;
    11'b01000101011: data <= 32'hbc34bb7a;
    11'b01000101100: data <= 32'hbb44b9a8;
    11'b01000101101: data <= 32'h38ffb70a;
    11'b01000101110: data <= 32'h3d733793;
    11'b01000101111: data <= 32'hb0e73cc0;
    11'b01000110000: data <= 32'hc0a03ab1;
    11'b01000110001: data <= 32'hc1273151;
    11'b01000110010: data <= 32'hbb74356e;
    11'b01000110011: data <= 32'h37383af0;
    11'b01000110100: data <= 32'h38053652;
    11'b01000110101: data <= 32'h3588b9ed;
    11'b01000110110: data <= 32'h3b90b8ec;
    11'b01000110111: data <= 32'h3dfc3cef;
    11'b01000111000: data <= 32'h3c194133;
    11'b01000111001: data <= 32'h31063e2d;
    11'b01000111010: data <= 32'h23afba78;
    11'b01000111011: data <= 32'h34c8bf71;
    11'b01000111100: data <= 32'h1e5dbc8b;
    11'b01000111101: data <= 32'hb7feb7e9;
    11'b01000111110: data <= 32'h2dd9bbeb;
    11'b01000111111: data <= 32'h3e15bdcc;
    11'b01001000000: data <= 32'h3ed5b997;
    11'b01001000001: data <= 32'hb3e9379e;
    11'b01001000010: data <= 32'hc0be39a8;
    11'b01001000011: data <= 32'hc0bf31c6;
    11'b01001000100: data <= 32'hba63a413;
    11'b01001000101: data <= 32'ha40c2e21;
    11'b01001000110: data <= 32'hb949b524;
    11'b01001000111: data <= 32'hbbe4bb40;
    11'b01001001000: data <= 32'h3010b321;
    11'b01001001001: data <= 32'h3d9c3eea;
    11'b01001001010: data <= 32'h3cfd41a9;
    11'b01001001011: data <= 32'h30273ea9;
    11'b01001001100: data <= 32'hb695b4b2;
    11'b01001001101: data <= 32'hb065b9e9;
    11'b01001001110: data <= 32'h2bff314c;
    11'b01001001111: data <= 32'h306f3462;
    11'b01001010000: data <= 32'h3b41bc46;
    11'b01001010001: data <= 32'h4020c002;
    11'b01001010010: data <= 32'h3fe6bc5a;
    11'b01001010011: data <= 32'h31753831;
    11'b01001010100: data <= 32'hbdf93aff;
    11'b01001010101: data <= 32'hbd38a9fa;
    11'b01001010110: data <= 32'hb2deba55;
    11'b01001010111: data <= 32'hb53cbaf4;
    11'b01001011000: data <= 32'hbe4fbbe9;
    11'b01001011001: data <= 32'hbf37bca7;
    11'b01001011010: data <= 32'hb167b6a7;
    11'b01001011011: data <= 32'h3d9a3cf1;
    11'b01001011100: data <= 32'h3bf1404a;
    11'b01001011101: data <= 32'hb8f83d6f;
    11'b01001011110: data <= 32'hbd66339f;
    11'b01001011111: data <= 32'hb9fa3744;
    11'b01001100000: data <= 32'ha7e63d42;
    11'b01001100001: data <= 32'h34433a8b;
    11'b01001100010: data <= 32'h3accbc21;
    11'b01001100011: data <= 32'h3f34bfa3;
    11'b01001100100: data <= 32'h3fd4b870;
    11'b01001100101: data <= 32'h3ad33d1d;
    11'b01001100110: data <= 32'hb1ea3d3c;
    11'b01001100111: data <= 32'ha197b27d;
    11'b01001101000: data <= 32'h36ccbd1c;
    11'b01001101001: data <= 32'hb629bce6;
    11'b01001101010: data <= 32'hbf28bc53;
    11'b01001101011: data <= 32'hbe9ebd60;
    11'b01001101100: data <= 32'h3471bc82;
    11'b01001101101: data <= 32'h3e7aa0fd;
    11'b01001101110: data <= 32'h38e43b5c;
    11'b01001101111: data <= 32'hbda43a6e;
    11'b01001110000: data <= 32'hc00f37f7;
    11'b01001110001: data <= 32'hbc3f3c2c;
    11'b01001110010: data <= 32'hb3ea3e81;
    11'b01001110011: data <= 32'hb4ed39e4;
    11'b01001110100: data <= 32'hb153bc3b;
    11'b01001110101: data <= 32'h3a84bdad;
    11'b01001110110: data <= 32'h3e853616;
    11'b01001110111: data <= 32'h3d884045;
    11'b01001111000: data <= 32'h3a283ecc;
    11'b01001111001: data <= 32'h39b9af68;
    11'b01001111010: data <= 32'h3950bc09;
    11'b01001111011: data <= 32'hb4c1b895;
    11'b01001111100: data <= 32'hbd65b6c0;
    11'b01001111101: data <= 32'hba4bbd2b;
    11'b01001111110: data <= 32'h3c79bfaf;
    11'b01001111111: data <= 32'h3fcebd01;
    11'b01010000000: data <= 32'h3771ada3;
    11'b01010000001: data <= 32'hbe363628;
    11'b01010000010: data <= 32'hbf4c36d1;
    11'b01010000011: data <= 32'hb9ef3a70;
    11'b01010000100: data <= 32'hb68c3c13;
    11'b01010000101: data <= 32'hbd0a2e53;
    11'b01010000110: data <= 32'hbe3dbce6;
    11'b01010000111: data <= 32'hb4eabc12;
    11'b01010001000: data <= 32'h3cdb3b65;
    11'b01010001001: data <= 32'h3df240ba;
    11'b01010001010: data <= 32'h3ae03eaf;
    11'b01010001011: data <= 32'h37ca3045;
    11'b01010001100: data <= 32'h356bad66;
    11'b01010001101: data <= 32'hb3d73a45;
    11'b01010001110: data <= 32'hb9e83932;
    11'b01010001111: data <= 32'h298cbc1b;
    11'b01010010000: data <= 32'h3ea7c0a8;
    11'b01010010001: data <= 32'h4037bf05;
    11'b01010010010: data <= 32'h394ab456;
    11'b01010010011: data <= 32'hbad0366b;
    11'b01010010100: data <= 32'hb9aa3232;
    11'b01010010101: data <= 32'h30582d7c;
    11'b01010010110: data <= 32'hb5e22cb8;
    11'b01010010111: data <= 32'hc005b890;
    11'b01010011000: data <= 32'hc0fabda4;
    11'b01010011001: data <= 32'hbaeabc25;
    11'b01010011010: data <= 32'h3c1138b0;
    11'b01010011011: data <= 32'h3cd43e90;
    11'b01010011100: data <= 32'h31f33c5b;
    11'b01010011101: data <= 32'hb655350c;
    11'b01010011110: data <= 32'hb43a3b73;
    11'b01010011111: data <= 32'hb4cd4016;
    11'b01010100000: data <= 32'hb7c13dee;
    11'b01010100001: data <= 32'h2f9dba03;
    11'b01010100010: data <= 32'h3d83c05d;
    11'b01010100011: data <= 32'h3f60bd41;
    11'b01010100100: data <= 32'h3c09363c;
    11'b01010100101: data <= 32'h34693a79;
    11'b01010100110: data <= 32'h399425a6;
    11'b01010100111: data <= 32'h3c59b7b2;
    11'b01010101000: data <= 32'hb0bdb63b;
    11'b01010101001: data <= 32'hc04bb942;
    11'b01010101010: data <= 32'hc0e3bd89;
    11'b01010101011: data <= 32'hb868bdc2;
    11'b01010101100: data <= 32'h3cb8b7a8;
    11'b01010101101: data <= 32'h3a9034f6;
    11'b01010101110: data <= 32'hb92932a4;
    11'b01010101111: data <= 32'hbca0343e;
    11'b01010110000: data <= 32'hb8b23db2;
    11'b01010110001: data <= 32'hb5a840f2;
    11'b01010110010: data <= 32'hba493e4d;
    11'b01010110011: data <= 32'hb9c6b97f;
    11'b01010110100: data <= 32'h34c0bec1;
    11'b01010110101: data <= 32'h3cc0b5e5;
    11'b01010110110: data <= 32'h3cd23d32;
    11'b01010110111: data <= 32'h3c763cdd;
    11'b01010111000: data <= 32'h3e38a235;
    11'b01010111001: data <= 32'h3e2db720;
    11'b01010111010: data <= 32'h2c9e2e28;
    11'b01010111011: data <= 32'hbec72d27;
    11'b01010111100: data <= 32'hbe60bc0f;
    11'b01010111101: data <= 32'h34fdbf8f;
    11'b01010111110: data <= 32'h3e1ebe5c;
    11'b01010111111: data <= 32'h38b5bab8;
    11'b01011000000: data <= 32'hbbd7b78f;
    11'b01011000001: data <= 32'hbc6b2401;
    11'b01011000010: data <= 32'hb2b23ca5;
    11'b01011000011: data <= 32'hb3293fa4;
    11'b01011000100: data <= 32'hbd983b9b;
    11'b01011000101: data <= 32'hbfe6bae8;
    11'b01011000110: data <= 32'hbbc8bcea;
    11'b01011000111: data <= 32'h3795354b;
    11'b01011001000: data <= 32'h3c583eaf;
    11'b01011001001: data <= 32'h3ca93c9b;
    11'b01011001010: data <= 32'h3d98a570;
    11'b01011001011: data <= 32'h3d1a3100;
    11'b01011001100: data <= 32'h303f3d3b;
    11'b01011001101: data <= 32'hbc2f3d32;
    11'b01011001110: data <= 32'hb923b6d3;
    11'b01011001111: data <= 32'h3be7c012;
    11'b01011010000: data <= 32'h3eb1c013;
    11'b01011010001: data <= 32'h3883bc7e;
    11'b01011010010: data <= 32'hb8a4b881;
    11'b01011010011: data <= 32'hb05cb414;
    11'b01011010100: data <= 32'h3a7936ae;
    11'b01011010101: data <= 32'h30e63b06;
    11'b01011010110: data <= 32'hbf6f314c;
    11'b01011010111: data <= 32'hc1aabc3a;
    11'b01011011000: data <= 32'hbe9fbc43;
    11'b01011011001: data <= 32'h2f7a344f;
    11'b01011011010: data <= 32'h39d63c64;
    11'b01011011011: data <= 32'h378a3714;
    11'b01011011100: data <= 32'h376bb195;
    11'b01011011101: data <= 32'h38a53aeb;
    11'b01011011110: data <= 32'h2b1140fa;
    11'b01011011111: data <= 32'hb931408f;
    11'b01011100000: data <= 32'hb50f2b8d;
    11'b01011100001: data <= 32'h3adebf13;
    11'b01011100010: data <= 32'h3d37be4b;
    11'b01011100011: data <= 32'h38b3b71e;
    11'b01011100100: data <= 32'h3372ae3b;
    11'b01011100101: data <= 32'h3cbab66e;
    11'b01011100110: data <= 32'h3fb4b427;
    11'b01011100111: data <= 32'h39063229;
    11'b01011101000: data <= 32'hbf55ad30;
    11'b01011101001: data <= 32'hc185bba3;
    11'b01011101010: data <= 32'hbd70bcab;
    11'b01011101011: data <= 32'h34bbb7af;
    11'b01011101100: data <= 32'h35b3b06c;
    11'b01011101101: data <= 32'hb71cb8ef;
    11'b01011101110: data <= 32'hb7d7b823;
    11'b01011101111: data <= 32'h2e3e3ca1;
    11'b01011110000: data <= 32'h29f741c5;
    11'b01011110001: data <= 32'hb97040da;
    11'b01011110010: data <= 32'hbac73104;
    11'b01011110011: data <= 32'haf80bd10;
    11'b01011110100: data <= 32'h377fb87c;
    11'b01011110101: data <= 32'h37703903;
    11'b01011110110: data <= 32'h3abb3769;
    11'b01011110111: data <= 32'h4003b741;
    11'b01011111000: data <= 32'h40f4b75a;
    11'b01011111001: data <= 32'h3b7b3614;
    11'b01011111010: data <= 32'hbd5f384b;
    11'b01011111011: data <= 32'hbf6cb6ad;
    11'b01011111100: data <= 32'hb5ddbd23;
    11'b01011111101: data <= 32'h3a47bd58;
    11'b01011111110: data <= 32'h300cbd04;
    11'b01011111111: data <= 32'hbbd9bdb7;
    11'b01100000000: data <= 32'hb9c7bb47;
    11'b01100000001: data <= 32'h35723a99;
    11'b01100000010: data <= 32'h352c408e;
    11'b01100000011: data <= 32'hbbae3ed5;
    11'b01100000100: data <= 32'hbf4eb057;
    11'b01100000101: data <= 32'hbd64ba8c;
    11'b01100000110: data <= 32'hb69034fd;
    11'b01100000111: data <= 32'h30be3d11;
    11'b01100001000: data <= 32'h3a4b3863;
    11'b01100001001: data <= 32'h3f44b8a7;
    11'b01100001010: data <= 32'h4050b1b1;
    11'b01100001011: data <= 32'h3b4d3d3b;
    11'b01100001100: data <= 32'hb9a93ed6;
    11'b01100001101: data <= 32'hba0a35b9;
    11'b01100001110: data <= 32'h387fbcbf;
    11'b01100001111: data <= 32'h3c5cbe93;
    11'b01100010000: data <= 32'h2220be0e;
    11'b01100010001: data <= 32'hbb0fbe0f;
    11'b01100010010: data <= 32'ha94fbc91;
    11'b01100010011: data <= 32'h3d332d78;
    11'b01100010100: data <= 32'h3b2b3c79;
    11'b01100010101: data <= 32'hbc903984;
    11'b01100010110: data <= 32'hc107b7fd;
    11'b01100010111: data <= 32'hc008b8c0;
    11'b01100011000: data <= 32'hba81383d;
    11'b01100011001: data <= 32'hb3303be2;
    11'b01100011010: data <= 32'h2d0ead8c;
    11'b01100011011: data <= 32'h3a36bb6e;
    11'b01100011100: data <= 32'h3d053355;
    11'b01100011101: data <= 32'h39534096;
    11'b01100011110: data <= 32'hb464415c;
    11'b01100011111: data <= 32'hb1773b7d;
    11'b01100100000: data <= 32'h39d2bac3;
    11'b01100100001: data <= 32'h3a86bc91;
    11'b01100100010: data <= 32'hb0b0ba03;
    11'b01100100011: data <= 32'hb61ebb09;
    11'b01100100100: data <= 32'h3c40bc87;
    11'b01100100101: data <= 32'h40d4b8de;
    11'b01100100110: data <= 32'h3e053258;
    11'b01100100111: data <= 32'hbbe530ae;
    11'b01100101000: data <= 32'hc0c1b822;
    11'b01100101001: data <= 32'hbe9fb844;
    11'b01100101010: data <= 32'hb8112e39;
    11'b01100101011: data <= 32'hb77ba544;
    11'b01100101100: data <= 32'hbac1bc93;
    11'b01100101101: data <= 32'hb638bdc2;
    11'b01100101110: data <= 32'h37a6358c;
    11'b01100101111: data <= 32'h38184133;
    11'b01100110000: data <= 32'hb1734192;
    11'b01100110001: data <= 32'hb6363baa;
    11'b01100110010: data <= 32'h9074b6f2;
    11'b01100110011: data <= 32'ha149afa7;
    11'b01100110100: data <= 32'hb75f3814;
    11'b01100110101: data <= 32'h211da892;
    11'b01100110110: data <= 32'h3f1bbc14;
    11'b01100110111: data <= 32'h41e3bb4f;
    11'b01100111000: data <= 32'h3f282d20;
    11'b01100111001: data <= 32'hb85937fa;
    11'b01100111010: data <= 32'hbdd19e38;
    11'b01100111011: data <= 32'hb7ebb72c;
    11'b01100111100: data <= 32'h33d5b813;
    11'b01100111101: data <= 32'hb834bc06;
    11'b01100111110: data <= 32'hbdd8bfd3;
    11'b01100111111: data <= 32'hbb51bf74;
    11'b01101000000: data <= 32'h370421dd;
    11'b01101000001: data <= 32'h39e43fdb;
    11'b01101000010: data <= 32'hb4053fb0;
    11'b01101000011: data <= 32'hbc6036dc;
    11'b01101000100: data <= 32'hbc53b0f7;
    11'b01101000101: data <= 32'hbb423a85;
    11'b01101000110: data <= 32'hbae53db9;
    11'b01101000111: data <= 32'hae3f3587;
    11'b01101001000: data <= 32'h3e30bc45;
    11'b01101001001: data <= 32'h4104ba8b;
    11'b01101001010: data <= 32'h3e4539c0;
    11'b01101001011: data <= 32'hac023dfe;
    11'b01101001100: data <= 32'hb4d93a5c;
    11'b01101001101: data <= 32'h39a0b310;
    11'b01101001110: data <= 32'h3ad9b9b9;
    11'b01101001111: data <= 32'hb840bcdb;
    11'b01101010000: data <= 32'hbe1ebfd9;
    11'b01101010001: data <= 32'hb840bfc7;
    11'b01101010010: data <= 32'h3cd1b8c9;
    11'b01101010011: data <= 32'h3d543a18;
    11'b01101010100: data <= 32'hb450392f;
    11'b01101010101: data <= 32'hbe8bb3e0;
    11'b01101010110: data <= 32'hbebcac17;
    11'b01101010111: data <= 32'hbd0f3cb9;
    11'b01101011000: data <= 32'hbc8f3dd0;
    11'b01101011001: data <= 32'hb9adac93;
    11'b01101011010: data <= 32'h377abdb3;
    11'b01101011011: data <= 32'h3d7cb8bd;
    11'b01101011100: data <= 32'h3c0d3e16;
    11'b01101011101: data <= 32'h330340c8;
    11'b01101011110: data <= 32'h36933d70;
    11'b01101011111: data <= 32'h3cb52d64;
    11'b01101100000: data <= 32'h3a9bb443;
    11'b01101100001: data <= 32'hb973b69d;
    11'b01101100010: data <= 32'hbce1bc79;
    11'b01101100011: data <= 32'h35ccbe94;
    11'b01101100100: data <= 32'h4073bc86;
    11'b01101100101: data <= 32'h3fd0b45c;
    11'b01101100110: data <= 32'hae2bb2ad;
    11'b01101100111: data <= 32'hbe08b849;
    11'b01101101000: data <= 32'hbd23a8d0;
    11'b01101101001: data <= 32'hba4b3b84;
    11'b01101101010: data <= 32'hbc7f3974;
    11'b01101101011: data <= 32'hbde7bc13;
    11'b01101101100: data <= 32'hba61bfde;
    11'b01101101101: data <= 32'h347fb857;
    11'b01101101110: data <= 32'h387d3f30;
    11'b01101101111: data <= 32'h342340e9;
    11'b01101110000: data <= 32'h36173cfc;
    11'b01101110001: data <= 32'h39a9347f;
    11'b01101110010: data <= 32'h303438e8;
    11'b01101110011: data <= 32'hbc243b7d;
    11'b01101110100: data <= 32'hbb7b2801;
    11'b01101110101: data <= 32'h3c07bcdd;
    11'b01101110110: data <= 32'h416ebd5e;
    11'b01101110111: data <= 32'h4049b88c;
    11'b01101111000: data <= 32'h31d6b063;
    11'b01101111001: data <= 32'hb99eb1f3;
    11'b01101111010: data <= 32'ha98a2d7c;
    11'b01101111011: data <= 32'h3421378e;
    11'b01101111100: data <= 32'hbae2b26c;
    11'b01101111101: data <= 32'hbfe6bf2b;
    11'b01101111110: data <= 32'hbdf6c0ad;
    11'b01101111111: data <= 32'haba8ba22;
    11'b01110000000: data <= 32'h38b73d00;
    11'b01110000001: data <= 32'h32773e14;
    11'b01110000010: data <= 32'hb13c3729;
    11'b01110000011: data <= 32'hb39133d6;
    11'b01110000100: data <= 32'hb9c63dac;
    11'b01110000101: data <= 32'hbdb14007;
    11'b01110000110: data <= 32'hbbe239d8;
    11'b01110000111: data <= 32'h3ab2bc1f;
    11'b01110001000: data <= 32'h406ebcfe;
    11'b01110001001: data <= 32'h3ebaaeac;
    11'b01110001010: data <= 32'h35e1398c;
    11'b01110001011: data <= 32'h350d3879;
    11'b01110001100: data <= 32'h3d383547;
    11'b01110001101: data <= 32'h3ccd342d;
    11'b01110001110: data <= 32'hb8ceb703;
    11'b01110001111: data <= 32'hc009beff;
    11'b01110010000: data <= 32'hbd26c070;
    11'b01110010001: data <= 32'h3808bc71;
    11'b01110010010: data <= 32'h3c6e31a9;
    11'b01110010011: data <= 32'h33022e8f;
    11'b01110010100: data <= 32'hb951b885;
    11'b01110010101: data <= 32'hbab52997;
    11'b01110010110: data <= 32'hbc2e3ef0;
    11'b01110010111: data <= 32'hbe314071;
    11'b01110011000: data <= 32'hbd7d385e;
    11'b01110011001: data <= 32'hafddbd22;
    11'b01110011010: data <= 32'h3b91bc40;
    11'b01110011011: data <= 32'h3a5338f8;
    11'b01110011100: data <= 32'h35693e38;
    11'b01110011101: data <= 32'h3bae3c67;
    11'b01110011110: data <= 32'h3fde383f;
    11'b01110011111: data <= 32'h3dbd3842;
    11'b01110100000: data <= 32'hb8e3341c;
    11'b01110100001: data <= 32'hbefaba4d;
    11'b01110100010: data <= 32'hb7ffbe62;
    11'b01110100011: data <= 32'h3ddabd4c;
    11'b01110100100: data <= 32'h3ed7ba2d;
    11'b01110100101: data <= 32'h3551bb94;
    11'b01110100110: data <= 32'hb950bc9c;
    11'b01110100111: data <= 32'hb837aedf;
    11'b01110101000: data <= 32'hb7813e12;
    11'b01110101001: data <= 32'hbcf23e50;
    11'b01110101010: data <= 32'hbf4db4ed;
    11'b01110101011: data <= 32'hbd2bbf36;
    11'b01110101100: data <= 32'hb56bbbe9;
    11'b01110101101: data <= 32'h21fa3bd0;
    11'b01110101110: data <= 32'h31253ebf;
    11'b01110101111: data <= 32'h3b833b4a;
    11'b01110110000: data <= 32'h3e973784;
    11'b01110110001: data <= 32'h3af23c7a;
    11'b01110110010: data <= 32'hbb753e06;
    11'b01110110011: data <= 32'hbdd9386d;
    11'b01110110100: data <= 32'h31dcba8d;
    11'b01110110101: data <= 32'h4001bd21;
    11'b01110110110: data <= 32'h3f62bc3d;
    11'b01110110111: data <= 32'h365abc30;
    11'b01110111000: data <= 32'hafb1bbc5;
    11'b01110111001: data <= 32'h38eda8de;
    11'b01110111010: data <= 32'h3a113c48;
    11'b01110111011: data <= 32'hb8eb3990;
    11'b01110111100: data <= 32'hc016bc73;
    11'b01110111101: data <= 32'hbfd5c048;
    11'b01110111110: data <= 32'hbaf4bc2e;
    11'b01110111111: data <= 32'hb18b393f;
    11'b01111000000: data <= 32'h24bf3ac1;
    11'b01111000001: data <= 32'h36c9ab40;
    11'b01111000010: data <= 32'h39e92d27;
    11'b01111000011: data <= 32'h1d703e83;
    11'b01111000100: data <= 32'hbd384117;
    11'b01111000101: data <= 32'hbd8f3dd5;
    11'b01111000110: data <= 32'h327fb604;
    11'b01111000111: data <= 32'h3e5fbc40;
    11'b01111001000: data <= 32'h3cf1b8fe;
    11'b01111001001: data <= 32'h33dbb490;
    11'b01111001010: data <= 32'h38c9b3d9;
    11'b01111001011: data <= 32'h3fa93271;
    11'b01111001100: data <= 32'h3fac3a3c;
    11'b01111001101: data <= 32'hab7034e1;
    11'b01111001110: data <= 32'hbfafbca0;
    11'b01111001111: data <= 32'hbf1cbf9a;
    11'b01111010000: data <= 32'hb680bc51;
    11'b01111010001: data <= 32'h34a0b002;
    11'b01111010010: data <= 32'h2728b828;
    11'b01111010011: data <= 32'hafcebd2e;
    11'b01111010100: data <= 32'h259db731;
    11'b01111010101: data <= 32'hb66c3ef9;
    11'b01111010110: data <= 32'hbd5c4187;
    11'b01111010111: data <= 32'hbe033d9f;
    11'b01111011000: data <= 32'hb7a9b83b;
    11'b01111011001: data <= 32'h3619bad7;
    11'b01111011010: data <= 32'h2f7c2fbf;
    11'b01111011011: data <= 32'hb054393c;
    11'b01111011100: data <= 32'h3c0c35f3;
    11'b01111011101: data <= 32'h412c3582;
    11'b01111011110: data <= 32'h40a13a90;
    11'b01111011111: data <= 32'h2d0039ef;
    11'b01111100000: data <= 32'hbe65b42a;
    11'b01111100001: data <= 32'hbbe3bc3c;
    11'b01111100010: data <= 32'h38c2bb73;
    11'b01111100011: data <= 32'h3b9fba92;
    11'b01111100100: data <= 32'h2f00be4b;
    11'b01111100101: data <= 32'hb4e7c027;
    11'b01111100110: data <= 32'h2e6bba5e;
    11'b01111100111: data <= 32'h2e703dca;
    11'b01111101000: data <= 32'hbaa54041;
    11'b01111101001: data <= 32'hbe633858;
    11'b01111101010: data <= 32'hbd86bc5a;
    11'b01111101011: data <= 32'hbb3cba20;
    11'b01111101100: data <= 32'hbb1438f7;
    11'b01111101101: data <= 32'hb8753bef;
    11'b01111101110: data <= 32'h3b0a343d;
    11'b01111101111: data <= 32'h408f2f54;
    11'b01111110000: data <= 32'h3f1d3c44;
    11'b01111110001: data <= 32'hb4103ee0;
    11'b01111110010: data <= 32'hbd3b3c4d;
    11'b01111110011: data <= 32'hb22aa8d7;
    11'b01111110100: data <= 32'h3d40b8ca;
    11'b01111110101: data <= 32'h3cb6bbb7;
    11'b01111110110: data <= 32'h28fcbec7;
    11'b01111110111: data <= 32'hacdabfde;
    11'b01111111000: data <= 32'h3bcbba09;
    11'b01111111001: data <= 32'h3d423be9;
    11'b01111111010: data <= 32'h29a33ca7;
    11'b01111111011: data <= 32'hbdf7b69e;
    11'b01111111100: data <= 32'hbf7cbe15;
    11'b01111111101: data <= 32'hbddab9c1;
    11'b01111111110: data <= 32'hbcbf38a5;
    11'b01111111111: data <= 32'hba33368f;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    