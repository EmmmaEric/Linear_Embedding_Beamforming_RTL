
module memory_rom_43(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hb0f43e4b;
    11'b00000000001: data <= 32'ha7453b4b;
    11'b00000000010: data <= 32'h2f92bb40;
    11'b00000000011: data <= 32'h3bf0be5a;
    11'b00000000100: data <= 32'h3ee5a252;
    11'b00000000101: data <= 32'h3d8f3f93;
    11'b00000000110: data <= 32'h392d3efa;
    11'b00000000111: data <= 32'h3855ab5d;
    11'b00000001000: data <= 32'h38e5bcd2;
    11'b00000001001: data <= 32'hb36abb50;
    11'b00000001010: data <= 32'hbda3b8d8;
    11'b00000001011: data <= 32'hbc74bce5;
    11'b00000001100: data <= 32'h3a06bf02;
    11'b00000001101: data <= 32'h3f79bc69;
    11'b00000001110: data <= 32'h38f72b9a;
    11'b00000001111: data <= 32'hbe103845;
    11'b00000010000: data <= 32'hc01f3819;
    11'b00000010001: data <= 32'hbbd93ade;
    11'b00000010010: data <= 32'hb5413cba;
    11'b00000010011: data <= 32'hbb4f3612;
    11'b00000010100: data <= 32'hbd04bc3b;
    11'b00000010101: data <= 32'hb1e0bc8c;
    11'b00000010110: data <= 32'h3d1b399d;
    11'b00000010111: data <= 32'h3e6540b5;
    11'b00000011000: data <= 32'h3bd63f6d;
    11'b00000011001: data <= 32'h388c30f2;
    11'b00000011010: data <= 32'h36cab6e2;
    11'b00000011011: data <= 32'hb1673523;
    11'b00000011100: data <= 32'hba6b36fc;
    11'b00000011101: data <= 32'hb23ebbc4;
    11'b00000011110: data <= 32'h3dd1c08d;
    11'b00000011111: data <= 32'h4039bf64;
    11'b00000100000: data <= 32'h39d9b60a;
    11'b00000100001: data <= 32'hbc2136bc;
    11'b00000100010: data <= 32'hbc9934e5;
    11'b00000100011: data <= 32'hb24132fa;
    11'b00000100100: data <= 32'hb50433ea;
    11'b00000100101: data <= 32'hbeffb5b5;
    11'b00000100110: data <= 32'hc0c2bd19;
    11'b00000100111: data <= 32'hbba5bc26;
    11'b00000101000: data <= 32'h3be938ed;
    11'b00000101001: data <= 32'h3d9c3f85;
    11'b00000101010: data <= 32'h377d3d96;
    11'b00000101011: data <= 32'hb2a6358a;
    11'b00000101100: data <= 32'hb15938d6;
    11'b00000101101: data <= 32'hb2e43ec6;
    11'b00000101110: data <= 32'hb6d13daa;
    11'b00000101111: data <= 32'h300ab940;
    11'b00000110000: data <= 32'h3dabc089;
    11'b00000110001: data <= 32'h3fdabe90;
    11'b00000110010: data <= 32'h3c2f2e74;
    11'b00000110011: data <= 32'h27123a22;
    11'b00000110100: data <= 32'h34352f9d;
    11'b00000110101: data <= 32'h3a8eb70b;
    11'b00000110110: data <= 32'hae72b6a5;
    11'b00000110111: data <= 32'hc01cb931;
    11'b00000111000: data <= 32'hc138bd4b;
    11'b00000111001: data <= 32'hbaf0bd66;
    11'b00000111010: data <= 32'h3c4ab4b3;
    11'b00000111011: data <= 32'h3c1f3922;
    11'b00000111100: data <= 32'hb62d3837;
    11'b00000111101: data <= 32'hbc5c354d;
    11'b00000111110: data <= 32'hb9083d0c;
    11'b00000111111: data <= 32'hb4a540c7;
    11'b00001000000: data <= 32'hb8a53ef1;
    11'b00001000001: data <= 32'hb7d3b835;
    11'b00001000010: data <= 32'h3805bf5f;
    11'b00001000011: data <= 32'h3d78ba20;
    11'b00001000100: data <= 32'h3d1d3c22;
    11'b00001000101: data <= 32'h3bea3cf6;
    11'b00001000110: data <= 32'h3d582bf8;
    11'b00001000111: data <= 32'h3ddbb8b0;
    11'b00001001000: data <= 32'h30b3b23c;
    11'b00001001001: data <= 32'hbef2af59;
    11'b00001001010: data <= 32'hbfb3bc1a;
    11'b00001001011: data <= 32'had08bf35;
    11'b00001001100: data <= 32'h3db6bdd2;
    11'b00001001101: data <= 32'h3a11b920;
    11'b00001001110: data <= 32'hbb31b45d;
    11'b00001001111: data <= 32'hbd352eab;
    11'b00001010000: data <= 32'hb7423cbf;
    11'b00001010001: data <= 32'hb29b4022;
    11'b00001010010: data <= 32'hbc873d09;
    11'b00001010011: data <= 32'hbecbb95c;
    11'b00001010100: data <= 32'hba6fbd70;
    11'b00001010101: data <= 32'h38d72c24;
    11'b00001010110: data <= 32'h3ce53e7f;
    11'b00001010111: data <= 32'h3d093d61;
    11'b00001011000: data <= 32'h3dd22b04;
    11'b00001011001: data <= 32'h3d83afbe;
    11'b00001011010: data <= 32'h33d43b00;
    11'b00001011011: data <= 32'hbc6f3c35;
    11'b00001011100: data <= 32'hbb65b713;
    11'b00001011101: data <= 32'h39e0c00f;
    11'b00001011110: data <= 32'h3ebac03c;
    11'b00001011111: data <= 32'h3983bcc5;
    11'b00001100000: data <= 32'hb994b84d;
    11'b00001100001: data <= 32'hb86eb197;
    11'b00001100010: data <= 32'h371d383f;
    11'b00001100011: data <= 32'h307c3c55;
    11'b00001100100: data <= 32'hbe9936ec;
    11'b00001100101: data <= 32'hc173bb49;
    11'b00001100110: data <= 32'hbed7bc79;
    11'b00001100111: data <= 32'h2f573361;
    11'b00001101000: data <= 32'h3b493d40;
    11'b00001101001: data <= 32'h39d33a52;
    11'b00001101010: data <= 32'h394facc8;
    11'b00001101011: data <= 32'h39d138b3;
    11'b00001101100: data <= 32'h316d4048;
    11'b00001101101: data <= 32'hb902405c;
    11'b00001101110: data <= 32'hb61b2fbd;
    11'b00001101111: data <= 32'h3ae4bf6e;
    11'b00001110000: data <= 32'h3dd9bf87;
    11'b00001110001: data <= 32'h39a0b9da;
    11'b00001110010: data <= 32'h28cbb18d;
    11'b00001110011: data <= 32'h39f5b575;
    11'b00001110100: data <= 32'h3e7bb28f;
    11'b00001110101: data <= 32'h391d3367;
    11'b00001110110: data <= 32'hbf02a5ab;
    11'b00001110111: data <= 32'hc1d5bb58;
    11'b00001111000: data <= 32'hbeb0bca4;
    11'b00001111001: data <= 32'h316db5c6;
    11'b00001111010: data <= 32'h384d3249;
    11'b00001111011: data <= 32'hb1e3b3cf;
    11'b00001111100: data <= 32'hb602b676;
    11'b00001111101: data <= 32'h2f023c07;
    11'b00001111110: data <= 32'h2ee24195;
    11'b00001111111: data <= 32'hb85e412b;
    11'b00010000000: data <= 32'hb988354f;
    11'b00010000001: data <= 32'h2d09bd9c;
    11'b00010000010: data <= 32'h39acbbaf;
    11'b00010000011: data <= 32'h38d53535;
    11'b00010000100: data <= 32'h39e03712;
    11'b00010000101: data <= 32'h3f12b639;
    11'b00010000110: data <= 32'h40c3b864;
    11'b00010000111: data <= 32'h3c16313b;
    11'b00010001000: data <= 32'hbd7835e1;
    11'b00010001001: data <= 32'hc062b7ad;
    11'b00010001010: data <= 32'hba57bd1c;
    11'b00010001011: data <= 32'h3925bcf3;
    11'b00010001100: data <= 32'h3494bc1f;
    11'b00010001101: data <= 32'hbae5bcc6;
    11'b00010001110: data <= 32'hbad9ba90;
    11'b00010001111: data <= 32'h301d3aa1;
    11'b00010010000: data <= 32'h34de40de;
    11'b00010010001: data <= 32'hba30401b;
    11'b00010010010: data <= 32'hbe6a2e7f;
    11'b00010010011: data <= 32'hbca8bb84;
    11'b00010010100: data <= 32'hb343201e;
    11'b00010010101: data <= 32'h34fc3ca7;
    11'b00010010110: data <= 32'h3ae739b1;
    11'b00010010111: data <= 32'h3f6eb7aa;
    11'b00010011000: data <= 32'h4092b62d;
    11'b00010011001: data <= 32'h3c4c3b77;
    11'b00010011010: data <= 32'hba043dd6;
    11'b00010011011: data <= 32'hbc4d349c;
    11'b00010011100: data <= 32'h33ecbce8;
    11'b00010011101: data <= 32'h3c46bee5;
    11'b00010011110: data <= 32'h313abe3c;
    11'b00010011111: data <= 32'hbb7fbdfa;
    11'b00010100000: data <= 32'hb684bc6c;
    11'b00010100001: data <= 32'h3b813160;
    11'b00010100010: data <= 32'h3aaf3d69;
    11'b00010100011: data <= 32'hbbe73c1a;
    11'b00010100100: data <= 32'hc0dab4f8;
    11'b00010100101: data <= 32'hc019b95d;
    11'b00010100110: data <= 32'hba6636cf;
    11'b00010100111: data <= 32'hac3c3c99;
    11'b00010101000: data <= 32'h34d53433;
    11'b00010101001: data <= 32'h3be6ba42;
    11'b00010101010: data <= 32'h3ddd1e94;
    11'b00010101011: data <= 32'h3ab33fe2;
    11'b00010101100: data <= 32'hb4304123;
    11'b00010101101: data <= 32'hb4e53bcd;
    11'b00010101110: data <= 32'h395bbb78;
    11'b00010101111: data <= 32'h3bcdbdb6;
    11'b00010110000: data <= 32'h25d2bc25;
    11'b00010110001: data <= 32'hb82bbc02;
    11'b00010110010: data <= 32'h392dbc88;
    11'b00010110011: data <= 32'h4030b882;
    11'b00010110100: data <= 32'h3df734c7;
    11'b00010110101: data <= 32'hbb54347a;
    11'b00010110110: data <= 32'hc10db777;
    11'b00010110111: data <= 32'hbfdeb8aa;
    11'b00010111000: data <= 32'hb95230be;
    11'b00010111001: data <= 32'hb56234a9;
    11'b00010111010: data <= 32'hb8d6b9f9;
    11'b00010111011: data <= 32'hb35dbd2c;
    11'b00010111100: data <= 32'h388932ae;
    11'b00010111101: data <= 32'h38db4101;
    11'b00010111110: data <= 32'had3e41e3;
    11'b00010111111: data <= 32'hb4fb3ca0;
    11'b00011000000: data <= 32'h3117b846;
    11'b00011000001: data <= 32'h3426b804;
    11'b00011000010: data <= 32'hb45431aa;
    11'b00011000011: data <= 32'hacd3affc;
    11'b00011000100: data <= 32'h3e1ebc01;
    11'b00011000101: data <= 32'h41b0bbd3;
    11'b00011000110: data <= 32'h3f96ab98;
    11'b00011000111: data <= 32'hb84b3620;
    11'b00011001000: data <= 32'hbf20ada5;
    11'b00011001001: data <= 32'hbb9fb80c;
    11'b00011001010: data <= 32'h29a9b738;
    11'b00011001011: data <= 32'hb690ba31;
    11'b00011001100: data <= 32'hbd52becd;
    11'b00011001101: data <= 32'hbbe0bf22;
    11'b00011001110: data <= 32'h349ca42a;
    11'b00011001111: data <= 32'h39bb4038;
    11'b00011010000: data <= 32'hb00d409a;
    11'b00011010001: data <= 32'hbb7139cf;
    11'b00011010010: data <= 32'hbb35b38d;
    11'b00011010011: data <= 32'hb9853801;
    11'b00011010100: data <= 32'hb9793d17;
    11'b00011010101: data <= 32'ha9cc3735;
    11'b00011010110: data <= 32'h3e45bbce;
    11'b00011010111: data <= 32'h4154bbd2;
    11'b00011011000: data <= 32'h3f2c368a;
    11'b00011011001: data <= 32'habf33d14;
    11'b00011011010: data <= 32'hb918398b;
    11'b00011011011: data <= 32'h3545b4c6;
    11'b00011011100: data <= 32'h3a3aba55;
    11'b00011011101: data <= 32'hb646bcef;
    11'b00011011110: data <= 32'hbe2ebfcc;
    11'b00011011111: data <= 32'hbab7bfdc;
    11'b00011100000: data <= 32'h3af6b88f;
    11'b00011100001: data <= 32'h3cff3c02;
    11'b00011100010: data <= 32'hb12c3c33;
    11'b00011100011: data <= 32'hbe4320a7;
    11'b00011100100: data <= 32'hbecdb010;
    11'b00011100101: data <= 32'hbcf73c24;
    11'b00011100110: data <= 32'hbc103e40;
    11'b00011100111: data <= 32'hb8543405;
    11'b00011101000: data <= 32'h395bbd0c;
    11'b00011101001: data <= 32'h3e93ba30;
    11'b00011101010: data <= 32'h3d0f3cea;
    11'b00011101011: data <= 32'h3420408d;
    11'b00011101100: data <= 32'h336b3d88;
    11'b00011101101: data <= 32'h3c381f92;
    11'b00011101110: data <= 32'h3ba9b81c;
    11'b00011101111: data <= 32'hb7dab971;
    11'b00011110000: data <= 32'hbd45bd26;
    11'b00011110001: data <= 32'ha6a6beea;
    11'b00011110010: data <= 32'h3f9fbc86;
    11'b00011110011: data <= 32'h3fb5b059;
    11'b00011110100: data <= 32'ha6c416b8;
    11'b00011110101: data <= 32'hbe8cb719;
    11'b00011110110: data <= 32'hbe53af07;
    11'b00011110111: data <= 32'hbbc63b85;
    11'b00011111000: data <= 32'hbc413bb8;
    11'b00011111001: data <= 32'hbd29b8ee;
    11'b00011111010: data <= 32'hb8f5bf36;
    11'b00011111011: data <= 32'h3730b969;
    11'b00011111100: data <= 32'h39c13ec2;
    11'b00011111101: data <= 32'h35644137;
    11'b00011111110: data <= 32'h365c3ddf;
    11'b00011111111: data <= 32'h3a993380;
    11'b00100000000: data <= 32'h368c3476;
    11'b00100000001: data <= 32'hba8538c5;
    11'b00100000010: data <= 32'hbc09b00f;
    11'b00100000011: data <= 32'h39fbbd17;
    11'b00100000100: data <= 32'h4137bdac;
    11'b00100000101: data <= 32'h408cb935;
    11'b00100000110: data <= 32'h3387b22a;
    11'b00100000111: data <= 32'hbbf2b439;
    11'b00100001000: data <= 32'hb811a285;
    11'b00100001001: data <= 32'h95103802;
    11'b00100001010: data <= 32'hba8a2946;
    11'b00100001011: data <= 32'hbf7cbe11;
    11'b00100001100: data <= 32'hbe11c08a;
    11'b00100001101: data <= 32'hb08abab5;
    11'b00100001110: data <= 32'h38c03d72;
    11'b00100001111: data <= 32'h34a63fa7;
    11'b00100010000: data <= 32'haa023a6d;
    11'b00100010001: data <= 32'habe23360;
    11'b00100010010: data <= 32'hb7a13c86;
    11'b00100010011: data <= 32'hbcf33f4b;
    11'b00100010100: data <= 32'hbbbf3a2a;
    11'b00100010101: data <= 32'h3a8cbbd4;
    11'b00100010110: data <= 32'h40c3bd8d;
    11'b00100010111: data <= 32'h3fe2b5cd;
    11'b00100011000: data <= 32'h36fc37d3;
    11'b00100011001: data <= 32'h1d6e36f4;
    11'b00100011010: data <= 32'h3b2d3335;
    11'b00100011011: data <= 32'h3c3d3260;
    11'b00100011100: data <= 32'hb808b6ad;
    11'b00100011101: data <= 32'hc00dbeec;
    11'b00100011110: data <= 32'hbe34c097;
    11'b00100011111: data <= 32'h3296bca1;
    11'b00100100000: data <= 32'h3c12363d;
    11'b00100100001: data <= 32'h34b5385c;
    11'b00100100010: data <= 32'hb8d2b3af;
    11'b00100100011: data <= 32'hba9d2669;
    11'b00100100100: data <= 32'hbc013e55;
    11'b00100100101: data <= 32'hbdd74095;
    11'b00100100110: data <= 32'hbd1c3aac;
    11'b00100100111: data <= 32'h2904bc7c;
    11'b00100101000: data <= 32'h3d07bcdf;
    11'b00100101001: data <= 32'h3c81358e;
    11'b00100101010: data <= 32'h36ec3db6;
    11'b00100101011: data <= 32'h3a313c68;
    11'b00100101100: data <= 32'h3f333779;
    11'b00100101101: data <= 32'h3e1f357a;
    11'b00100101110: data <= 32'hb6c428cd;
    11'b00100101111: data <= 32'hbf48bbd5;
    11'b00100110000: data <= 32'hbaf5bf10;
    11'b00100110001: data <= 32'h3c90bd97;
    11'b00100110010: data <= 32'h3eacb916;
    11'b00100110011: data <= 32'h3676b971;
    11'b00100110100: data <= 32'hba0ebc0b;
    11'b00100110101: data <= 32'hba42b1a0;
    11'b00100110110: data <= 32'hb94b3df7;
    11'b00100110111: data <= 32'hbcfe3f5e;
    11'b00100111000: data <= 32'hbee32e54;
    11'b00100111001: data <= 32'hbc87be80;
    11'b00100111010: data <= 32'haf2cbc7e;
    11'b00100111011: data <= 32'h33af3ac2;
    11'b00100111100: data <= 32'h341c3f3e;
    11'b00100111101: data <= 32'h3b633c8b;
    11'b00100111110: data <= 32'h3ef037a6;
    11'b00100111111: data <= 32'h3c9a3ae2;
    11'b00101000000: data <= 32'hb9853cc9;
    11'b00101000001: data <= 32'hbe203590;
    11'b00101000010: data <= 32'hae59bba9;
    11'b00101000011: data <= 32'h3f7cbd98;
    11'b00101000100: data <= 32'h3fedbc75;
    11'b00101000101: data <= 32'h37eebc38;
    11'b00101000110: data <= 32'hb599bc28;
    11'b00101000111: data <= 32'h31c1b144;
    11'b00101001000: data <= 32'h37683c53;
    11'b00101001001: data <= 32'hb9373ba7;
    11'b00101001010: data <= 32'hbffdba72;
    11'b00101001011: data <= 32'hbfe6c026;
    11'b00101001100: data <= 32'hbb2cbca5;
    11'b00101001101: data <= 32'hb05c39b2;
    11'b00101001110: data <= 32'h2d933cde;
    11'b00101001111: data <= 32'h38103559;
    11'b00101010000: data <= 32'h3b593070;
    11'b00101010001: data <= 32'h34973d9a;
    11'b00101010010: data <= 32'hbc6b40b6;
    11'b00101010011: data <= 32'hbda43dca;
    11'b00101010100: data <= 32'h3008b5f6;
    11'b00101010101: data <= 32'h3ef3bcd0;
    11'b00101010110: data <= 32'h3e41bac7;
    11'b00101010111: data <= 32'h3632b796;
    11'b00101011000: data <= 32'h357eb65e;
    11'b00101011001: data <= 32'h3e0b2c34;
    11'b00101011010: data <= 32'h3eee39e1;
    11'b00101011011: data <= 32'ha3a43623;
    11'b00101011100: data <= 32'hbfcabc6a;
    11'b00101011101: data <= 32'hc008c006;
    11'b00101011110: data <= 32'hb96cbcd2;
    11'b00101011111: data <= 32'h320b27af;
    11'b00101100000: data <= 32'h2c84acbb;
    11'b00101100001: data <= 32'hac1fbb5b;
    11'b00101100010: data <= 32'h2cf2b69d;
    11'b00101100011: data <= 32'hb5033e75;
    11'b00101100100: data <= 32'hbd1341a4;
    11'b00101100101: data <= 32'hbdf13eab;
    11'b00101100110: data <= 32'hb629b5f3;
    11'b00101100111: data <= 32'h398bbbe9;
    11'b00101101000: data <= 32'h381db070;
    11'b00101101001: data <= 32'h26323806;
    11'b00101101010: data <= 32'h3aca354a;
    11'b00101101011: data <= 32'h40cd346d;
    11'b00101101100: data <= 32'h40c53986;
    11'b00101101101: data <= 32'h341f38c7;
    11'b00101101110: data <= 32'hbea7b703;
    11'b00101101111: data <= 32'hbd61bd2b;
    11'b00101110000: data <= 32'h3428bc58;
    11'b00101110001: data <= 32'h3b07b9bd;
    11'b00101110010: data <= 32'h315ebd20;
    11'b00101110011: data <= 32'hb5c9bf96;
    11'b00101110100: data <= 32'hada7bad3;
    11'b00101110101: data <= 32'hac213da4;
    11'b00101110110: data <= 32'hbb2740c5;
    11'b00101110111: data <= 32'hbe573bb5;
    11'b00101111000: data <= 32'hbd15bb14;
    11'b00101111001: data <= 32'hb938bb1c;
    11'b00101111010: data <= 32'hb8cc376b;
    11'b00101111011: data <= 32'hb6f53c41;
    11'b00101111100: data <= 32'h3ace3759;
    11'b00101111101: data <= 32'h40b43103;
    11'b00101111110: data <= 32'h40253b20;
    11'b00101111111: data <= 32'h24523de4;
    11'b00110000000: data <= 32'hbd783adb;
    11'b00110000001: data <= 32'hb7feb3d3;
    11'b00110000010: data <= 32'h3c8eba22;
    11'b00110000011: data <= 32'h3d27bc0e;
    11'b00110000100: data <= 32'h312fbeb2;
    11'b00110000101: data <= 32'hb397c011;
    11'b00110000110: data <= 32'h38cdbb4c;
    11'b00110000111: data <= 32'h3c143bd6;
    11'b00110001000: data <= 32'hab543dca;
    11'b00110001001: data <= 32'hbe0eaba5;
    11'b00110001010: data <= 32'hbf9bbdb7;
    11'b00110001011: data <= 32'hbdd4bae0;
    11'b00110001100: data <= 32'hbc81389c;
    11'b00110001101: data <= 32'hb9d039d6;
    11'b00110001110: data <= 32'h364cb4a7;
    11'b00110001111: data <= 32'h3e04b696;
    11'b00110010000: data <= 32'h3c7e3c4d;
    11'b00110010001: data <= 32'hb7b940cc;
    11'b00110010010: data <= 32'hbcd03fe9;
    11'b00110010011: data <= 32'hac2b383c;
    11'b00110010100: data <= 32'h3cfeb64d;
    11'b00110010101: data <= 32'h3b7ab96c;
    11'b00110010110: data <= 32'hb0f4bc51;
    11'b00110010111: data <= 32'h2eaabd62;
    11'b00110011000: data <= 32'h3ebfb8eb;
    11'b00110011001: data <= 32'h409e38e1;
    11'b00110011010: data <= 32'h3a673997;
    11'b00110011011: data <= 32'hbcf2b8b0;
    11'b00110011100: data <= 32'hbf60bdc8;
    11'b00110011101: data <= 32'hbcf5b9c8;
    11'b00110011110: data <= 32'hba653373;
    11'b00110011111: data <= 32'hb9a8b4fb;
    11'b00110100000: data <= 32'hb22cbe3e;
    11'b00110100001: data <= 32'h3828bcd4;
    11'b00110100010: data <= 32'h35013c12;
    11'b00110100011: data <= 32'hb9f24178;
    11'b00110100100: data <= 32'hbc86406c;
    11'b00110100101: data <= 32'hb41e389d;
    11'b00110100110: data <= 32'h374db187;
    11'b00110100111: data <= 32'hafe72a30;
    11'b00110101000: data <= 32'hba312204;
    11'b00110101001: data <= 32'h34e7b6de;
    11'b00110101010: data <= 32'h40d8b4bf;
    11'b00110101011: data <= 32'h41f9373d;
    11'b00110101100: data <= 32'h3cac38f2;
    11'b00110101101: data <= 32'hbb2bb19c;
    11'b00110101110: data <= 32'hbc91b9d9;
    11'b00110101111: data <= 32'hb2d5b58a;
    11'b00110110000: data <= 32'h2a41b211;
    11'b00110110001: data <= 32'hb802bd62;
    11'b00110110010: data <= 32'hb893c128;
    11'b00110110011: data <= 32'h2da7bf29;
    11'b00110110100: data <= 32'h34e339a6;
    11'b00110110101: data <= 32'hb650407f;
    11'b00110110110: data <= 32'hbbe13dc5;
    11'b00110110111: data <= 32'hba72ab82;
    11'b00110111000: data <= 32'hb99bb178;
    11'b00110111001: data <= 32'hbd2939ad;
    11'b00110111010: data <= 32'hbdaf3a7b;
    11'b00110111011: data <= 32'h30cba9ee;
    11'b00110111100: data <= 32'h409cb5d8;
    11'b00110111101: data <= 32'h414536e2;
    11'b00110111110: data <= 32'h3ac83c9f;
    11'b00110111111: data <= 32'hb9683b57;
    11'b00111000000: data <= 32'hb40035fc;
    11'b00111000001: data <= 32'h3b01325d;
    11'b00111000010: data <= 32'h39a6b481;
    11'b00111000011: data <= 32'hb6e8be9e;
    11'b00111000100: data <= 32'hb91ec168;
    11'b00111000101: data <= 32'h3723bf46;
    11'b00111000110: data <= 32'h3cb1351d;
    11'b00111000111: data <= 32'h37e83d16;
    11'b00111001000: data <= 32'hb94e337b;
    11'b00111001001: data <= 32'hbcc4bab7;
    11'b00111001010: data <= 32'hbd9eb388;
    11'b00111001011: data <= 32'hbf563bdf;
    11'b00111001100: data <= 32'hbef43a57;
    11'b00111001101: data <= 32'hb4d7b88a;
    11'b00111001110: data <= 32'h3dabbbc4;
    11'b00111001111: data <= 32'h3e1b35a8;
    11'b00111010000: data <= 32'h301d3f3a;
    11'b00111010001: data <= 32'hb8f03fae;
    11'b00111010010: data <= 32'h35193cc4;
    11'b00111010011: data <= 32'h3d27393d;
    11'b00111010100: data <= 32'h38bf2e39;
    11'b00111010101: data <= 32'hba1ebc0f;
    11'b00111010110: data <= 32'hb874bf8b;
    11'b00111010111: data <= 32'h3cf2bd50;
    11'b00111011000: data <= 32'h40a82b5c;
    11'b00111011001: data <= 32'h3daa3693;
    11'b00111011010: data <= 32'hb3ecb8a7;
    11'b00111011011: data <= 32'hbc2bbc6e;
    11'b00111011100: data <= 32'hbc8baee1;
    11'b00111011101: data <= 32'hbda63b17;
    11'b00111011110: data <= 32'hbe422b9c;
    11'b00111011111: data <= 32'hba53bec3;
    11'b00111100000: data <= 32'h3570bf5f;
    11'b00111100001: data <= 32'h37112f4e;
    11'b00111100010: data <= 32'hb6504001;
    11'b00111100011: data <= 32'hb8a54030;
    11'b00111100100: data <= 32'h35ad3cbb;
    11'b00111100101: data <= 32'h3a7c3a2e;
    11'b00111100110: data <= 32'hb4d639f9;
    11'b00111100111: data <= 32'hbddb30f7;
    11'b00111101000: data <= 32'hb88fb9b9;
    11'b00111101001: data <= 32'h3f2fb9f2;
    11'b00111101010: data <= 32'h41e2a8bc;
    11'b00111101011: data <= 32'h3f102fe0;
    11'b00111101100: data <= 32'h29d3b7d7;
    11'b00111101101: data <= 32'hb626b89c;
    11'b00111101110: data <= 32'ha9143580;
    11'b00111101111: data <= 32'hb55f399e;
    11'b00111110000: data <= 32'hbc64ba23;
    11'b00111110001: data <= 32'hbc57c146;
    11'b00111110010: data <= 32'hb46cc0e3;
    11'b00111110011: data <= 32'h2f2eb2b2;
    11'b00111110100: data <= 32'hb40a3e19;
    11'b00111110101: data <= 32'hb6033d0b;
    11'b00111110110: data <= 32'h2b433599;
    11'b00111110111: data <= 32'haf273842;
    11'b00111111000: data <= 32'hbd903d40;
    11'b00111111001: data <= 32'hc0533c77;
    11'b00111111010: data <= 32'hba59a1a9;
    11'b00111111011: data <= 32'h3e96b8a2;
    11'b00111111100: data <= 32'h410eadee;
    11'b00111111101: data <= 32'h3d223687;
    11'b00111111110: data <= 32'h2b263582;
    11'b00111111111: data <= 32'h36a0370a;
    11'b01000000000: data <= 32'h3cc83bbc;
    11'b01000000001: data <= 32'h391a39d3;
    11'b01000000010: data <= 32'hba31bc06;
    11'b01000000011: data <= 32'hbca1c16a;
    11'b01000000100: data <= 32'hb142c0b4;
    11'b01000000101: data <= 32'h399bb6d3;
    11'b01000000110: data <= 32'h383b3904;
    11'b01000000111: data <= 32'h2900ad32;
    11'b01000001000: data <= 32'hb159b9e5;
    11'b01000001001: data <= 32'hb9b03263;
    11'b01000001010: data <= 32'hbf8d3e41;
    11'b01000001011: data <= 32'hc0d03d55;
    11'b01000001100: data <= 32'hbc81b38d;
    11'b01000001101: data <= 32'h3a8fbc35;
    11'b01000001110: data <= 32'h3d31b438;
    11'b01000001111: data <= 32'h345d3ae7;
    11'b01000010000: data <= 32'hb11a3cd7;
    11'b01000010001: data <= 32'h3b803cde;
    11'b01000010010: data <= 32'h3f523d98;
    11'b01000010011: data <= 32'h3ab03c2b;
    11'b01000010100: data <= 32'hbb91b67f;
    11'b01000010101: data <= 32'hbca1bf20;
    11'b01000010110: data <= 32'h3689be61;
    11'b01000010111: data <= 32'h3ec2b6b8;
    11'b01000011000: data <= 32'h3da4b18f;
    11'b01000011001: data <= 32'h3796bc6f;
    11'b01000011010: data <= 32'ha675bd53;
    11'b01000011011: data <= 32'hb749305c;
    11'b01000011100: data <= 32'hbd813e20;
    11'b01000011101: data <= 32'hc0003aa3;
    11'b01000011110: data <= 32'hbd74bca8;
    11'b01000011111: data <= 32'hb21dbf83;
    11'b01000100000: data <= 32'h2127b876;
    11'b01000100001: data <= 32'hb8b33c0d;
    11'b01000100010: data <= 32'hb5803d79;
    11'b01000100011: data <= 32'h3c123c8c;
    11'b01000100100: data <= 32'h3e5b3d51;
    11'b01000100101: data <= 32'h31273de3;
    11'b01000100110: data <= 32'hbe583994;
    11'b01000100111: data <= 32'hbcfeb6b5;
    11'b01000101000: data <= 32'h3b03b954;
    11'b01000101001: data <= 32'h4084b445;
    11'b01000101010: data <= 32'h3ed5b7bc;
    11'b01000101011: data <= 32'h390dbd09;
    11'b01000101100: data <= 32'h374cbc31;
    11'b01000101101: data <= 32'h38a73812;
    11'b01000101110: data <= 32'hafe93dbf;
    11'b01000101111: data <= 32'hbcc83035;
    11'b01000110000: data <= 32'hbd91c015;
    11'b01000110001: data <= 32'hba76c0e2;
    11'b01000110010: data <= 32'hb885ba5f;
    11'b01000110011: data <= 32'hb9cc394d;
    11'b01000110100: data <= 32'hb3df38a5;
    11'b01000110101: data <= 32'h3a8030b3;
    11'b01000110110: data <= 32'h3a9a3a27;
    11'b01000110111: data <= 32'hbaab3f10;
    11'b01000111000: data <= 32'hc0853e91;
    11'b01000111001: data <= 32'hbdbe3841;
    11'b01000111010: data <= 32'h3a72b22b;
    11'b01000111011: data <= 32'h3f80b1c8;
    11'b01000111100: data <= 32'h3c5cb48e;
    11'b01000111101: data <= 32'h359fb8e0;
    11'b01000111110: data <= 32'h3beeb0e0;
    11'b01000111111: data <= 32'h3f283c75;
    11'b01001000000: data <= 32'h3c613de0;
    11'b01001000001: data <= 32'hb84bb07b;
    11'b01001000010: data <= 32'hbd23c041;
    11'b01001000011: data <= 32'hba25c07b;
    11'b01001000100: data <= 32'hb1e2ba19;
    11'b01001000101: data <= 32'hae2a200f;
    11'b01001000110: data <= 32'h30beb9d7;
    11'b01001000111: data <= 32'h3909bcb8;
    11'b01001001000: data <= 32'h33972d68;
    11'b01001001001: data <= 32'hbd563f38;
    11'b01001001010: data <= 32'hc0d93fa8;
    11'b01001001011: data <= 32'hbe403843;
    11'b01001001100: data <= 32'h322eb79e;
    11'b01001001101: data <= 32'h3968b50b;
    11'b01001001110: data <= 32'hb0de2eb1;
    11'b01001001111: data <= 32'hb31b328b;
    11'b01001010000: data <= 32'h3d1e38e9;
    11'b01001010001: data <= 32'h40ed3dfb;
    11'b01001010010: data <= 32'h3e243e84;
    11'b01001010011: data <= 32'hb7ae347d;
    11'b01001010100: data <= 32'hbce3bced;
    11'b01001010101: data <= 32'hb45ebd12;
    11'b01001010110: data <= 32'h39bbb66e;
    11'b01001010111: data <= 32'h3a0bb85c;
    11'b01001011000: data <= 32'h3874bf26;
    11'b01001011001: data <= 32'h395cc010;
    11'b01001011010: data <= 32'h35a0b3e1;
    11'b01001011011: data <= 32'hbad33eb6;
    11'b01001011100: data <= 32'hbf4f3df6;
    11'b01001011101: data <= 32'hbddab461;
    11'b01001011110: data <= 32'hb888bcfc;
    11'b01001011111: data <= 32'hb913b8c8;
    11'b01001100000: data <= 32'hbd2134ee;
    11'b01001100001: data <= 32'hb9ae376d;
    11'b01001100010: data <= 32'h3ced3884;
    11'b01001100011: data <= 32'h409a3d11;
    11'b01001100100: data <= 32'h3c0c3f02;
    11'b01001100101: data <= 32'hbc233c8e;
    11'b01001100110: data <= 32'hbd3830aa;
    11'b01001100111: data <= 32'h32b5abaf;
    11'b01001101000: data <= 32'h3d632d82;
    11'b01001101001: data <= 32'h3c53b98f;
    11'b01001101010: data <= 32'h38bdc007;
    11'b01001101011: data <= 32'h3b18bfb8;
    11'b01001101100: data <= 32'h3ca31cce;
    11'b01001101101: data <= 32'h36883e47;
    11'b01001101110: data <= 32'hb9f33a75;
    11'b01001101111: data <= 32'hbc89bcb5;
    11'b01001110000: data <= 32'hbbf7bf57;
    11'b01001110001: data <= 32'hbd22ba00;
    11'b01001110010: data <= 32'hbe8a3199;
    11'b01001110011: data <= 32'hba34af83;
    11'b01001110100: data <= 32'h3bf9b6d4;
    11'b01001110101: data <= 32'h3e4c3710;
    11'b01001110110: data <= 32'h262d3eba;
    11'b01001110111: data <= 32'hbee63f7f;
    11'b01001111000: data <= 32'hbdbe3cab;
    11'b01001111001: data <= 32'h34f03948;
    11'b01001111010: data <= 32'h3c93361f;
    11'b01001111011: data <= 32'h3786b717;
    11'b01001111100: data <= 32'h2c77bdab;
    11'b01001111101: data <= 32'h3c41bc4e;
    11'b01001111110: data <= 32'h404a38e5;
    11'b01001111111: data <= 32'h3ec53e48;
    11'b01010000000: data <= 32'h320d368c;
    11'b01010000001: data <= 32'hba28bdab;
    11'b01010000010: data <= 32'hbafdbe99;
    11'b01010000011: data <= 32'hbbc0b807;
    11'b01010000100: data <= 32'hbc59b091;
    11'b01010000101: data <= 32'hb675bcd2;
    11'b01010000110: data <= 32'h3a64bf43;
    11'b01010000111: data <= 32'h3b31b849;
    11'b01010001000: data <= 32'hb8d53db0;
    11'b01010001001: data <= 32'hbfa94011;
    11'b01010001010: data <= 32'hbd8b3cfb;
    11'b01010001011: data <= 32'h1c023802;
    11'b01010001100: data <= 32'h312634e1;
    11'b01010001101: data <= 32'hbaa0a99e;
    11'b01010001110: data <= 32'hba71b86a;
    11'b01010001111: data <= 32'h3c1ab2af;
    11'b01010010000: data <= 32'h415d3c1f;
    11'b01010010001: data <= 32'h406f3e5e;
    11'b01010010010: data <= 32'h369d3874;
    11'b01010010011: data <= 32'hb8d9b9d5;
    11'b01010010100: data <= 32'hb5cab907;
    11'b01010010101: data <= 32'haa2b3105;
    11'b01010010110: data <= 32'hb14ab59b;
    11'b01010010111: data <= 32'h2a37c035;
    11'b01010011000: data <= 32'h39ebc184;
    11'b01010011001: data <= 32'h3a3abc4d;
    11'b01010011010: data <= 32'hb5273c96;
    11'b01010011011: data <= 32'hbd243e4f;
    11'b01010011100: data <= 32'hbbfe3719;
    11'b01010011101: data <= 32'hb677b4de;
    11'b01010011110: data <= 32'hbbd4a3de;
    11'b01010011111: data <= 32'hc01e333d;
    11'b01010100000: data <= 32'hbe2aae34;
    11'b01010100001: data <= 32'h3a3fac82;
    11'b01010100010: data <= 32'h40ee3a53;
    11'b01010100011: data <= 32'h3ee33dcf;
    11'b01010100100: data <= 32'hb0593c45;
    11'b01010100101: data <= 32'hb9ad3782;
    11'b01010100110: data <= 32'h3147397b;
    11'b01010100111: data <= 32'h39ed3b69;
    11'b01010101000: data <= 32'h3558b429;
    11'b01010101001: data <= 32'h2e0fc084;
    11'b01010101010: data <= 32'h39d3c16a;
    11'b01010101011: data <= 32'h3d03baff;
    11'b01010101100: data <= 32'h3a073c1f;
    11'b01010101101: data <= 32'hae493ae3;
    11'b01010101110: data <= 32'hb5d4b8ab;
    11'b01010101111: data <= 32'hb870bc31;
    11'b01010110000: data <= 32'hbe27b256;
    11'b01010110001: data <= 32'hc0f83485;
    11'b01010110010: data <= 32'hbed2b5eb;
    11'b01010110011: data <= 32'h3805baf9;
    11'b01010110100: data <= 32'h3ed6b01c;
    11'b01010110101: data <= 32'h391f3c42;
    11'b01010110110: data <= 32'hbbb03dfb;
    11'b01010110111: data <= 32'hbb133d8b;
    11'b01010111000: data <= 32'h36a93e02;
    11'b01010111001: data <= 32'h3a8a3d80;
    11'b01010111010: data <= 32'had672cec;
    11'b01010111011: data <= 32'hb806be86;
    11'b01010111100: data <= 32'h38bfbf29;
    11'b01010111101: data <= 32'h3fa9b116;
    11'b01010111110: data <= 32'h3fad3c52;
    11'b01010111111: data <= 32'h3b9e357c;
    11'b01011000000: data <= 32'h3288bc4e;
    11'b01011000001: data <= 32'hb4d1bc3a;
    11'b01011000010: data <= 32'hbcbe2e75;
    11'b01011000011: data <= 32'hbfa03428;
    11'b01011000100: data <= 32'hbd0bbc83;
    11'b01011000101: data <= 32'h3595c042;
    11'b01011000110: data <= 32'h3b83bcf1;
    11'b01011000111: data <= 32'hb2e13875;
    11'b01011001000: data <= 32'hbd613de8;
    11'b01011001001: data <= 32'hba763dab;
    11'b01011001010: data <= 32'h361b3d64;
    11'b01011001011: data <= 32'h31273d14;
    11'b01011001100: data <= 32'hbcf9372b;
    11'b01011001101: data <= 32'hbe0eb987;
    11'b01011001110: data <= 32'h345bb9c7;
    11'b01011001111: data <= 32'h4077373c;
    11'b01011010000: data <= 32'h40c63c68;
    11'b01011010001: data <= 32'h3cdf33f9;
    11'b01011010010: data <= 32'h364fb9a8;
    11'b01011010011: data <= 32'h32bdb1ed;
    11'b01011010100: data <= 32'hb2913b26;
    11'b01011010101: data <= 32'hba8335ae;
    11'b01011010110: data <= 32'hb8fdbf1b;
    11'b01011010111: data <= 32'h3505c204;
    11'b01011011000: data <= 32'h38debf68;
    11'b01011011001: data <= 32'hb3b6324d;
    11'b01011011010: data <= 32'hbb063bde;
    11'b01011011011: data <= 32'hb4cc3881;
    11'b01011011100: data <= 32'h34913682;
    11'b01011011101: data <= 32'hb9a63a45;
    11'b01011011110: data <= 32'hc0cf396c;
    11'b01011011111: data <= 32'hc0b6ab5d;
    11'b01011100000: data <= 32'haf28b49b;
    11'b01011100001: data <= 32'h3fc13640;
    11'b01011100010: data <= 32'h3f5f3ae7;
    11'b01011100011: data <= 32'h388d3734;
    11'b01011100100: data <= 32'h30fa3281;
    11'b01011100101: data <= 32'h398b3c35;
    11'b01011100110: data <= 32'h39df3f30;
    11'b01011100111: data <= 32'ha8733916;
    11'b01011101000: data <= 32'hb623bf42;
    11'b01011101001: data <= 32'h3371c1d2;
    11'b01011101010: data <= 32'h3a4abe5d;
    11'b01011101011: data <= 32'h3847319b;
    11'b01011101100: data <= 32'h332a34d9;
    11'b01011101101: data <= 32'h37ccb8be;
    11'b01011101110: data <= 32'h35e8b8c9;
    11'b01011101111: data <= 32'hbc753659;
    11'b01011110000: data <= 32'hc1933a2e;
    11'b01011110001: data <= 32'hc103aad1;
    11'b01011110010: data <= 32'hb581ba42;
    11'b01011110011: data <= 32'h3cccb6d3;
    11'b01011110100: data <= 32'h39313511;
    11'b01011110101: data <= 32'hb7e938e0;
    11'b01011110110: data <= 32'hb3363b7f;
    11'b01011110111: data <= 32'h3ba43f57;
    11'b01011111000: data <= 32'h3c42408e;
    11'b01011111001: data <= 32'hb0953bd9;
    11'b01011111010: data <= 32'hbadfbcb8;
    11'b01011111011: data <= 32'haadcbf96;
    11'b01011111100: data <= 32'h3ca1b950;
    11'b01011111101: data <= 32'h3df636c7;
    11'b01011111110: data <= 32'h3cf9b2a0;
    11'b01011111111: data <= 32'h3c88bd43;
    11'b01100000000: data <= 32'h3982bb56;
    11'b01100000001: data <= 32'hb9d33866;
    11'b01100000010: data <= 32'hc0423b10;
    11'b01100000011: data <= 32'hbf89b81b;
    11'b01100000100: data <= 32'hb510bf3a;
    11'b01100000101: data <= 32'h372fbe01;
    11'b01100000110: data <= 32'hb6adb4eb;
    11'b01100000111: data <= 32'hbcc0377f;
    11'b01100001000: data <= 32'hb5133b3d;
    11'b01100001001: data <= 32'h3c1e3e78;
    11'b01100001010: data <= 32'h39a44014;
    11'b01100001011: data <= 32'hbc333ccd;
    11'b01100001100: data <= 32'hbf51b435;
    11'b01100001101: data <= 32'hb826b915;
    11'b01100001110: data <= 32'h3d36340b;
    11'b01100001111: data <= 32'h3f763913;
    11'b01100010000: data <= 32'h3ddab626;
    11'b01100010001: data <= 32'h3cf8bcf3;
    11'b01100010010: data <= 32'h3c5cb503;
    11'b01100010011: data <= 32'h33863d28;
    11'b01100010100: data <= 32'hbae73c8c;
    11'b01100010101: data <= 32'hbb9bbb9b;
    11'b01100010110: data <= 32'hb0aec121;
    11'b01100010111: data <= 32'h2bbfc02d;
    11'b01100011000: data <= 32'hb9d0b920;
    11'b01100011001: data <= 32'hbc05284e;
    11'b01100011010: data <= 32'h2f8a2b1d;
    11'b01100011011: data <= 32'h3c623830;
    11'b01100011100: data <= 32'h2cef3d1b;
    11'b01100011101: data <= 32'hc0223ce0;
    11'b01100011110: data <= 32'hc150367d;
    11'b01100011111: data <= 32'hbb6a2cb0;
    11'b01100100000: data <= 32'h3c0e37e7;
    11'b01100100001: data <= 32'h3d3937eb;
    11'b01100100010: data <= 32'h397cb571;
    11'b01100100011: data <= 32'h3a13b8b2;
    11'b01100100100: data <= 32'h3d793a12;
    11'b01100100101: data <= 32'h3cc5405f;
    11'b01100100110: data <= 32'h31bf3df4;
    11'b01100100111: data <= 32'hb645bb87;
    11'b01100101000: data <= 32'hae41c0de;
    11'b01100101001: data <= 32'h2e1bbee4;
    11'b01100101010: data <= 32'hb339b75c;
    11'b01100101011: data <= 32'hade6b76b;
    11'b01100101100: data <= 32'h3b38bc70;
    11'b01100101101: data <= 32'h3d28b9d8;
    11'b01100101110: data <= 32'hb38e387e;
    11'b01100101111: data <= 32'hc0cd3c9c;
    11'b01100110000: data <= 32'hc1753841;
    11'b01100110001: data <= 32'hbc06b05a;
    11'b01100110010: data <= 32'h36cdaef0;
    11'b01100110011: data <= 32'h2eaea95a;
    11'b01100110100: data <= 32'hb8e4b518;
    11'b01100110101: data <= 32'h2a642107;
    11'b01100110110: data <= 32'h3dc93de8;
    11'b01100110111: data <= 32'h3e7d413d;
    11'b01100111000: data <= 32'h35c93eef;
    11'b01100111001: data <= 32'hb8fcb6b1;
    11'b01100111010: data <= 32'hb5b0bda1;
    11'b01100111011: data <= 32'h3502b8a6;
    11'b01100111100: data <= 32'h38722edb;
    11'b01100111101: data <= 32'h3ac4ba37;
    11'b01100111110: data <= 32'h3e1dbfa7;
    11'b01100111111: data <= 32'h3e42bd5e;
    11'b01101000000: data <= 32'h2d2b3715;
    11'b01101000001: data <= 32'hbee73cd4;
    11'b01101000010: data <= 32'hbfa9335a;
    11'b01101000011: data <= 32'hb970bba7;
    11'b01101000100: data <= 32'hb00abc54;
    11'b01101000101: data <= 32'hbc1eb959;
    11'b01101000110: data <= 32'hbe66b785;
    11'b01101000111: data <= 32'hb57215fe;
    11'b01101001000: data <= 32'h3dbd3cf5;
    11'b01101001001: data <= 32'h3da94071;
    11'b01101001010: data <= 32'hb50f3ebe;
    11'b01101001011: data <= 32'hbddf34ed;
    11'b01101001100: data <= 32'hbaacada8;
    11'b01101001101: data <= 32'h3669390c;
    11'b01101001110: data <= 32'h3b48391d;
    11'b01101001111: data <= 32'h3c2bbab4;
    11'b01101010000: data <= 32'h3e10bfe9;
    11'b01101010001: data <= 32'h3efabbe7;
    11'b01101010010: data <= 32'h3af73c1d;
    11'b01101010011: data <= 32'hb6893de5;
    11'b01101010100: data <= 32'hb989af65;
    11'b01101010101: data <= 32'hb183be9c;
    11'b01101010110: data <= 32'hb5f5be8e;
    11'b01101010111: data <= 32'hbde3bb5a;
    11'b01101011000: data <= 32'hbebfb9e2;
    11'b01101011001: data <= 32'hadceb99c;
    11'b01101011010: data <= 32'h3e042e8c;
    11'b01101011011: data <= 32'h3b3a3cbc;
    11'b01101011100: data <= 32'hbcf13d72;
    11'b01101011101: data <= 32'hc0843a81;
    11'b01101011110: data <= 32'hbcc839f6;
    11'b01101011111: data <= 32'h33353ca6;
    11'b01101100000: data <= 32'h376e39c4;
    11'b01101100001: data <= 32'h334cba39;
    11'b01101100010: data <= 32'h3a43bdd7;
    11'b01101100011: data <= 32'h3ec1a9d1;
    11'b01101100100: data <= 32'h3e9b3f82;
    11'b01101100101: data <= 32'h39fe3f3c;
    11'b01101100110: data <= 32'h319eb153;
    11'b01101100111: data <= 32'h3058be65;
    11'b01101101000: data <= 32'hb4bdbcf9;
    11'b01101101001: data <= 32'hbc74b82b;
    11'b01101101010: data <= 32'hbb7abb64;
    11'b01101101011: data <= 32'h3908bec1;
    11'b01101101100: data <= 32'h3ecebd08;
    11'b01101101101: data <= 32'h389b30b9;
    11'b01101101110: data <= 32'hbe743c00;
    11'b01101101111: data <= 32'hc09c3af3;
    11'b01101110000: data <= 32'hbc613979;
    11'b01101110001: data <= 32'hadc93a0a;
    11'b01101110010: data <= 32'hb88d3461;
    11'b01101110011: data <= 32'hbcabba30;
    11'b01101110100: data <= 32'hb405bb1c;
    11'b01101110101: data <= 32'h3dc7397c;
    11'b01101110110: data <= 32'h3fee4096;
    11'b01101110111: data <= 32'h3c533faa;
    11'b01101111000: data <= 32'h31913006;
    11'b01101111001: data <= 32'h18dcb9cd;
    11'b01101111010: data <= 32'hae2da1b6;
    11'b01101111011: data <= 32'hb64935d7;
    11'b01101111100: data <= 32'ha38bbb34;
    11'b01101111101: data <= 32'h3cfcc0be;
    11'b01101111110: data <= 32'h3f87c00a;
    11'b01101111111: data <= 32'h39abb384;
    11'b01110000000: data <= 32'hbc4a3b1e;
    11'b01110000001: data <= 32'hbda73896;
    11'b01110000010: data <= 32'hb774aa34;
    11'b01110000011: data <= 32'hb4dab156;
    11'b01110000100: data <= 32'hbe46b57f;
    11'b01110000101: data <= 32'hc09dbaf7;
    11'b01110000110: data <= 32'hbb7bba16;
    11'b01110000111: data <= 32'h3ce63884;
    11'b01110001000: data <= 32'h3f0d3f55;
    11'b01110001001: data <= 32'h38193e5e;
    11'b01110001010: data <= 32'hb8a83830;
    11'b01110001011: data <= 32'hb74c3740;
    11'b01110001100: data <= 32'h22ee3d69;
    11'b01110001101: data <= 32'h2a7f3cdd;
    11'b01110001110: data <= 32'h3471b9b6;
    11'b01110001111: data <= 32'h3cc3c0cd;
    11'b01110010000: data <= 32'h3f49bf2a;
    11'b01110010001: data <= 32'h3cc3332c;
    11'b01110010010: data <= 32'h2e8a3c76;
    11'b01110010011: data <= 32'ha91d3337;
    11'b01110010100: data <= 32'h3613ba54;
    11'b01110010101: data <= 32'hb449ba60;
    11'b01110010110: data <= 32'hbfd4b894;
    11'b01110010111: data <= 32'hc111bb86;
    11'b01110011000: data <= 32'hbad3bcbf;
    11'b01110011001: data <= 32'h3ce4b6ec;
    11'b01110011010: data <= 32'h3d07393a;
    11'b01110011011: data <= 32'hb6ac3b5d;
    11'b01110011100: data <= 32'hbdae39c4;
    11'b01110011101: data <= 32'hba7f3cdd;
    11'b01110011110: data <= 32'ha2504015;
    11'b01110011111: data <= 32'hb0ff3e08;
    11'b01110100000: data <= 32'hb66cb85f;
    11'b01110100001: data <= 32'h354ebf8e;
    11'b01110100010: data <= 32'h3db3baf4;
    11'b01110100011: data <= 32'h3e993c60;
    11'b01110100100: data <= 32'h3cb43dcf;
    11'b01110100101: data <= 32'h3c012c45;
    11'b01110100110: data <= 32'h3b8cbb7e;
    11'b01110100111: data <= 32'ha99fb83c;
    11'b01110101000: data <= 32'hbe65ac81;
    11'b01110101001: data <= 32'hbf54ba77;
    11'b01110101010: data <= 32'hb09bbf66;
    11'b01110101011: data <= 32'h3db1becb;
    11'b01110101100: data <= 32'h3ad9b889;
    11'b01110101101: data <= 32'hbba73435;
    11'b01110101110: data <= 32'hbe5a38af;
    11'b01110101111: data <= 32'hb9103c95;
    11'b01110110000: data <= 32'ha8f63edc;
    11'b01110110001: data <= 32'hbb003c71;
    11'b01110110010: data <= 32'hbec7b849;
    11'b01110110011: data <= 32'hbb1fbd16;
    11'b01110110100: data <= 32'h3ad4a239;
    11'b01110110101: data <= 32'h3eff3e7c;
    11'b01110110110: data <= 32'h3df33e07;
    11'b01110110111: data <= 32'h3c722ed9;
    11'b01110111000: data <= 32'h3b3fb5ba;
    11'b01110111001: data <= 32'h31d838c6;
    11'b01110111010: data <= 32'hbacf3c00;
    11'b01110111011: data <= 32'hba90b704;
    11'b01110111100: data <= 32'h3898c08a;
    11'b01110111101: data <= 32'h3e4fc0db;
    11'b01110111110: data <= 32'h3a36bc5d;
    11'b01110111111: data <= 32'hb9811c4a;
    11'b01111000000: data <= 32'hba71336d;
    11'b01111000001: data <= 32'h316f3663;
    11'b01111000010: data <= 32'h2e5939e5;
    11'b01111000011: data <= 32'hbe5e368c;
    11'b01111000100: data <= 32'hc196b905;
    11'b01111000101: data <= 32'hbef9bbc6;
    11'b01111000110: data <= 32'h36ed2f60;
    11'b01111000111: data <= 32'h3dbb3d1c;
    11'b01111001000: data <= 32'h3b453c1d;
    11'b01111001001: data <= 32'h35613124;
    11'b01111001010: data <= 32'h363d3839;
    11'b01111001011: data <= 32'h34943fa9;
    11'b01111001100: data <= 32'hb45f4015;
    11'b01111001101: data <= 32'hb4e09bd4;
    11'b01111001110: data <= 32'h3925c053;
    11'b01111001111: data <= 32'h3d8fc061;
    11'b01111010000: data <= 32'h3b76b936;
    11'b01111010001: data <= 32'h321f33fc;
    11'b01111010010: data <= 32'h3824af0d;
    11'b01111010011: data <= 32'h3ce5b720;
    11'b01111010100: data <= 32'h36c6ada4;
    11'b01111010101: data <= 32'hbf3c2a69;
    11'b01111010110: data <= 32'hc207b8d5;
    11'b01111010111: data <= 32'hbee0bc64;
    11'b01111011000: data <= 32'h367db8b5;
    11'b01111011001: data <= 32'h3b5a3100;
    11'b01111011010: data <= 32'hae473081;
    11'b01111011011: data <= 32'hb95528e4;
    11'b01111011100: data <= 32'hae2a3c5a;
    11'b01111011101: data <= 32'h35214132;
    11'b01111011110: data <= 32'hb2e340de;
    11'b01111011111: data <= 32'hb99533a8;
    11'b01111100000: data <= 32'hb09abe7c;
    11'b01111100001: data <= 32'h3a3fbcd5;
    11'b01111100010: data <= 32'h3c3435a0;
    11'b01111100011: data <= 32'h3c2739ab;
    11'b01111100100: data <= 32'h3e3ab4d8;
    11'b01111100101: data <= 32'h3fb7ba90;
    11'b01111100110: data <= 32'h3a37ae19;
    11'b01111100111: data <= 32'hbd933769;
    11'b01111101000: data <= 32'hc088b46d;
    11'b01111101001: data <= 32'hbb4abda9;
    11'b01111101010: data <= 32'h39b0be6e;
    11'b01111101011: data <= 32'h3801bc41;
    11'b01111101100: data <= 32'hbaaeb992;
    11'b01111101101: data <= 32'hbc61b47f;
    11'b01111101110: data <= 32'ha5d63b76;
    11'b01111101111: data <= 32'h3769407c;
    11'b01111110000: data <= 32'hb8c43fe9;
    11'b01111110001: data <= 32'hbeee317a;
    11'b01111110010: data <= 32'hbd72bbf5;
    11'b01111110011: data <= 32'h0e24b1d1;
    11'b01111110100: data <= 32'h3b553c80;
    11'b01111110101: data <= 32'h3cef3b14;
    11'b01111110110: data <= 32'h3e9eb66c;
    11'b01111110111: data <= 32'h3f86b882;
    11'b01111111000: data <= 32'h3bb23a1f;
    11'b01111111001: data <= 32'hb9173e15;
    11'b01111111010: data <= 32'hbc703519;
    11'b01111111011: data <= 32'h28adbe3e;
    11'b01111111100: data <= 32'h3bfec063;
    11'b01111111101: data <= 32'h3503be5c;
    11'b01111111110: data <= 32'hbaf2bbfa;
    11'b01111111111: data <= 32'hb8a7b921;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    