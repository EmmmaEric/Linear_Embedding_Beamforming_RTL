
module memory_rom_23(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3e28b615;
    11'b00000000001: data <= 32'h3a9cb3fd;
    11'b00000000010: data <= 32'hbb9b31d2;
    11'b00000000011: data <= 32'hbf44b766;
    11'b00000000100: data <= 32'hb808bea0;
    11'b00000000101: data <= 32'h3d87bfa9;
    11'b00000000110: data <= 32'h3d9fbc97;
    11'b00000000111: data <= 32'hb495b7b3;
    11'b00000001000: data <= 32'hbd60b1a8;
    11'b00000001001: data <= 32'hba123862;
    11'b00000001010: data <= 32'haf6a3e35;
    11'b00000001011: data <= 32'hbab23dab;
    11'b00000001100: data <= 32'hbfafb28b;
    11'b00000001101: data <= 32'hbe73bdae;
    11'b00000001110: data <= 32'hae0db867;
    11'b00000001111: data <= 32'h3c0d3d3c;
    11'b00000010000: data <= 32'h3c983f11;
    11'b00000010001: data <= 32'h3c8838df;
    11'b00000010010: data <= 32'h3ce2ac4f;
    11'b00000010011: data <= 32'h38f63a3e;
    11'b00000010100: data <= 32'hb90c3e1d;
    11'b00000010101: data <= 32'hbc0037b9;
    11'b00000010110: data <= 32'h34ebbdf4;
    11'b00000010111: data <= 32'h3eeec08a;
    11'b00000011000: data <= 32'h3d9abdf8;
    11'b00000011001: data <= 32'had0cb88c;
    11'b00000011010: data <= 32'hb83fb41b;
    11'b00000011011: data <= 32'h363e2ca5;
    11'b00000011100: data <= 32'h3936390b;
    11'b00000011101: data <= 32'hbb613799;
    11'b00000011110: data <= 32'hc14fb96f;
    11'b00000011111: data <= 32'hc0c7bd9a;
    11'b00000100000: data <= 32'hb843b82e;
    11'b00000100001: data <= 32'h39ff3af8;
    11'b00000100010: data <= 32'h392b3bbe;
    11'b00000100011: data <= 32'h343d2ded;
    11'b00000100100: data <= 32'h357033fd;
    11'b00000100101: data <= 32'h32d73f4b;
    11'b00000100110: data <= 32'hb754414f;
    11'b00000100111: data <= 32'hb9483ca8;
    11'b00000101000: data <= 32'h34ddbcc7;
    11'b00000101001: data <= 32'h3d5ebfb1;
    11'b00000101010: data <= 32'h3c95bad0;
    11'b00000101011: data <= 32'h36162e33;
    11'b00000101100: data <= 32'h393eaa9f;
    11'b00000101101: data <= 32'h3ec9b581;
    11'b00000101110: data <= 32'h3dbda94f;
    11'b00000101111: data <= 32'hb9f02d56;
    11'b00000110000: data <= 32'hc143b919;
    11'b00000110001: data <= 32'hc046bd57;
    11'b00000110010: data <= 32'hb1f4bbfc;
    11'b00000110011: data <= 32'h39b8b426;
    11'b00000110100: data <= 32'h9d56b4d1;
    11'b00000110101: data <= 32'hb97eb90b;
    11'b00000110110: data <= 32'hb5723487;
    11'b00000110111: data <= 32'h2a6c406b;
    11'b00000111000: data <= 32'hb6ec41c2;
    11'b00000111001: data <= 32'hbc023cb9;
    11'b00000111010: data <= 32'hb8c9bbb9;
    11'b00000111011: data <= 32'h34bfbc9d;
    11'b00000111100: data <= 32'h38fe33a8;
    11'b00000111101: data <= 32'h39673b5b;
    11'b00000111110: data <= 32'h3dba30ed;
    11'b00000111111: data <= 32'h40bdb802;
    11'b00001000000: data <= 32'h3f1e2407;
    11'b00001000001: data <= 32'hb69d3919;
    11'b00001000010: data <= 32'hbfae2d87;
    11'b00001000011: data <= 32'hbc73bc4f;
    11'b00001000100: data <= 32'h38d7be2d;
    11'b00001000101: data <= 32'h3aa3bd52;
    11'b00001000110: data <= 32'hb6a1bd26;
    11'b00001000111: data <= 32'hbc16bcb8;
    11'b00001001000: data <= 32'hb24ca592;
    11'b00001001001: data <= 32'h373b3ee7;
    11'b00001001010: data <= 32'hb6454043;
    11'b00001001011: data <= 32'hbed538c2;
    11'b00001001100: data <= 32'hbf47bb38;
    11'b00001001101: data <= 32'hba88b77f;
    11'b00001001110: data <= 32'h2a9a3bcc;
    11'b00001001111: data <= 32'h384b3cb4;
    11'b00001010000: data <= 32'h3d331f0b;
    11'b00001010001: data <= 32'h4010b75d;
    11'b00001010010: data <= 32'h3e1139b4;
    11'b00001010011: data <= 32'hb0623f57;
    11'b00001010100: data <= 32'hbc193c9b;
    11'b00001010101: data <= 32'had8fb92d;
    11'b00001010110: data <= 32'h3ca5bec9;
    11'b00001010111: data <= 32'h3aa2be77;
    11'b00001011000: data <= 32'hb736bd91;
    11'b00001011001: data <= 32'hb845bd04;
    11'b00001011010: data <= 32'h3a57b7a4;
    11'b00001011011: data <= 32'h3d5a39ec;
    11'b00001011100: data <= 32'hb2103c01;
    11'b00001011101: data <= 32'hc068ad22;
    11'b00001011110: data <= 32'hc10dbb49;
    11'b00001011111: data <= 32'hbd3ab343;
    11'b00001100000: data <= 32'hb4393ad1;
    11'b00001100001: data <= 32'h24e63861;
    11'b00001100010: data <= 32'h3608b8f4;
    11'b00001100011: data <= 32'h3bf4b71a;
    11'b00001100100: data <= 32'h3b643df5;
    11'b00001100101: data <= 32'ha1be41c4;
    11'b00001100110: data <= 32'hb8013fab;
    11'b00001100111: data <= 32'h32d9b3cd;
    11'b00001101000: data <= 32'h3ba3bd2b;
    11'b00001101001: data <= 32'h37b6bb67;
    11'b00001101010: data <= 32'hb4b3b8d7;
    11'b00001101011: data <= 32'h35e0bb1b;
    11'b00001101100: data <= 32'h4007bab4;
    11'b00001101101: data <= 32'h4077ad93;
    11'b00001101110: data <= 32'h30e7351a;
    11'b00001101111: data <= 32'hc029b3a8;
    11'b00001110000: data <= 32'hc073ba3a;
    11'b00001110001: data <= 32'hbb05b686;
    11'b00001110010: data <= 32'hb19e250f;
    11'b00001110011: data <= 32'hb8a4b906;
    11'b00001110100: data <= 32'hb9a6bde6;
    11'b00001110101: data <= 32'h291eb8f5;
    11'b00001110110: data <= 32'h385e3ef4;
    11'b00001110111: data <= 32'h2a67421f;
    11'b00001111000: data <= 32'hb8853f92;
    11'b00001111001: data <= 32'hb618add1;
    11'b00001111010: data <= 32'h242ab877;
    11'b00001111011: data <= 32'hb1de3477;
    11'b00001111100: data <= 32'hb3dc3786;
    11'b00001111101: data <= 32'h3bcab766;
    11'b00001111110: data <= 32'h4149bc01;
    11'b00001111111: data <= 32'h4129b491;
    11'b00010000000: data <= 32'h3758387a;
    11'b00010000001: data <= 32'hbd8535ba;
    11'b00010000010: data <= 32'hbc67b612;
    11'b00010000011: data <= 32'h3084b970;
    11'b00010000100: data <= 32'h30f7bacf;
    11'b00010000101: data <= 32'hbbc9be4c;
    11'b00010000110: data <= 32'hbd18c025;
    11'b00010000111: data <= 32'hb034bbaa;
    11'b00010001000: data <= 32'h3a613cf3;
    11'b00010001001: data <= 32'h32fa4073;
    11'b00010001010: data <= 32'hbbdd3c70;
    11'b00010001011: data <= 32'hbd81b354;
    11'b00010001100: data <= 32'hbc3a2e35;
    11'b00010001101: data <= 32'hbac53ce7;
    11'b00010001110: data <= 32'hb79a3c2a;
    11'b00010001111: data <= 32'h3a5bb6f8;
    11'b00010010000: data <= 32'h4077bc42;
    11'b00010010001: data <= 32'h40522fbf;
    11'b00010010010: data <= 32'h387a3e0a;
    11'b00010010011: data <= 32'hb8273d82;
    11'b00010010100: data <= 32'h2f8d318e;
    11'b00010010101: data <= 32'h3c09b980;
    11'b00010010110: data <= 32'h3598bc3c;
    11'b00010010111: data <= 32'hbc59be7f;
    11'b00010011000: data <= 32'hbc49c012;
    11'b00010011001: data <= 32'h38bdbd19;
    11'b00010011010: data <= 32'h3e80348a;
    11'b00010011011: data <= 32'h387f3b59;
    11'b00010011100: data <= 32'hbd273026;
    11'b00010011101: data <= 32'hbfe6b735;
    11'b00010011110: data <= 32'hbe083641;
    11'b00010011111: data <= 32'hbc6b3d86;
    11'b00010100000: data <= 32'hbb37398e;
    11'b00010100001: data <= 32'haeecbbe0;
    11'b00010100010: data <= 32'h3c27bcca;
    11'b00010100011: data <= 32'h3d1b3968;
    11'b00010100100: data <= 32'h376540d8;
    11'b00010100101: data <= 32'h2851403c;
    11'b00010100110: data <= 32'h39823895;
    11'b00010100111: data <= 32'h3c68b51f;
    11'b00010101000: data <= 32'h2ea4b5f1;
    11'b00010101001: data <= 32'hbc4db99d;
    11'b00010101010: data <= 32'hb6a2bda0;
    11'b00010101011: data <= 32'h3e9ebda7;
    11'b00010101100: data <= 32'h4101b86e;
    11'b00010101101: data <= 32'h3b98a645;
    11'b00010101110: data <= 32'hbc97b588;
    11'b00010101111: data <= 32'hbe9fb72d;
    11'b00010110000: data <= 32'hbbbc3581;
    11'b00010110001: data <= 32'hba523a7a;
    11'b00010110010: data <= 32'hbd2eb4cd;
    11'b00010110011: data <= 32'hbcc2bf4f;
    11'b00010110100: data <= 32'hb142bdd4;
    11'b00010110101: data <= 32'h388c3ad9;
    11'b00010110110: data <= 32'h35c8411f;
    11'b00010110111: data <= 32'h2d754002;
    11'b00010111000: data <= 32'h35de385e;
    11'b00010111001: data <= 32'h35e83392;
    11'b00010111010: data <= 32'hb85d3a9f;
    11'b00010111011: data <= 32'hbc9338dc;
    11'b00010111100: data <= 32'h2d13b929;
    11'b00010111101: data <= 32'h4074bd8c;
    11'b00010111110: data <= 32'h4194bac4;
    11'b00010111111: data <= 32'h3c82ac23;
    11'b00011000000: data <= 32'hb8b22449;
    11'b00011000001: data <= 32'hb845ad1a;
    11'b00011000010: data <= 32'h344d32ad;
    11'b00011000011: data <= 32'hb0262dc1;
    11'b00011000100: data <= 32'hbdebbcb2;
    11'b00011000101: data <= 32'hbf50c0c8;
    11'b00011000110: data <= 32'hb8f8bee3;
    11'b00011000111: data <= 32'h3871373b;
    11'b00011001000: data <= 32'h37963ee3;
    11'b00011001001: data <= 32'hb1ff3c1a;
    11'b00011001010: data <= 32'hb7182e0f;
    11'b00011001011: data <= 32'hb8e5396c;
    11'b00011001100: data <= 32'hbccb3f52;
    11'b00011001101: data <= 32'hbd693ddd;
    11'b00011001110: data <= 32'haa26b532;
    11'b00011001111: data <= 32'h3f3cbd74;
    11'b00011010000: data <= 32'h4066b8a8;
    11'b00011010001: data <= 32'h3b883962;
    11'b00011010010: data <= 32'h2c303b5d;
    11'b00011010011: data <= 32'h39da37a5;
    11'b00011010100: data <= 32'h3db23364;
    11'b00011010101: data <= 32'h3620affe;
    11'b00011010110: data <= 32'hbde6bcd6;
    11'b00011010111: data <= 32'hbf0ac070;
    11'b00011011000: data <= 32'hb039bf2a;
    11'b00011011001: data <= 32'h3cf5b4ed;
    11'b00011011010: data <= 32'h3a9b3603;
    11'b00011011011: data <= 32'hb6c4b3af;
    11'b00011011100: data <= 32'hbc06b76a;
    11'b00011011101: data <= 32'hbc2c3a98;
    11'b00011011110: data <= 32'hbd6f4037;
    11'b00011011111: data <= 32'hbe533d7e;
    11'b00011100000: data <= 32'hba3db996;
    11'b00011100001: data <= 32'h38a4bdfa;
    11'b00011100010: data <= 32'h3c28b002;
    11'b00011100011: data <= 32'h37f33e0a;
    11'b00011100100: data <= 32'h372b3e86;
    11'b00011100101: data <= 32'h3da83a87;
    11'b00011100110: data <= 32'h3f2a3747;
    11'b00011100111: data <= 32'h358e36c5;
    11'b00011101000: data <= 32'hbdc7b424;
    11'b00011101001: data <= 32'hbce0bd54;
    11'b00011101010: data <= 32'h3a90be56;
    11'b00011101011: data <= 32'h4027bbac;
    11'b00011101100: data <= 32'h3cbbb95f;
    11'b00011101101: data <= 32'hb5efbc0a;
    11'b00011101110: data <= 32'hba52b9ad;
    11'b00011101111: data <= 32'hb7ae39e1;
    11'b00011110000: data <= 32'hba873ea6;
    11'b00011110001: data <= 32'hbe973829;
    11'b00011110010: data <= 32'hbeacbdf0;
    11'b00011110011: data <= 32'hb9bfbefe;
    11'b00011110100: data <= 32'h25752e0a;
    11'b00011110101: data <= 32'h2f113ede;
    11'b00011110110: data <= 32'h36db3e02;
    11'b00011110111: data <= 32'h3ce738c8;
    11'b00011111000: data <= 32'h3cee39ba;
    11'b00011111001: data <= 32'hb3233dbc;
    11'b00011111010: data <= 32'hbe143c8d;
    11'b00011111011: data <= 32'hb9d1b40a;
    11'b00011111100: data <= 32'h3db6bcf6;
    11'b00011111101: data <= 32'h40b4bc9a;
    11'b00011111110: data <= 32'h3cd5bac8;
    11'b00011111111: data <= 32'hac1fbad7;
    11'b00100000000: data <= 32'h3106b738;
    11'b00100000001: data <= 32'h3aad38e3;
    11'b00100000010: data <= 32'h31253bd8;
    11'b00100000011: data <= 32'hbdf9b5b4;
    11'b00100000100: data <= 32'hc05cc015;
    11'b00100000101: data <= 32'hbd3fbf9b;
    11'b00100000110: data <= 32'hb388ae6d;
    11'b00100000111: data <= 32'h2ca93c21;
    11'b00100001000: data <= 32'h311e3741;
    11'b00100001001: data <= 32'h37b8b111;
    11'b00100001010: data <= 32'h347b3a7d;
    11'b00100001011: data <= 32'hbaf84095;
    11'b00100001100: data <= 32'hbea24043;
    11'b00100001101: data <= 32'hb989357f;
    11'b00100001110: data <= 32'h3c94bc16;
    11'b00100001111: data <= 32'h3ed1bafc;
    11'b00100010000: data <= 32'h39ebb267;
    11'b00100010001: data <= 32'h33eea431;
    11'b00100010010: data <= 32'h3d122e21;
    11'b00100010011: data <= 32'h404038c6;
    11'b00100010100: data <= 32'h3bd03933;
    11'b00100010101: data <= 32'hbd01b80e;
    11'b00100010110: data <= 32'hc026bf52;
    11'b00100010111: data <= 32'hbb71bee0;
    11'b00100011000: data <= 32'h3584b84b;
    11'b00100011001: data <= 32'h3654b107;
    11'b00100011010: data <= 32'had9cbb96;
    11'b00100011011: data <= 32'hb0dabc2a;
    11'b00100011100: data <= 32'hb3d53977;
    11'b00100011101: data <= 32'hbc0c4104;
    11'b00100011110: data <= 32'hbeb44053;
    11'b00100011111: data <= 32'hbc812f55;
    11'b00100100000: data <= 32'h2c87bc62;
    11'b00100100001: data <= 32'h369ab6a7;
    11'b00100100010: data <= 32'ha96f395b;
    11'b00100100011: data <= 32'h35393a1c;
    11'b00100100100: data <= 32'h3f7e36e6;
    11'b00100100101: data <= 32'h4143393d;
    11'b00100100110: data <= 32'h3c833b7d;
    11'b00100100111: data <= 32'hbc8234a9;
    11'b00100101000: data <= 32'hbe22ba96;
    11'b00100101001: data <= 32'h258dbcb1;
    11'b00100101010: data <= 32'h3ce4baea;
    11'b00100101011: data <= 32'h3a15bc71;
    11'b00100101100: data <= 32'hb10fbf7b;
    11'b00100101101: data <= 32'hb112be13;
    11'b00100101110: data <= 32'h3189375b;
    11'b00100101111: data <= 32'hb5e8401e;
    11'b00100110000: data <= 32'hbda93d59;
    11'b00100110001: data <= 32'hbebbb975;
    11'b00100110010: data <= 32'hbc7dbd6f;
    11'b00100110011: data <= 32'hba2caf12;
    11'b00100110100: data <= 32'hb99f3c3c;
    11'b00100110101: data <= 32'h302a3a2d;
    11'b00100110110: data <= 32'h3ead3062;
    11'b00100110111: data <= 32'h404238f0;
    11'b00100111000: data <= 32'h38aa3e7a;
    11'b00100111001: data <= 32'hbcd13e4a;
    11'b00100111010: data <= 32'hbbe136df;
    11'b00100111011: data <= 32'h3a35b826;
    11'b00100111100: data <= 32'h3e81bab1;
    11'b00100111101: data <= 32'h39e3bd0b;
    11'b00100111110: data <= 32'haf56bf37;
    11'b00100111111: data <= 32'h37a2bd50;
    11'b00101000000: data <= 32'h3d773521;
    11'b00101000001: data <= 32'h3a3e3d5b;
    11'b00101000010: data <= 32'hbb693590;
    11'b00101000011: data <= 32'hbfc1bd6d;
    11'b00101000100: data <= 32'hbeb5bdf2;
    11'b00101000101: data <= 32'hbc96ad31;
    11'b00101000110: data <= 32'hbae0394f;
    11'b00101000111: data <= 32'hb1d2b0e6;
    11'b00101001000: data <= 32'h3b38ba43;
    11'b00101001001: data <= 32'h3c6335dd;
    11'b00101001010: data <= 32'hb15c4063;
    11'b00101001011: data <= 32'hbd5b4109;
    11'b00101001100: data <= 32'hba1e3cb0;
    11'b00101001101: data <= 32'h3a0fb015;
    11'b00101001110: data <= 32'h3c6db7a7;
    11'b00101001111: data <= 32'h2fa6b8c7;
    11'b00101010000: data <= 32'hb0a6bb5e;
    11'b00101010001: data <= 32'h3d29b99e;
    11'b00101010010: data <= 32'h41333512;
    11'b00101010011: data <= 32'h3f113ae3;
    11'b00101010100: data <= 32'hb75da988;
    11'b00101010101: data <= 32'hbed8bd1d;
    11'b00101010110: data <= 32'hbd1fbcb7;
    11'b00101010111: data <= 32'hb87cb208;
    11'b00101011000: data <= 32'hb7dbb324;
    11'b00101011001: data <= 32'hb6a5bdf6;
    11'b00101011010: data <= 32'h30edbf6b;
    11'b00101011011: data <= 32'h35baa78e;
    11'b00101011100: data <= 32'hb7304080;
    11'b00101011101: data <= 32'hbd0b4110;
    11'b00101011110: data <= 32'hbb253bcf;
    11'b00101011111: data <= 32'ha376b281;
    11'b00101100000: data <= 32'haf52a682;
    11'b00101100001: data <= 32'hbae835c3;
    11'b00101100010: data <= 32'hb5eb29b4;
    11'b00101100011: data <= 32'h3eccb31c;
    11'b00101100100: data <= 32'h422d3502;
    11'b00101100101: data <= 32'h3ff63af8;
    11'b00101100110: data <= 32'hb49d3755;
    11'b00101100111: data <= 32'hbc9db5a8;
    11'b00101101000: data <= 32'hb42ab6eb;
    11'b00101101001: data <= 32'h378db206;
    11'b00101101010: data <= 32'h22dbbba1;
    11'b00101101011: data <= 32'hb825c0cb;
    11'b00101101100: data <= 32'hae05c0e3;
    11'b00101101101: data <= 32'h37ceb5ab;
    11'b00101101110: data <= 32'h2e2c3f05;
    11'b00101101111: data <= 32'hba7d3e9c;
    11'b00101110000: data <= 32'hbc702b75;
    11'b00101110001: data <= 32'hbbb3b8ba;
    11'b00101110010: data <= 32'hbd2434ab;
    11'b00101110011: data <= 32'hbeb43ba6;
    11'b00101110100: data <= 32'hb9c6353e;
    11'b00101110101: data <= 32'h3dafb66e;
    11'b00101110110: data <= 32'h41172ef0;
    11'b00101110111: data <= 32'h3d723cdc;
    11'b00101111000: data <= 32'hb7753dea;
    11'b00101111001: data <= 32'hb8d23b12;
    11'b00101111010: data <= 32'h39603687;
    11'b00101111011: data <= 32'h3c8a2a27;
    11'b00101111100: data <= 32'h2fa8bbfc;
    11'b00101111101: data <= 32'hb8e5c09b;
    11'b00101111110: data <= 32'h32e7c06e;
    11'b00101111111: data <= 32'h3da4b6d4;
    11'b00110000000: data <= 32'h3ce43c23;
    11'b00110000001: data <= 32'haf4b3812;
    11'b00110000010: data <= 32'hbc72bae1;
    11'b00110000011: data <= 32'hbd86bae6;
    11'b00110000100: data <= 32'hbe9836d8;
    11'b00110000101: data <= 32'hbf5f3af1;
    11'b00110000110: data <= 32'hbc0bb520;
    11'b00110000111: data <= 32'h392abd24;
    11'b00110001000: data <= 32'h3d87b5be;
    11'b00110001001: data <= 32'h36303e02;
    11'b00110001010: data <= 32'hba044085;
    11'b00110001011: data <= 32'hb4de3e82;
    11'b00110001100: data <= 32'h3b813ae5;
    11'b00110001101: data <= 32'h3b2b36fc;
    11'b00110001110: data <= 32'hb719b4f8;
    11'b00110001111: data <= 32'hbad9bd41;
    11'b00110010000: data <= 32'h39c5bd90;
    11'b00110010001: data <= 32'h40eab477;
    11'b00110010010: data <= 32'h40703804;
    11'b00110010011: data <= 32'h376eb0a8;
    11'b00110010100: data <= 32'hba5fbc44;
    11'b00110010101: data <= 32'hbb86b90a;
    11'b00110010110: data <= 32'hbbd53829;
    11'b00110010111: data <= 32'hbd4234c6;
    11'b00110011000: data <= 32'hbc6cbdd1;
    11'b00110011001: data <= 32'hb066c0bf;
    11'b00110011010: data <= 32'h3669bb46;
    11'b00110011011: data <= 32'hb1d53dac;
    11'b00110011100: data <= 32'hba324069;
    11'b00110011101: data <= 32'hb40d3d7d;
    11'b00110011110: data <= 32'h37c93963;
    11'b00110011111: data <= 32'haecf3a37;
    11'b00110100000: data <= 32'hbdc7395f;
    11'b00110100001: data <= 32'hbd11b021;
    11'b00110100010: data <= 32'h3b8eb901;
    11'b00110100011: data <= 32'h41b6b10f;
    11'b00110100100: data <= 32'h40d135be;
    11'b00110100101: data <= 32'h389b28d8;
    11'b00110100110: data <= 32'hb504b606;
    11'b00110100111: data <= 32'h2ea4301b;
    11'b00110101000: data <= 32'h33fa39d6;
    11'b00110101001: data <= 32'hb847b2a9;
    11'b00110101010: data <= 32'hbc42c082;
    11'b00110101011: data <= 32'hb815c1e9;
    11'b00110101100: data <= 32'h3304bce9;
    11'b00110101101: data <= 32'h2f003b9e;
    11'b00110101110: data <= 32'hb5473d2f;
    11'b00110101111: data <= 32'hb400348b;
    11'b00110110000: data <= 32'hb2a127c2;
    11'b00110110001: data <= 32'hbc9e3b88;
    11'b00110110010: data <= 32'hc08b3d78;
    11'b00110110011: data <= 32'hbeac3749;
    11'b00110110100: data <= 32'h392db843;
    11'b00110110101: data <= 32'h408cb54d;
    11'b00110110110: data <= 32'h3e8c37c9;
    11'b00110110111: data <= 32'h31873a3f;
    11'b00110111000: data <= 32'h2db039c3;
    11'b00110111001: data <= 32'h3c783c04;
    11'b00110111010: data <= 32'h3cce3c45;
    11'b00110111011: data <= 32'hb082b1f9;
    11'b00110111100: data <= 32'hbc63c03a;
    11'b00110111101: data <= 32'hb678c13a;
    11'b00110111110: data <= 32'h3ac9bc75;
    11'b00110111111: data <= 32'h3c4c35d7;
    11'b00111000000: data <= 32'h36982d56;
    11'b00111000001: data <= 32'haec8bb49;
    11'b00111000010: data <= 32'hb81db84e;
    11'b00111000011: data <= 32'hbdda3be7;
    11'b00111000100: data <= 32'hc0ba3dda;
    11'b00111000101: data <= 32'hbf492f0a;
    11'b00111000110: data <= 32'ha503bcee;
    11'b00111000111: data <= 32'h3c31baba;
    11'b00111001000: data <= 32'h366638c1;
    11'b00111001001: data <= 32'hb6a13da2;
    11'b00111001010: data <= 32'h34643d9b;
    11'b00111001011: data <= 32'h3e323daf;
    11'b00111001100: data <= 32'h3d163d81;
    11'b00111001101: data <= 32'hb7ed36cb;
    11'b00111001110: data <= 32'hbd7bbc44;
    11'b00111001111: data <= 32'hae34be32;
    11'b00111010000: data <= 32'h3ed5b95f;
    11'b00111010001: data <= 32'h3ffea8d7;
    11'b00111010010: data <= 32'h3beab9c4;
    11'b00111010011: data <= 32'h3208bdbb;
    11'b00111010100: data <= 32'haf14b854;
    11'b00111010101: data <= 32'hb9ef3c5b;
    11'b00111010110: data <= 32'hbe7f3c66;
    11'b00111010111: data <= 32'hbe8dba77;
    11'b00111011000: data <= 32'hb953c078;
    11'b00111011001: data <= 32'hac5cbdac;
    11'b00111011010: data <= 32'hb7d63798;
    11'b00111011011: data <= 32'hb9983d66;
    11'b00111011100: data <= 32'h34f33c65;
    11'b00111011101: data <= 32'h3d383c3c;
    11'b00111011110: data <= 32'h38113de2;
    11'b00111011111: data <= 32'hbd943d17;
    11'b00111100000: data <= 32'hbf4f33ac;
    11'b00111100001: data <= 32'h2972b762;
    11'b00111100010: data <= 32'h401fb432;
    11'b00111100011: data <= 32'h4049b060;
    11'b00111100100: data <= 32'h3bc2b9ee;
    11'b00111100101: data <= 32'h378bbc05;
    11'b00111100110: data <= 32'h3a832e03;
    11'b00111100111: data <= 32'h38c43d6a;
    11'b00111101000: data <= 32'hb83e39b9;
    11'b00111101001: data <= 32'hbd29be1e;
    11'b00111101010: data <= 32'hbbbbc18c;
    11'b00111101011: data <= 32'hb726be99;
    11'b00111101100: data <= 32'hb7be3105;
    11'b00111101101: data <= 32'hb682384c;
    11'b00111101110: data <= 32'h35dcadad;
    11'b00111101111: data <= 32'h3a1b2f97;
    11'b00111110000: data <= 32'hb6de3d4c;
    11'b00111110001: data <= 32'hc05d3f7f;
    11'b00111110010: data <= 32'hc05e3c0d;
    11'b00111110011: data <= 32'hb11dabc0;
    11'b00111110100: data <= 32'h3e32b3f3;
    11'b00111110101: data <= 32'h3d21aa70;
    11'b00111110110: data <= 32'h34b6b187;
    11'b00111110111: data <= 32'h3893aa46;
    11'b00111111000: data <= 32'h3ee23b6e;
    11'b00111111001: data <= 32'h3ee93ebf;
    11'b00111111010: data <= 32'h3211398f;
    11'b00111111011: data <= 32'hbc65bdb9;
    11'b00111111100: data <= 32'hbb0ac0b6;
    11'b00111111101: data <= 32'h9ee6bd31;
    11'b00111111110: data <= 32'h34edb0ca;
    11'b00111111111: data <= 32'h3490b889;
    11'b01000000000: data <= 32'h384dbdd2;
    11'b01000000001: data <= 32'h376bba4f;
    11'b01000000010: data <= 32'hba083c75;
    11'b01000000011: data <= 32'hc06f3fdb;
    11'b01000000100: data <= 32'hc0473aea;
    11'b01000000101: data <= 32'hb89eb86e;
    11'b01000000110: data <= 32'h36d9b980;
    11'b01000000111: data <= 32'haf9f2152;
    11'b01000001000: data <= 32'hb919366f;
    11'b01000001001: data <= 32'h379b38f8;
    11'b01000001010: data <= 32'h403f3d3a;
    11'b01000001011: data <= 32'h40003f63;
    11'b01000001100: data <= 32'h2cc53c63;
    11'b01000001101: data <= 32'hbd18b7ad;
    11'b01000001110: data <= 32'hb902bc8e;
    11'b01000001111: data <= 32'h3a1ab819;
    11'b01000010000: data <= 32'h3cc5b412;
    11'b01000010001: data <= 32'h3ab3bd4c;
    11'b01000010010: data <= 32'h39dfc05f;
    11'b01000010011: data <= 32'h39a4bc41;
    11'b01000010100: data <= 32'haf7e3c54;
    11'b01000010101: data <= 32'hbd5d3e9a;
    11'b01000010110: data <= 32'hbe852c29;
    11'b01000010111: data <= 32'hbb5cbdf3;
    11'b01000011000: data <= 32'hb907bcfc;
    11'b01000011001: data <= 32'hbce4ab4b;
    11'b01000011010: data <= 32'hbce8374d;
    11'b01000011011: data <= 32'h35713636;
    11'b01000011100: data <= 32'h3fac3aa8;
    11'b01000011101: data <= 32'h3d843e93;
    11'b01000011110: data <= 32'hb9cb3e98;
    11'b01000011111: data <= 32'hbed63a11;
    11'b01000100000: data <= 32'hb7893149;
    11'b01000100001: data <= 32'h3cbb3361;
    11'b01000100010: data <= 32'h3d90b0ab;
    11'b01000100011: data <= 32'h39d9bd7b;
    11'b01000100100: data <= 32'h3a13bfb0;
    11'b01000100101: data <= 32'h3d6ab882;
    11'b01000100110: data <= 32'h3c973d42;
    11'b01000100111: data <= 32'ha83f3d1b;
    11'b01000101000: data <= 32'hbb6cb974;
    11'b01000101001: data <= 32'hbbd5c020;
    11'b01000101010: data <= 32'hbc13bdab;
    11'b01000101011: data <= 32'hbd9eb140;
    11'b01000101100: data <= 32'hbc6faf10;
    11'b01000101101: data <= 32'h3586b9ce;
    11'b01000101110: data <= 32'h3d9fb4ff;
    11'b01000101111: data <= 32'h373d3c89;
    11'b01000110000: data <= 32'hbe223fee;
    11'b01000110001: data <= 32'hc00e3e1d;
    11'b01000110010: data <= 32'hb8153a34;
    11'b01000110011: data <= 32'h3b0c376e;
    11'b01000110100: data <= 32'h38ce259a;
    11'b01000110101: data <= 32'hb033baba;
    11'b01000110110: data <= 32'h3807bc0c;
    11'b01000110111: data <= 32'h3fea3459;
    11'b01000111000: data <= 32'h40873e84;
    11'b01000111001: data <= 32'h3b503c8e;
    11'b01000111010: data <= 32'hb78aba10;
    11'b01000111011: data <= 32'hba31bedc;
    11'b01000111100: data <= 32'hb8f6bb34;
    11'b01000111101: data <= 32'hb98ab047;
    11'b01000111110: data <= 32'hb71bbb74;
    11'b01000111111: data <= 32'h3812c023;
    11'b01001000000: data <= 32'h3c1fbdd6;
    11'b01001000001: data <= 32'ha21838f4;
    11'b01001000010: data <= 32'hbe8b3fa9;
    11'b01001000011: data <= 32'hbf653dac;
    11'b01001000100: data <= 32'hb8f53659;
    11'b01001000101: data <= 32'h28582db0;
    11'b01001000110: data <= 32'hba302dd9;
    11'b01001000111: data <= 32'hbd3db336;
    11'b01001001000: data <= 32'h2c9db397;
    11'b01001001001: data <= 32'h406139be;
    11'b01001001010: data <= 32'h41233ec0;
    11'b01001001011: data <= 32'h3b943d14;
    11'b01001001100: data <= 32'hb84cac3a;
    11'b01001001101: data <= 32'hb7f5b83c;
    11'b01001001110: data <= 32'h31383037;
    11'b01001001111: data <= 32'h34292f77;
    11'b01001010000: data <= 32'h317cbde2;
    11'b01001010001: data <= 32'h391ac1a8;
    11'b01001010010: data <= 32'h3c2dbfaa;
    11'b01001010011: data <= 32'h362636e9;
    11'b01001010100: data <= 32'hba673e38;
    11'b01001010101: data <= 32'hbc6838fa;
    11'b01001010110: data <= 32'hb8cbb88c;
    11'b01001010111: data <= 32'hba4ab82a;
    11'b01001011000: data <= 32'hbf9e2c06;
    11'b01001011001: data <= 32'hc039220d;
    11'b01001011010: data <= 32'hb448b408;
    11'b01001011011: data <= 32'h3fa334b8;
    11'b01001011100: data <= 32'h3fdb3d14;
    11'b01001011101: data <= 32'h30e63dd9;
    11'b01001011110: data <= 32'hbc033b63;
    11'b01001011111: data <= 32'hb5243a6a;
    11'b01001100000: data <= 32'h39cd3c78;
    11'b01001100001: data <= 32'h393537a1;
    11'b01001100010: data <= 32'h301cbda5;
    11'b01001100011: data <= 32'h37afc12e;
    11'b01001100100: data <= 32'h3d68bdd5;
    11'b01001100101: data <= 32'h3d953950;
    11'b01001100110: data <= 32'h383d3caa;
    11'b01001100111: data <= 32'hb058b36b;
    11'b01001101000: data <= 32'hb5d3bd3f;
    11'b01001101001: data <= 32'hbc29ba1d;
    11'b01001101010: data <= 32'hc03f2e9a;
    11'b01001101011: data <= 32'hc029b3c8;
    11'b01001101100: data <= 32'hb4d2bc75;
    11'b01001101101: data <= 32'h3d84bae7;
    11'b01001101110: data <= 32'h3baa37cc;
    11'b01001101111: data <= 32'hba5f3de0;
    11'b01001110000: data <= 32'hbd9a3e1f;
    11'b01001110001: data <= 32'hb3f13dd6;
    11'b01001110010: data <= 32'h399b3df0;
    11'b01001110011: data <= 32'h2eba39d7;
    11'b01001110100: data <= 32'hb9dfbad4;
    11'b01001110101: data <= 32'ha9bcbe82;
    11'b01001110110: data <= 32'h3e85b817;
    11'b01001110111: data <= 32'h40a73c3a;
    11'b01001111000: data <= 32'h3e213b93;
    11'b01001111001: data <= 32'h3800b86a;
    11'b01001111010: data <= 32'ha569bcca;
    11'b01001111011: data <= 32'hb8c4b436;
    11'b01001111100: data <= 32'hbd873632;
    11'b01001111101: data <= 32'hbd5cb9b5;
    11'b01001111110: data <= 32'hac50c084;
    11'b01001111111: data <= 32'h3b93c024;
    11'b01010000000: data <= 32'h3484b3f2;
    11'b01010000001: data <= 32'hbc803cd8;
    11'b01010000010: data <= 32'hbd053d68;
    11'b01010000011: data <= 32'hb01a3c4d;
    11'b01010000100: data <= 32'h325d3c4d;
    11'b01010000101: data <= 32'hbc3d39ff;
    11'b01010000110: data <= 32'hbfe7b260;
    11'b01010000111: data <= 32'hb9d3b960;
    11'b01010001000: data <= 32'h3e6b30d4;
    11'b01010001001: data <= 32'h41143caf;
    11'b01010001010: data <= 32'h3e553b07;
    11'b01010001011: data <= 32'h3736b223;
    11'b01010001100: data <= 32'h33a8b34a;
    11'b01010001101: data <= 32'h32fb3aa1;
    11'b01010001110: data <= 32'hb47b3b47;
    11'b01010001111: data <= 32'hb82ebbd4;
    11'b01010010000: data <= 32'h305fc1ce;
    11'b01010010001: data <= 32'h3a5dc121;
    11'b01010010010: data <= 32'h35d4b80a;
    11'b01010010011: data <= 32'hb8193a97;
    11'b01010010100: data <= 32'hb758382e;
    11'b01010010101: data <= 32'h3198a0fd;
    11'b01010010110: data <= 32'hb51f3499;
    11'b01010010111: data <= 32'hc01f3913;
    11'b01010011000: data <= 32'hc1ad3167;
    11'b01010011001: data <= 32'hbcc2b650;
    11'b01010011010: data <= 32'h3cfea95a;
    11'b01010011011: data <= 32'h3f9239c9;
    11'b01010011100: data <= 32'h39963a55;
    11'b01010011101: data <= 32'hb12f37a9;
    11'b01010011110: data <= 32'h35423bb0;
    11'b01010011111: data <= 32'h3b0f3f93;
    11'b01010100000: data <= 32'h36113dc4;
    11'b01010100001: data <= 32'hb544ba5f;
    11'b01010100010: data <= 32'ha648c13a;
    11'b01010100011: data <= 32'h3ab7c018;
    11'b01010100100: data <= 32'h3c30b146;
    11'b01010100101: data <= 32'h394d3814;
    11'b01010100110: data <= 32'h38ccb69d;
    11'b01010100111: data <= 32'h3903bbf8;
    11'b01010101000: data <= 32'hb683b23b;
    11'b01010101001: data <= 32'hc06f3933;
    11'b01010101010: data <= 32'hc18e30e3;
    11'b01010101011: data <= 32'hbca5bb6c;
    11'b01010101100: data <= 32'h3a28bc1e;
    11'b01010101101: data <= 32'h3a88b0f7;
    11'b01010101110: data <= 32'hb78a3860;
    11'b01010101111: data <= 32'hba5b3b03;
    11'b01010110000: data <= 32'h35a33e31;
    11'b01010110001: data <= 32'h3c464089;
    11'b01010110010: data <= 32'h31053ec0;
    11'b01010110011: data <= 32'hbc05b424;
    11'b01010110100: data <= 32'hb918be59;
    11'b01010110101: data <= 32'h3ac5bb3d;
    11'b01010110110: data <= 32'h3ef13741;
    11'b01010110111: data <= 32'h3e5735b8;
    11'b01010111000: data <= 32'h3d1fbb54;
    11'b01010111001: data <= 32'h3c15bcca;
    11'b01010111010: data <= 32'h2b202ea4;
    11'b01010111011: data <= 32'hbdae3c04;
    11'b01010111100: data <= 32'hbf7da90e;
    11'b01010111101: data <= 32'hb9c5bf36;
    11'b01010111110: data <= 32'h36a6c04b;
    11'b01010111111: data <= 32'ha4d4bbbb;
    11'b01011000000: data <= 32'hbc6c31bd;
    11'b01011000001: data <= 32'hbaf23918;
    11'b01011000010: data <= 32'h38263c70;
    11'b01011000011: data <= 32'h3ab83eee;
    11'b01011000100: data <= 32'hb9c73e20;
    11'b01011000101: data <= 32'hc04a3513;
    11'b01011000110: data <= 32'hbdacb7e4;
    11'b01011000111: data <= 32'h39452aee;
    11'b01011001000: data <= 32'h3f603a6c;
    11'b01011001001: data <= 32'h3e553451;
    11'b01011001010: data <= 32'h3c96ba8c;
    11'b01011001011: data <= 32'h3c99b833;
    11'b01011001100: data <= 32'h3a6b3c52;
    11'b01011001101: data <= 32'hb24b3e8c;
    11'b01011001110: data <= 32'hba2dae85;
    11'b01011001111: data <= 32'hb44fc09d;
    11'b01011010000: data <= 32'h345ec12e;
    11'b01011010001: data <= 32'hb1e5bcbb;
    11'b01011010010: data <= 32'hba69b02a;
    11'b01011010011: data <= 32'hb297b0ad;
    11'b01011010100: data <= 32'h3b7aad27;
    11'b01011010101: data <= 32'h386d3976;
    11'b01011010110: data <= 32'hbe343ca8;
    11'b01011010111: data <= 32'hc1ea3935;
    11'b01011011000: data <= 32'hbf882329;
    11'b01011011001: data <= 32'h352d31bb;
    11'b01011011010: data <= 32'h3cda381a;
    11'b01011011011: data <= 32'h38d82d07;
    11'b01011011100: data <= 32'h34d1b669;
    11'b01011011101: data <= 32'h3bf9376c;
    11'b01011011110: data <= 32'h3da84031;
    11'b01011011111: data <= 32'h3962406d;
    11'b01011100000: data <= 32'hb40e2f6c;
    11'b01011100001: data <= 32'hb3cfc000;
    11'b01011100010: data <= 32'h3363bff6;
    11'b01011100011: data <= 32'h3385b92a;
    11'b01011100100: data <= 32'h30c5b330;
    11'b01011100101: data <= 32'h3a69bc17;
    11'b01011100110: data <= 32'h3dddbd0a;
    11'b01011100111: data <= 32'h3870b00e;
    11'b01011101000: data <= 32'hbea53bba;
    11'b01011101001: data <= 32'hc1a9398e;
    11'b01011101010: data <= 32'hbecdb40e;
    11'b01011101011: data <= 32'h27a9b879;
    11'b01011101100: data <= 32'h3227b4d8;
    11'b01011101101: data <= 32'hb9f0b45b;
    11'b01011101110: data <= 32'hb93fb070;
    11'b01011101111: data <= 32'h3a473bcd;
    11'b01011110000: data <= 32'h3e8740d7;
    11'b01011110001: data <= 32'h39b340b4;
    11'b01011110010: data <= 32'hb9433817;
    11'b01011110011: data <= 32'hba2fbc12;
    11'b01011110100: data <= 32'h2fa0b978;
    11'b01011110101: data <= 32'h39fa3496;
    11'b01011110110: data <= 32'h3bbfb01c;
    11'b01011110111: data <= 32'h3dc9be23;
    11'b01011111000: data <= 32'h3f3abede;
    11'b01011111001: data <= 32'h3b65afc4;
    11'b01011111010: data <= 32'hbb243cd6;
    11'b01011111011: data <= 32'hbf1a38f5;
    11'b01011111100: data <= 32'hbbb6bb61;
    11'b01011111101: data <= 32'hacabbe2e;
    11'b01011111110: data <= 32'hb913bc5c;
    11'b01011111111: data <= 32'hbe81b91a;
    11'b01100000000: data <= 32'hbc2bb56e;
    11'b01100000001: data <= 32'h3a7b3867;
    11'b01100000010: data <= 32'h3e0a3f08;
    11'b01100000011: data <= 32'h2b9b3fb8;
    11'b01100000100: data <= 32'hbe8e3ac1;
    11'b01100000101: data <= 32'hbe222b2d;
    11'b01100000110: data <= 32'haf0c3828;
    11'b01100000111: data <= 32'h3abb3bbc;
    11'b01100001000: data <= 32'h3bada9a3;
    11'b01100001001: data <= 32'h3cdabe1c;
    11'b01100001010: data <= 32'h3ed8bd22;
    11'b01100001011: data <= 32'h3dcc395b;
    11'b01100001100: data <= 32'h34e13f44;
    11'b01100001101: data <= 32'hb709390e;
    11'b01100001110: data <= 32'hb157bd74;
    11'b01100001111: data <= 32'ha325bfd8;
    11'b01100010000: data <= 32'hbafbbcef;
    11'b01100010001: data <= 32'hbe4bba30;
    11'b01100010010: data <= 32'hb8c0bb79;
    11'b01100010011: data <= 32'h3cbfb8e9;
    11'b01100010100: data <= 32'h3d4737c3;
    11'b01100010101: data <= 32'hb9573cdb;
    11'b01100010110: data <= 32'hc0cf3b9d;
    11'b01100010111: data <= 32'hbfcd38f1;
    11'b01100011000: data <= 32'hb5373b42;
    11'b01100011001: data <= 32'h35b43b64;
    11'b01100011010: data <= 32'h1ab1b197;
    11'b01100011011: data <= 32'h313dbcde;
    11'b01100011100: data <= 32'h3cdfb6e3;
    11'b01100011101: data <= 32'h3f493e7a;
    11'b01100011110: data <= 32'h3cd940bb;
    11'b01100011111: data <= 32'h359d3a42;
    11'b01100100000: data <= 32'h307abca3;
    11'b01100100001: data <= 32'h2868bd81;
    11'b01100100010: data <= 32'hb884b823;
    11'b01100100011: data <= 32'hba4fb869;
    11'b01100100100: data <= 32'h3538be48;
    11'b01100100101: data <= 32'h3ed5bf46;
    11'b01100100110: data <= 32'h3d35b8cf;
    11'b01100100111: data <= 32'hbaae399c;
    11'b01100101000: data <= 32'hc0913af5;
    11'b01100101001: data <= 32'hbe783750;
    11'b01100101010: data <= 32'hb56635d1;
    11'b01100101011: data <= 32'hb6f63325;
    11'b01100101100: data <= 32'hbd72b82e;
    11'b01100101101: data <= 32'hbc47bbd1;
    11'b01100101110: data <= 32'h39562e49;
    11'b01100101111: data <= 32'h3f843fc9;
    11'b01100110000: data <= 32'h3d6540c7;
    11'b01100110001: data <= 32'h315a3b81;
    11'b01100110010: data <= 32'hb3a6b628;
    11'b01100110011: data <= 32'hac6dab25;
    11'b01100110100: data <= 32'haee13980;
    11'b01100110101: data <= 32'h2093ae82;
    11'b01100110110: data <= 32'h3bc0bf94;
    11'b01100110111: data <= 32'h3fdfc0b9;
    11'b01100111000: data <= 32'h3decbab9;
    11'b01100111001: data <= 32'hb3f23a09;
    11'b01100111010: data <= 32'hbce13a28;
    11'b01100111011: data <= 32'hb8f7b04c;
    11'b01100111100: data <= 32'had52b881;
    11'b01100111101: data <= 32'hbc3ab868;
    11'b01100111110: data <= 32'hc0a6babb;
    11'b01100111111: data <= 32'hbee4bc28;
    11'b01101000000: data <= 32'h3762b19d;
    11'b01101000001: data <= 32'h3ed23d1f;
    11'b01101000010: data <= 32'h3a493ee9;
    11'b01101000011: data <= 32'hb9bf3b61;
    11'b01101000100: data <= 32'hbbc1379c;
    11'b01101000101: data <= 32'hb4723ce2;
    11'b01101000110: data <= 32'h2cc63e9d;
    11'b01101000111: data <= 32'h2f95340e;
    11'b01101001000: data <= 32'h39e9bf3a;
    11'b01101001001: data <= 32'h3ea9c00c;
    11'b01101001010: data <= 32'h3eb7b1b2;
    11'b01101001011: data <= 32'h39e03d3a;
    11'b01101001100: data <= 32'h31eb3a35;
    11'b01101001101: data <= 32'h37a7b8f3;
    11'b01101001110: data <= 32'h3486bc40;
    11'b01101001111: data <= 32'hbcbeb9a6;
    11'b01101010000: data <= 32'hc0beba7a;
    11'b01101010001: data <= 32'hbdbfbd5e;
    11'b01101010010: data <= 32'h3a04bc87;
    11'b01101010011: data <= 32'h3e0caaf5;
    11'b01101010100: data <= 32'h2a94399e;
    11'b01101010101: data <= 32'hbe24398e;
    11'b01101010110: data <= 32'hbd9b3b36;
    11'b01101010111: data <= 32'hb5e03edc;
    11'b01101011000: data <= 32'hb1293f3e;
    11'b01101011001: data <= 32'hb92833e6;
    11'b01101011010: data <= 32'hb5c8bdf3;
    11'b01101011011: data <= 32'h3af3bcc4;
    11'b01101011100: data <= 32'h3ec93a55;
    11'b01101011101: data <= 32'h3def3f7e;
    11'b01101011110: data <= 32'h3c573ab3;
    11'b01101011111: data <= 32'h3c18b8f1;
    11'b01101100000: data <= 32'h37fdb937;
    11'b01101100001: data <= 32'hbad62a3b;
    11'b01101100010: data <= 32'hbe87b4d3;
    11'b01101100011: data <= 32'hb83ebe7d;
    11'b01101100100: data <= 32'h3d23c053;
    11'b01101100101: data <= 32'h3dbfbd03;
    11'b01101100110: data <= 32'hb46bad6f;
    11'b01101100111: data <= 32'hbe473658;
    11'b01101101000: data <= 32'hbc2e3994;
    11'b01101101001: data <= 32'hafb63cf2;
    11'b01101101010: data <= 32'hb8e03ca5;
    11'b01101101011: data <= 32'hbf50ae41;
    11'b01101101100: data <= 32'hbed3bcdc;
    11'b01101101101: data <= 32'h23efb858;
    11'b01101101110: data <= 32'h3dfa3d04;
    11'b01101101111: data <= 32'h3e363f8e;
    11'b01101110000: data <= 32'h3be53a27;
    11'b01101110001: data <= 32'h39eab142;
    11'b01101110010: data <= 32'h36ca37cb;
    11'b01101110011: data <= 32'hb6173d72;
    11'b01101110100: data <= 32'hba03377a;
    11'b01101110101: data <= 32'h334fbe9a;
    11'b01101110110: data <= 32'h3e39c13a;
    11'b01101110111: data <= 32'h3db9be5f;
    11'b01101111000: data <= 32'h2496b18b;
    11'b01101111001: data <= 32'hb9783362;
    11'b01101111010: data <= 32'h2aa02dff;
    11'b01101111011: data <= 32'h37583431;
    11'b01101111100: data <= 32'hbb4934b7;
    11'b01101111101: data <= 32'hc15db714;
    11'b01101111110: data <= 32'hc0f3bc88;
    11'b01101111111: data <= 32'hb611b873;
    11'b01110000000: data <= 32'h3cd83a19;
    11'b01110000001: data <= 32'h3bc63c90;
    11'b01110000010: data <= 32'h2d7136f0;
    11'b01110000011: data <= 32'haaad35cf;
    11'b01110000100: data <= 32'h31e23e91;
    11'b01110000101: data <= 32'hadf840eb;
    11'b01110000110: data <= 32'hb6a93c39;
    11'b01110000111: data <= 32'h3172bda0;
    11'b01110001000: data <= 32'h3cc1c07f;
    11'b01110001001: data <= 32'h3d4ebb8d;
    11'b01110001010: data <= 32'h39513672;
    11'b01110001011: data <= 32'h38bb3431;
    11'b01110001100: data <= 32'h3d2db772;
    11'b01110001101: data <= 32'h3c65b6d9;
    11'b01110001110: data <= 32'hbab9a6f0;
    11'b01110001111: data <= 32'hc160b5fb;
    11'b01110010000: data <= 32'hc076bca6;
    11'b01110010001: data <= 32'haee3bcbb;
    11'b01110010010: data <= 32'h3c19b6f0;
    11'b01110010011: data <= 32'h31dda85a;
    11'b01110010100: data <= 32'hbb19ae76;
    11'b01110010101: data <= 32'hb9233868;
    11'b01110010110: data <= 32'h2eb8402a;
    11'b01110010111: data <= 32'hadec4160;
    11'b01110011000: data <= 32'hbaea3c77;
    11'b01110011001: data <= 32'hba43bc44;
    11'b01110011010: data <= 32'h33e7bd7e;
    11'b01110011011: data <= 32'h3c1230cd;
    11'b01110011100: data <= 32'h3c933c73;
    11'b01110011101: data <= 32'h3db8355a;
    11'b01110011110: data <= 32'h3fc6b94d;
    11'b01110011111: data <= 32'h3dbeb4f8;
    11'b01110100000: data <= 32'hb7433894;
    11'b01110100001: data <= 32'hbfa53439;
    11'b01110100010: data <= 32'hbcedbc71;
    11'b01110100011: data <= 32'h3862bfae;
    11'b01110100100: data <= 32'h3bcabe3e;
    11'b01110100101: data <= 32'hb4efbba2;
    11'b01110100110: data <= 32'hbcc6b899;
    11'b01110100111: data <= 32'hb72b3404;
    11'b01110101000: data <= 32'h37583e4a;
    11'b01110101001: data <= 32'hb2f53feb;
    11'b01110101010: data <= 32'hbef8396b;
    11'b01110101011: data <= 32'hc018ba97;
    11'b01110101100: data <= 32'hba19b8b8;
    11'b01110101101: data <= 32'h38b43ae4;
    11'b01110101110: data <= 32'h3c4c3d30;
    11'b01110101111: data <= 32'h3d3331f4;
    11'b01110110000: data <= 32'h3e90b81b;
    11'b01110110001: data <= 32'h3d383826;
    11'b01110110010: data <= 32'h9c6e3f2e;
    11'b01110110011: data <= 32'hbb5e3ccf;
    11'b01110110100: data <= 32'hb3e2baf4;
    11'b01110110101: data <= 32'h3bf4c063;
    11'b01110110110: data <= 32'h3b55bf7a;
    11'b01110110111: data <= 32'hb4b3bc45;
    11'b01110111000: data <= 32'hb8eab9e0;
    11'b01110111001: data <= 32'h3863b584;
    11'b01110111010: data <= 32'h3cd83812;
    11'b01110111011: data <= 32'hb3103b4d;
    11'b01110111100: data <= 32'hc0c530fc;
    11'b01110111101: data <= 32'hc191b9c0;
    11'b01110111110: data <= 32'hbce5b59d;
    11'b01110111111: data <= 32'h34113963;
    11'b01111000000: data <= 32'h37943950;
    11'b01111000001: data <= 32'h3534b511;
    11'b01111000010: data <= 32'h3971b4d1;
    11'b01111000011: data <= 32'h3b2c3dc2;
    11'b01111000100: data <= 32'h348541b8;
    11'b01111000101: data <= 32'hb5cd3f97;
    11'b01111000110: data <= 32'h9df1b825;
    11'b01111000111: data <= 32'h3a15bf1a;
    11'b01111001000: data <= 32'h3949bca3;
    11'b01111001001: data <= 32'h2815b5c0;
    11'b01111001010: data <= 32'h3686b873;
    11'b01111001011: data <= 32'h3f08bb1d;
    11'b01111001100: data <= 32'h3ff8b604;
    11'b01111001101: data <= 32'h219c34cc;
    11'b01111001110: data <= 32'hc09b2c81;
    11'b01111001111: data <= 32'hc0fbb8fb;
    11'b01111010000: data <= 32'hbae7b948;
    11'b01111010001: data <= 32'h31cbb412;
    11'b01111010010: data <= 32'hb4c6b792;
    11'b01111010011: data <= 32'hba89bc14;
    11'b01111010100: data <= 32'hb204b526;
    11'b01111010101: data <= 32'h39293f0e;
    11'b01111010110: data <= 32'h360b421a;
    11'b01111010111: data <= 32'hb80b3fa9;
    11'b01111011000: data <= 32'hb96cb3f5;
    11'b01111011001: data <= 32'hb036bb43;
    11'b01111011010: data <= 32'h31572d59;
    11'b01111011011: data <= 32'h343238e2;
    11'b01111011100: data <= 32'h3c68b4cf;
    11'b01111011101: data <= 32'h40c5bc9a;
    11'b01111011110: data <= 32'h40adb85e;
    11'b01111011111: data <= 32'h360538dd;
    11'b01111100000: data <= 32'hbe14391d;
    11'b01111100001: data <= 32'hbd71b61f;
    11'b01111100010: data <= 32'h27bbbc7a;
    11'b01111100011: data <= 32'h350abcd9;
    11'b01111100100: data <= 32'hbaa3bd8a;
    11'b01111100101: data <= 32'hbd90be37;
    11'b01111100110: data <= 32'hb4adb93b;
    11'b01111100111: data <= 32'h3b3f3ce8;
    11'b01111101000: data <= 32'h36e34078;
    11'b01111101001: data <= 32'hbc593d13;
    11'b01111101010: data <= 32'hbeffb1cd;
    11'b01111101011: data <= 32'hbc8fae71;
    11'b01111101100: data <= 32'hb5ee3c2e;
    11'b01111101101: data <= 32'h2ebb3c66;
    11'b01111101110: data <= 32'h3b66b547;
    11'b01111101111: data <= 32'h3ffdbca3;
    11'b01111110000: data <= 32'h4014a4cb;
    11'b01111110001: data <= 32'h395c3e78;
    11'b01111110010: data <= 32'hb8203e4f;
    11'b01111110011: data <= 32'hb07f1be7;
    11'b01111110100: data <= 32'h3a46bd03;
    11'b01111110101: data <= 32'h366dbdce;
    11'b01111110110: data <= 32'hbb9bbdc2;
    11'b01111110111: data <= 32'hbc75be64;
    11'b01111111000: data <= 32'h378dbc82;
    11'b01111111001: data <= 32'h3e9930de;
    11'b01111111010: data <= 32'h38c63b9c;
    11'b01111111011: data <= 32'hbe303711;
    11'b01111111100: data <= 32'hc0cab3be;
    11'b01111111101: data <= 32'hbe473400;
    11'b01111111110: data <= 32'hb9293ca2;
    11'b01111111111: data <= 32'hb6a539bf;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    