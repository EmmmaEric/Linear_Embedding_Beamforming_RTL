
module memory_rom_50(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3e4132fd;
    11'b00000000001: data <= 32'h3b6a2be1;
    11'b00000000010: data <= 32'hbb10b0a4;
    11'b00000000011: data <= 32'hbe39bc27;
    11'b00000000100: data <= 32'h26a9bee3;
    11'b00000000101: data <= 32'h3fbabd50;
    11'b00000000110: data <= 32'h3f20b8b3;
    11'b00000000111: data <= 32'ha469b853;
    11'b00000001000: data <= 32'hbcb7b945;
    11'b00000001001: data <= 32'hbb6d31de;
    11'b00000001010: data <= 32'hb93d3d84;
    11'b00000001011: data <= 32'hbd053c54;
    11'b00000001100: data <= 32'hbee6ba5d;
    11'b00000001101: data <= 32'hbc2fbfa2;
    11'b00000001110: data <= 32'h2ca5b923;
    11'b00000001111: data <= 32'h37a43e10;
    11'b00000010000: data <= 32'h36f7402b;
    11'b00000010001: data <= 32'h3a853c19;
    11'b00000010010: data <= 32'h3cae35f0;
    11'b00000010011: data <= 32'h35c83b59;
    11'b00000010100: data <= 32'hbc5d3ce0;
    11'b00000010101: data <= 32'hbc9e3115;
    11'b00000010110: data <= 32'h39c9bcf4;
    11'b00000010111: data <= 32'h40cebe0f;
    11'b00000011000: data <= 32'h3fa2bb56;
    11'b00000011001: data <= 32'h3221b882;
    11'b00000011010: data <= 32'hb6aeb717;
    11'b00000011011: data <= 32'h34e63179;
    11'b00000011100: data <= 32'h36a33a87;
    11'b00000011101: data <= 32'hbbab319a;
    11'b00000011110: data <= 32'hc06ebe14;
    11'b00000011111: data <= 32'hbf21c05e;
    11'b00000100000: data <= 32'hb5d5ba24;
    11'b00000100001: data <= 32'h36173c23;
    11'b00000100010: data <= 32'h34413cac;
    11'b00000100011: data <= 32'h32b432c3;
    11'b00000100100: data <= 32'h339e34fb;
    11'b00000100101: data <= 32'hb68e3ee1;
    11'b00000100110: data <= 32'hbd6c40ab;
    11'b00000100111: data <= 32'hbc573b84;
    11'b00000101000: data <= 32'h390cbb9b;
    11'b00000101001: data <= 32'h3fb4bd5a;
    11'b00000101010: data <= 32'h3db4b6d7;
    11'b00000101011: data <= 32'h358532fa;
    11'b00000101100: data <= 32'h38b13217;
    11'b00000101101: data <= 32'h3eb43464;
    11'b00000101110: data <= 32'h3da837a9;
    11'b00000101111: data <= 32'hb901b065;
    11'b00000110000: data <= 32'hc06abdf1;
    11'b00000110001: data <= 32'hbe56c00d;
    11'b00000110010: data <= 32'h2fe5bc3a;
    11'b00000110011: data <= 32'h3a279c94;
    11'b00000110100: data <= 32'h3067b3ff;
    11'b00000110101: data <= 32'hb685baae;
    11'b00000110110: data <= 32'hb6b22c36;
    11'b00000110111: data <= 32'hb9bd4006;
    11'b00000111000: data <= 32'hbda64122;
    11'b00000111001: data <= 32'hbd8e3abe;
    11'b00000111010: data <= 32'hb44dbc48;
    11'b00000111011: data <= 32'h3966bc12;
    11'b00000111100: data <= 32'h3825363e;
    11'b00000111101: data <= 32'h349b3c67;
    11'b00000111110: data <= 32'h3ce33974;
    11'b00000111111: data <= 32'h40be3609;
    11'b00001000000: data <= 32'h3eee3922;
    11'b00001000001: data <= 32'hb82737a2;
    11'b00001000010: data <= 32'hbf4ab874;
    11'b00001000011: data <= 32'hb9e3bd90;
    11'b00001000100: data <= 32'h3c44bcfa;
    11'b00001000101: data <= 32'h3d23bb8b;
    11'b00001000110: data <= 32'h2ff8bd4e;
    11'b00001000111: data <= 32'hb840bdf6;
    11'b00001001000: data <= 32'hb236b1a1;
    11'b00001001001: data <= 32'hb1873edd;
    11'b00001001010: data <= 32'hbc553f97;
    11'b00001001011: data <= 32'hbf3528ae;
    11'b00001001100: data <= 32'hbda4bde7;
    11'b00001001101: data <= 32'hb8f4ba64;
    11'b00001001110: data <= 32'hb4ea3afd;
    11'b00001001111: data <= 32'h2a283d3d;
    11'b00001010000: data <= 32'h3c9f380c;
    11'b00001010001: data <= 32'h401c346f;
    11'b00001010010: data <= 32'h3cf13caa;
    11'b00001010011: data <= 32'hb9b53eb3;
    11'b00001010100: data <= 32'hbd933a27;
    11'b00001010101: data <= 32'h2c23b8b9;
    11'b00001010110: data <= 32'h3ea3bca6;
    11'b00001010111: data <= 32'h3d9cbcd4;
    11'b00001011000: data <= 32'h2fa3bdcc;
    11'b00001011001: data <= 32'hacf1bd8d;
    11'b00001011010: data <= 32'h3afdb35a;
    11'b00001011011: data <= 32'h3c133c8d;
    11'b00001011100: data <= 32'hb7483b5e;
    11'b00001011101: data <= 32'hbff7ba50;
    11'b00001011110: data <= 32'hc01fbf0a;
    11'b00001011111: data <= 32'hbcb4ba01;
    11'b00001100000: data <= 32'hb8893958;
    11'b00001100001: data <= 32'hb26c3875;
    11'b00001100010: data <= 32'h384cb6b0;
    11'b00001100011: data <= 32'h3c5aaf53;
    11'b00001100100: data <= 32'h362e3e94;
    11'b00001100101: data <= 32'hbbfd4161;
    11'b00001100110: data <= 32'hbcc23ebf;
    11'b00001100111: data <= 32'h32ebadc4;
    11'b00001101000: data <= 32'h3d5ebae2;
    11'b00001101001: data <= 32'h3aa0b99b;
    11'b00001101010: data <= 32'haa0db950;
    11'b00001101011: data <= 32'h38c8b9a9;
    11'b00001101100: data <= 32'h4044ae77;
    11'b00001101101: data <= 32'h4056399c;
    11'b00001101110: data <= 32'h304a365b;
    11'b00001101111: data <= 32'hbf40bb52;
    11'b00001110000: data <= 32'hbf59be21;
    11'b00001110001: data <= 32'hb9bcb9ef;
    11'b00001110010: data <= 32'hb185a9a2;
    11'b00001110011: data <= 32'hb4feb9f2;
    11'b00001110100: data <= 32'hb0cdbe80;
    11'b00001110101: data <= 32'h340cb939;
    11'b00001110110: data <= 32'hacf53ee6;
    11'b00001110111: data <= 32'hbc1041c4;
    11'b00001111000: data <= 32'hbce73e9a;
    11'b00001111001: data <= 32'hb5d9b167;
    11'b00001111010: data <= 32'h32eab848;
    11'b00001111011: data <= 32'hb3c9315e;
    11'b00001111100: data <= 32'hb6c835d0;
    11'b00001111101: data <= 32'h3be7ac62;
    11'b00001111110: data <= 32'h4190a14b;
    11'b00001111111: data <= 32'h41283913;
    11'b00010000000: data <= 32'h355639ab;
    11'b00010000001: data <= 32'hbd90afa8;
    11'b00010000010: data <= 32'hbb95b9ef;
    11'b00010000011: data <= 32'h3567b8c2;
    11'b00010000100: data <= 32'h379ab9af;
    11'b00010000101: data <= 32'hb50ebf11;
    11'b00010000110: data <= 32'hb773c0ce;
    11'b00010000111: data <= 32'h3236bc29;
    11'b00010001000: data <= 32'h35283d6e;
    11'b00010001001: data <= 32'hb863405b;
    11'b00010001010: data <= 32'hbd363a21;
    11'b00010001011: data <= 32'hbcdeb973;
    11'b00010001100: data <= 32'hbc13b562;
    11'b00010001101: data <= 32'hbce33a78;
    11'b00010001110: data <= 32'hbae73aaa;
    11'b00010001111: data <= 32'h3a7badb6;
    11'b00010010000: data <= 32'h40deb316;
    11'b00010010001: data <= 32'h40153aae;
    11'b00010010010: data <= 32'h2c173e6b;
    11'b00010010011: data <= 32'hbbdc3c8e;
    11'b00010010100: data <= 32'ha4653387;
    11'b00010010101: data <= 32'h3cadb43a;
    11'b00010010110: data <= 32'h3a0bba9c;
    11'b00010010111: data <= 32'hb66fbf73;
    11'b00010011000: data <= 32'hb4fec09a;
    11'b00010011001: data <= 32'h3babbc3e;
    11'b00010011010: data <= 32'h3dbe3a52;
    11'b00010011011: data <= 32'h34443c60;
    11'b00010011100: data <= 32'hbcd2b469;
    11'b00010011101: data <= 32'hbebbbc87;
    11'b00010011110: data <= 32'hbe36b390;
    11'b00010011111: data <= 32'hbe1d3b04;
    11'b00010100000: data <= 32'hbc843617;
    11'b00010100001: data <= 32'h31ecbb5f;
    11'b00010100010: data <= 32'h3d82ba63;
    11'b00010100011: data <= 32'h3c013c03;
    11'b00010100100: data <= 32'hb62f40d0;
    11'b00010100101: data <= 32'hba044012;
    11'b00010100110: data <= 32'h36183a9d;
    11'b00010100111: data <= 32'h3c972f3a;
    11'b00010101000: data <= 32'h349eb494;
    11'b00010101001: data <= 32'hb9f1bc07;
    11'b00010101010: data <= 32'h293dbddc;
    11'b00010101011: data <= 32'h3fedba39;
    11'b00010101100: data <= 32'h41213590;
    11'b00010101101: data <= 32'h3be63599;
    11'b00010101110: data <= 32'hbb27b98a;
    11'b00010101111: data <= 32'hbd92bc20;
    11'b00010110000: data <= 32'hbc27acb4;
    11'b00010110001: data <= 32'hbc1337cc;
    11'b00010110010: data <= 32'hbc71b95a;
    11'b00010110011: data <= 32'hb7f2c036;
    11'b00010110100: data <= 32'h3590be00;
    11'b00010110101: data <= 32'h340d3b30;
    11'b00010110110: data <= 32'hb86a4101;
    11'b00010110111: data <= 32'hb9483fd5;
    11'b00010111000: data <= 32'h2f623971;
    11'b00010111001: data <= 32'h348f3585;
    11'b00010111010: data <= 32'hba0a389c;
    11'b00010111011: data <= 32'hbd38321b;
    11'b00010111100: data <= 32'h3280b86e;
    11'b00010111101: data <= 32'h4102b82a;
    11'b00010111110: data <= 32'h41e631dd;
    11'b00010111111: data <= 32'h3cad35b6;
    11'b00011000000: data <= 32'hb825b188;
    11'b00011000001: data <= 32'hb7ffb482;
    11'b00011000010: data <= 32'h313b3459;
    11'b00011000011: data <= 32'haf962d3e;
    11'b00011000100: data <= 32'hbb82be2d;
    11'b00011000101: data <= 32'hbb0ac1c0;
    11'b00011000110: data <= 32'h1505bfaf;
    11'b00011000111: data <= 32'h35d63833;
    11'b00011001000: data <= 32'hb0b13f1b;
    11'b00011001001: data <= 32'hb8513b96;
    11'b00011001010: data <= 32'hb733ab4c;
    11'b00011001011: data <= 32'hba3e35ec;
    11'b00011001100: data <= 32'hbef43d0c;
    11'b00011001101: data <= 32'hbf503b70;
    11'b00011001110: data <= 32'ha82bb46e;
    11'b00011001111: data <= 32'h403cb924;
    11'b00011010000: data <= 32'h409d3263;
    11'b00011010001: data <= 32'h39ae3b9f;
    11'b00011010010: data <= 32'hb44c3b29;
    11'b00011010011: data <= 32'h376339aa;
    11'b00011010100: data <= 32'h3cfb39db;
    11'b00011010101: data <= 32'h376f2cdd;
    11'b00011010110: data <= 32'hbb42be54;
    11'b00011010111: data <= 32'hbb1dc164;
    11'b00011011000: data <= 32'h3757bf30;
    11'b00011011001: data <= 32'h3d102ddf;
    11'b00011011010: data <= 32'h39713956;
    11'b00011011011: data <= 32'hb472b53e;
    11'b00011011100: data <= 32'hba11ba7d;
    11'b00011011101: data <= 32'hbcf53544;
    11'b00011011110: data <= 32'hbffe3de0;
    11'b00011011111: data <= 32'hc0013a45;
    11'b00011100000: data <= 32'hb878bb02;
    11'b00011100001: data <= 32'h3c26bce1;
    11'b00011100010: data <= 32'h3c3631c9;
    11'b00011100011: data <= 32'ha8e33e39;
    11'b00011100100: data <= 32'hb24f3ecb;
    11'b00011100101: data <= 32'h3bcd3d21;
    11'b00011100110: data <= 32'h3e1d3c4d;
    11'b00011100111: data <= 32'h3406387b;
    11'b00011101000: data <= 32'hbceab99a;
    11'b00011101001: data <= 32'hb9d8beac;
    11'b00011101010: data <= 32'h3d03bcec;
    11'b00011101011: data <= 32'h4091b1d2;
    11'b00011101100: data <= 32'h3da1b18b;
    11'b00011101101: data <= 32'h2b54bc2f;
    11'b00011101110: data <= 32'hb79ebbe4;
    11'b00011101111: data <= 32'hb98c372c;
    11'b00011110000: data <= 32'hbd4e3d16;
    11'b00011110001: data <= 32'hbeeba36f;
    11'b00011110010: data <= 32'hbc4abfba;
    11'b00011110011: data <= 32'hac9fbfc7;
    11'b00011110100: data <= 32'h1dbc1852;
    11'b00011110101: data <= 32'hb8013e71;
    11'b00011110110: data <= 32'hb1b33e54;
    11'b00011110111: data <= 32'h3b273c09;
    11'b00011111000: data <= 32'h3b7b3c61;
    11'b00011111001: data <= 32'hb9243d13;
    11'b00011111010: data <= 32'hbf4b3885;
    11'b00011111011: data <= 32'hb978b774;
    11'b00011111100: data <= 32'h3ec5b947;
    11'b00011111101: data <= 32'h413eb3d1;
    11'b00011111110: data <= 32'h3dffb568;
    11'b00011111111: data <= 32'h3457ba81;
    11'b00100000000: data <= 32'h349eb690;
    11'b00100000001: data <= 32'h388a3a99;
    11'b00100000010: data <= 32'hb0d43c0d;
    11'b00100000011: data <= 32'hbcf1ba25;
    11'b00100000100: data <= 32'hbd4fc14b;
    11'b00100000101: data <= 32'hb89ac0a0;
    11'b00100000110: data <= 32'hb1e4b43c;
    11'b00100000111: data <= 32'hb4cb3bd7;
    11'b00100001000: data <= 32'ha8d53823;
    11'b00100001001: data <= 32'h37f824a8;
    11'b00100001010: data <= 32'h265a3a70;
    11'b00100001011: data <= 32'hbe443f3c;
    11'b00100001100: data <= 32'hc0a83dc7;
    11'b00100001101: data <= 32'hbaf32ff7;
    11'b00100001110: data <= 32'h3d75b858;
    11'b00100001111: data <= 32'h3fb7b336;
    11'b00100010000: data <= 32'h3a852cd9;
    11'b00100010001: data <= 32'h33362c6a;
    11'b00100010010: data <= 32'h3c663813;
    11'b00100010011: data <= 32'h3f1d3d31;
    11'b00100010100: data <= 32'h3a073c09;
    11'b00100010101: data <= 32'hbb79baa3;
    11'b00100010110: data <= 32'hbd38c0d9;
    11'b00100010111: data <= 32'hb4d8bffe;
    11'b00100011000: data <= 32'h3802b6ec;
    11'b00100011001: data <= 32'h3700240c;
    11'b00100011010: data <= 32'h3422bb06;
    11'b00100011011: data <= 32'h33b0bc3e;
    11'b00100011100: data <= 32'hb6c23778;
    11'b00100011101: data <= 32'hbf283fd2;
    11'b00100011110: data <= 32'hc0b63ded;
    11'b00100011111: data <= 32'hbcadb365;
    11'b00100100000: data <= 32'h36a6bc03;
    11'b00100100001: data <= 32'h3880b493;
    11'b00100100010: data <= 32'hb41738b3;
    11'b00100100011: data <= 32'ha4923a9c;
    11'b00100100100: data <= 32'h3e1d3c37;
    11'b00100100101: data <= 32'h407b3e28;
    11'b00100100110: data <= 32'h3a7c3d44;
    11'b00100100111: data <= 32'hbc6cabfd;
    11'b00100101000: data <= 32'hbcbbbd2d;
    11'b00100101001: data <= 32'h35ebbc7c;
    11'b00100101010: data <= 32'h3dc2b624;
    11'b00100101011: data <= 32'h3c8db9c6;
    11'b00100101100: data <= 32'h384bbf18;
    11'b00100101101: data <= 32'h3663be20;
    11'b00100101110: data <= 32'h27d13668;
    11'b00100101111: data <= 32'hbc213f1f;
    11'b00100110000: data <= 32'hbf2d3a9a;
    11'b00100110001: data <= 32'hbd75bcb2;
    11'b00100110010: data <= 32'hb8a2beca;
    11'b00100110011: data <= 32'hb946b721;
    11'b00100110100: data <= 32'hbc2739b4;
    11'b00100110101: data <= 32'hb3173a39;
    11'b00100110110: data <= 32'h3dce39b4;
    11'b00100110111: data <= 32'h3f383d3a;
    11'b00100111000: data <= 32'h2bba3ee7;
    11'b00100111001: data <= 32'hbea13c55;
    11'b00100111010: data <= 32'hbc942d0a;
    11'b00100111011: data <= 32'h3aa9b2b5;
    11'b00100111100: data <= 32'h3f46b1ff;
    11'b00100111101: data <= 32'h3cb8baf5;
    11'b00100111110: data <= 32'h3857bed9;
    11'b00100111111: data <= 32'h3b2abc89;
    11'b00101000000: data <= 32'h3cb239b6;
    11'b00101000001: data <= 32'h34e53e31;
    11'b00101000010: data <= 32'hbb9a2dab;
    11'b00101000011: data <= 32'hbd52bfa1;
    11'b00101000100: data <= 32'hbc2dc010;
    11'b00101000101: data <= 32'hbc23b868;
    11'b00101000110: data <= 32'hbc3934f9;
    11'b00101000111: data <= 32'hb187b1b1;
    11'b00101001000: data <= 32'h3c5bb6d8;
    11'b00101001001: data <= 32'h3b90395b;
    11'b00101001010: data <= 32'hbada3fd4;
    11'b00101001011: data <= 32'hc0493f9f;
    11'b00101001100: data <= 32'hbcdb3aeb;
    11'b00101001101: data <= 32'h39853150;
    11'b00101001110: data <= 32'h3ce5a912;
    11'b00101001111: data <= 32'h35ccb7d1;
    11'b00101010000: data <= 32'h3149bb4d;
    11'b00101010001: data <= 32'h3d93b3fd;
    11'b00101010010: data <= 32'h40a03cb5;
    11'b00101010011: data <= 32'h3da73de2;
    11'b00101010100: data <= 32'hb59faf78;
    11'b00101010101: data <= 32'hbc8dbf16;
    11'b00101010110: data <= 32'hba5cbe6c;
    11'b00101010111: data <= 32'hb75fb6a1;
    11'b00101011000: data <= 32'hb632b595;
    11'b00101011001: data <= 32'h2f35bdfb;
    11'b00101011010: data <= 32'h3a5bbedb;
    11'b00101011011: data <= 32'h36541c18;
    11'b00101011100: data <= 32'hbca13f92;
    11'b00101011101: data <= 32'hc02b3fcf;
    11'b00101011110: data <= 32'hbcfb392f;
    11'b00101011111: data <= 32'h275db1e9;
    11'b00101100000: data <= 32'habf8ace1;
    11'b00101100001: data <= 32'hbb542810;
    11'b00101100010: data <= 32'hb6d5adf1;
    11'b00101100011: data <= 32'h3e5135cd;
    11'b00101100100: data <= 32'h418b3d73;
    11'b00101100101: data <= 32'h3e893e35;
    11'b00101100110: data <= 32'hb5e63633;
    11'b00101100111: data <= 32'hbbbbb9c9;
    11'b00101101000: data <= 32'hb02eb837;
    11'b00101101001: data <= 32'h38039dd4;
    11'b00101101010: data <= 32'h35d4ba8e;
    11'b00101101011: data <= 32'h35c8c0c1;
    11'b00101101100: data <= 32'h3a32c0be;
    11'b00101101101: data <= 32'h38eab437;
    11'b00101101110: data <= 32'hb7c43e8c;
    11'b00101101111: data <= 32'hbd5a3d3f;
    11'b00101110000: data <= 32'hbc54b48b;
    11'b00101110001: data <= 32'hb979bb41;
    11'b00101110010: data <= 32'hbd0eb32d;
    11'b00101110011: data <= 32'hbfa334a8;
    11'b00101110100: data <= 32'hbb052bb7;
    11'b00101110101: data <= 32'h3d892f13;
    11'b00101110110: data <= 32'h40b53bc3;
    11'b00101110111: data <= 32'h3b6d3e78;
    11'b00101111000: data <= 32'hbb5a3cfb;
    11'b00101111001: data <= 32'hbb6338fc;
    11'b00101111010: data <= 32'h36d538ea;
    11'b00101111011: data <= 32'h3c3237b2;
    11'b00101111100: data <= 32'h37f7ba82;
    11'b00101111101: data <= 32'h33aac0ab;
    11'b00101111110: data <= 32'h3ba7c01c;
    11'b00101111111: data <= 32'h3de42295;
    11'b00110000000: data <= 32'h3a8c3d94;
    11'b00110000001: data <= 32'hb40e3813;
    11'b00110000010: data <= 32'hb9c7bc9d;
    11'b00110000011: data <= 32'hbbb1bd55;
    11'b00110000100: data <= 32'hbea2b386;
    11'b00110000101: data <= 32'hc0173151;
    11'b00110000110: data <= 32'hbb48b8fc;
    11'b00110000111: data <= 32'h3bffbbe5;
    11'b00110001000: data <= 32'h3dcf2df6;
    11'b00110001001: data <= 32'hae003e00;
    11'b00110001010: data <= 32'hbdf83f67;
    11'b00110001011: data <= 32'hbb6d3db7;
    11'b00110001100: data <= 32'h382e3c98;
    11'b00110001101: data <= 32'h39ae3a17;
    11'b00110001110: data <= 32'hb443b637;
    11'b00110001111: data <= 32'hb5d8be0d;
    11'b00110010000: data <= 32'h3c62bc64;
    11'b00110010001: data <= 32'h40c0386d;
    11'b00110010010: data <= 32'h3fc83d1e;
    11'b00110010011: data <= 32'h38542e9e;
    11'b00110010100: data <= 32'hb57bbd05;
    11'b00110010101: data <= 32'hb91ebbc4;
    11'b00110010110: data <= 32'hbc502ee3;
    11'b00110010111: data <= 32'hbd5fb07e;
    11'b00110011000: data <= 32'hb889bec4;
    11'b00110011001: data <= 32'h397ac094;
    11'b00110011010: data <= 32'h39e6ba63;
    11'b00110011011: data <= 32'hb8ea3cca;
    11'b00110011100: data <= 32'hbe0c3f2b;
    11'b00110011101: data <= 32'hba413ce0;
    11'b00110011110: data <= 32'h32613a78;
    11'b00110011111: data <= 32'hb52b3996;
    11'b00110100000: data <= 32'hbe3b309f;
    11'b00110100001: data <= 32'hbcd1b87a;
    11'b00110100010: data <= 32'h3c02b490;
    11'b00110100011: data <= 32'h41653aa8;
    11'b00110100100: data <= 32'h405e3cdc;
    11'b00110100101: data <= 32'h38a834aa;
    11'b00110100110: data <= 32'hb0f5b762;
    11'b00110100111: data <= 32'h29452f4d;
    11'b00110101000: data <= 32'ha27f3a32;
    11'b00110101001: data <= 32'hb6a4b4cd;
    11'b00110101010: data <= 32'hb2dfc0d3;
    11'b00110101011: data <= 32'h3870c1f4;
    11'b00110101100: data <= 32'h3955bcb0;
    11'b00110101101: data <= 32'hb2503b00;
    11'b00110101110: data <= 32'hba2e3c7c;
    11'b00110101111: data <= 32'hb5c532b5;
    11'b00110110000: data <= 32'hb1d5ab8f;
    11'b00110110001: data <= 32'hbd623724;
    11'b00110110010: data <= 32'hc13037b5;
    11'b00110110011: data <= 32'hbf3bb0b9;
    11'b00110110100: data <= 32'h3983b48a;
    11'b00110110101: data <= 32'h4076377a;
    11'b00110110110: data <= 32'h3db13c24;
    11'b00110110111: data <= 32'hacf23a76;
    11'b00110111000: data <= 32'hb2863987;
    11'b00110111001: data <= 32'h393b3d3b;
    11'b00110111010: data <= 32'h3a1a3dd4;
    11'b00110111011: data <= 32'ha820b007;
    11'b00110111100: data <= 32'hb48dc09a;
    11'b00110111101: data <= 32'h3820c142;
    11'b00110111110: data <= 32'h3cbdbaa1;
    11'b00110111111: data <= 32'h3b30399f;
    11'b00111000000: data <= 32'h35e4346e;
    11'b00111000001: data <= 32'h336ebae1;
    11'b00111000010: data <= 32'hb3d2b9cf;
    11'b00111000011: data <= 32'hbe9b35c4;
    11'b00111000100: data <= 32'hc1723860;
    11'b00111000101: data <= 32'hbf4ab7ff;
    11'b00111000110: data <= 32'h3574bca4;
    11'b00111000111: data <= 32'h3d2ab75c;
    11'b00111001000: data <= 32'h333d394b;
    11'b00111001001: data <= 32'hbb083ca1;
    11'b00111001010: data <= 32'hb4d13d90;
    11'b00111001011: data <= 32'h3b433f75;
    11'b00111001100: data <= 32'h39eb3f19;
    11'b00111001101: data <= 32'hb88634da;
    11'b00111001110: data <= 32'hbb66bdc2;
    11'b00111001111: data <= 32'h363fbe18;
    11'b00111010000: data <= 32'h3f34ad09;
    11'b00111010001: data <= 32'h3f9c3984;
    11'b00111010010: data <= 32'h3cd7b425;
    11'b00111010011: data <= 32'h39a6bd0b;
    11'b00111010100: data <= 32'h301fb8d6;
    11'b00111010101: data <= 32'hbc1d39be;
    11'b00111010110: data <= 32'hbf9c3802;
    11'b00111010111: data <= 32'hbd30bd0e;
    11'b00111011000: data <= 32'h302bc0a6;
    11'b00111011001: data <= 32'h3780bdac;
    11'b00111011010: data <= 32'hb89e32c2;
    11'b00111011011: data <= 32'hbc983bfc;
    11'b00111011100: data <= 32'hb1463c85;
    11'b00111011101: data <= 32'h3aa73dc2;
    11'b00111011110: data <= 32'h253f3e47;
    11'b00111011111: data <= 32'hbed139ef;
    11'b00111100000: data <= 32'hbf5db662;
    11'b00111100001: data <= 32'h2eaab71c;
    11'b00111100010: data <= 32'h3fe73757;
    11'b00111100011: data <= 32'h4029394e;
    11'b00111100100: data <= 32'h3cd0b4c9;
    11'b00111100101: data <= 32'h3a6bba49;
    11'b00111100110: data <= 32'h39e734fe;
    11'b00111100111: data <= 32'h2f233ddc;
    11'b00111101000: data <= 32'hb9d73886;
    11'b00111101001: data <= 32'hb977bf31;
    11'b00111101010: data <= 32'h2c1bc1e3;
    11'b00111101011: data <= 32'h322abf1f;
    11'b00111101100: data <= 32'hb7b2ace9;
    11'b00111101101: data <= 32'hb8c435d7;
    11'b00111101110: data <= 32'h354c2ae6;
    11'b00111101111: data <= 32'h399035a8;
    11'b00111110000: data <= 32'hba443c41;
    11'b00111110001: data <= 32'hc1533bf5;
    11'b00111110010: data <= 32'hc0f0323b;
    11'b00111110011: data <= 32'hb36eafca;
    11'b00111110100: data <= 32'h3e0634da;
    11'b00111110101: data <= 32'h3d0736cd;
    11'b00111110110: data <= 32'h35b7a90e;
    11'b00111110111: data <= 32'h38292fcc;
    11'b00111111000: data <= 32'h3d063db0;
    11'b00111111001: data <= 32'h3c2f4069;
    11'b00111111010: data <= 32'ha76d3a8d;
    11'b00111111011: data <= 32'hb828be93;
    11'b00111111100: data <= 32'h9f8ac111;
    11'b00111111101: data <= 32'h3742bd25;
    11'b00111111110: data <= 32'h3591aa32;
    11'b00111111111: data <= 32'h3733b632;
    11'b01000000000: data <= 32'h3c06bca0;
    11'b01000000001: data <= 32'h3a1bb8fe;
    11'b01000000010: data <= 32'hbc0a39cb;
    11'b01000000011: data <= 32'hc17a3c3f;
    11'b01000000100: data <= 32'hc0bf2dcd;
    11'b01000000101: data <= 32'hb6bfb9b4;
    11'b01000000110: data <= 32'h392ab817;
    11'b01000000111: data <= 32'hac50a9cd;
    11'b01000001000: data <= 32'hb9f33066;
    11'b01000001001: data <= 32'h310339a8;
    11'b01000001010: data <= 32'h3df03fb9;
    11'b01000001011: data <= 32'h3d0740ea;
    11'b01000001100: data <= 32'hb42d3c8e;
    11'b01000001101: data <= 32'hbc17babb;
    11'b01000001110: data <= 32'hb359bd40;
    11'b01000001111: data <= 32'h3ae9b40e;
    11'b01000010000: data <= 32'h3cd032ac;
    11'b01000010001: data <= 32'h3cffbb03;
    11'b01000010010: data <= 32'h3ddabf1c;
    11'b01000010011: data <= 32'h3c55ba89;
    11'b01000010100: data <= 32'hb6bb3b55;
    11'b01000010101: data <= 32'hbf423c68;
    11'b01000010110: data <= 32'hbe5db727;
    11'b01000010111: data <= 32'hb5e7becb;
    11'b01000011000: data <= 32'haf64bdb3;
    11'b01000011001: data <= 32'hbc51b82e;
    11'b01000011010: data <= 32'hbd5ba706;
    11'b01000011011: data <= 32'h2e52373a;
    11'b01000011100: data <= 32'h3de63dae;
    11'b01000011101: data <= 32'h3a33400f;
    11'b01000011110: data <= 32'hbcc73d55;
    11'b01000011111: data <= 32'hbf8e3033;
    11'b01000100000: data <= 32'hb89da89b;
    11'b01000100001: data <= 32'h3bd638f4;
    11'b01000100010: data <= 32'h3d6d367a;
    11'b01000100011: data <= 32'h3cb2bbaf;
    11'b01000100100: data <= 32'h3d88be2d;
    11'b01000100101: data <= 32'h3decb026;
    11'b01000100110: data <= 32'h39373e67;
    11'b01000100111: data <= 32'hb74d3cff;
    11'b01000101000: data <= 32'hb919bb02;
    11'b01000101001: data <= 32'hb1fac086;
    11'b01000101010: data <= 32'hb699bef3;
    11'b01000101011: data <= 32'hbceab97b;
    11'b01000101100: data <= 32'hbc2bb7e1;
    11'b01000101101: data <= 32'h3817b886;
    11'b01000101110: data <= 32'h3dbb3140;
    11'b01000101111: data <= 32'h2f2f3cc4;
    11'b01000110000: data <= 32'hc0253d48;
    11'b01000110001: data <= 32'hc0f639c9;
    11'b01000110010: data <= 32'hbab53845;
    11'b01000110011: data <= 32'h390639fd;
    11'b01000110100: data <= 32'h389e3472;
    11'b01000110101: data <= 32'h31a4ba60;
    11'b01000110110: data <= 32'h3a4cba76;
    11'b01000110111: data <= 32'h3eea3b01;
    11'b01000111000: data <= 32'h3e4440a1;
    11'b01000111001: data <= 32'h37d93de7;
    11'b01000111010: data <= 32'hb126ba51;
    11'b01000111011: data <= 32'haf37bf86;
    11'b01000111100: data <= 32'hb3b1bc73;
    11'b01000111101: data <= 32'hb8c2b5fc;
    11'b01000111110: data <= 32'hb016bbe0;
    11'b01000111111: data <= 32'h3cabbefb;
    11'b01001000000: data <= 32'h3e11bc39;
    11'b01001000001: data <= 32'hb04b3821;
    11'b01001000010: data <= 32'hc0513cd2;
    11'b01001000011: data <= 32'hc08f398c;
    11'b01001000100: data <= 32'hba483112;
    11'b01001000101: data <= 32'h1dad2e35;
    11'b01001000110: data <= 32'hb9b4b16a;
    11'b01001000111: data <= 32'hbca4b95c;
    11'b01001001000: data <= 32'h2ca6b3e7;
    11'b01001001001: data <= 32'h3ef93d85;
    11'b01001001010: data <= 32'h3f5640fb;
    11'b01001001011: data <= 32'h37db3e66;
    11'b01001001100: data <= 32'hb770b23c;
    11'b01001001101: data <= 32'hb4bab989;
    11'b01001001110: data <= 32'h2e2f30b2;
    11'b01001001111: data <= 32'h323a33a3;
    11'b01001010000: data <= 32'h3936bcf2;
    11'b01001010001: data <= 32'h3e4dc0cf;
    11'b01001010010: data <= 32'h3ec5bdfa;
    11'b01001010011: data <= 32'h3488378d;
    11'b01001010100: data <= 32'hbd103cb7;
    11'b01001010101: data <= 32'hbd2433af;
    11'b01001010110: data <= 32'hb61fb9cd;
    11'b01001010111: data <= 32'hb80eba38;
    11'b01001011000: data <= 32'hbf03b8fa;
    11'b01001011001: data <= 32'hc007b9f3;
    11'b01001011010: data <= 32'hb424b5ed;
    11'b01001011011: data <= 32'h3e893b31;
    11'b01001011100: data <= 32'h3dc03f82;
    11'b01001011101: data <= 32'hb4ef3dda;
    11'b01001011110: data <= 32'hbd103837;
    11'b01001011111: data <= 32'hb90f38d6;
    11'b01001100000: data <= 32'h34143d28;
    11'b01001100001: data <= 32'h370139f2;
    11'b01001100010: data <= 32'h38d5bcc1;
    11'b01001100011: data <= 32'h3d5dc082;
    11'b01001100100: data <= 32'h3f28bbc3;
    11'b01001100101: data <= 32'h3c733c3d;
    11'b01001100110: data <= 32'h2ebc3d47;
    11'b01001100111: data <= 32'hab0fb22c;
    11'b01001101000: data <= 32'h3064bd5b;
    11'b01001101001: data <= 32'hb91ebc73;
    11'b01001101010: data <= 32'hbfebb955;
    11'b01001101011: data <= 32'hbfa3bb9d;
    11'b01001101100: data <= 32'h25c0bca5;
    11'b01001101101: data <= 32'h3e50b5d1;
    11'b01001101110: data <= 32'h3a663a1c;
    11'b01001101111: data <= 32'hbccc3c5d;
    11'b01001110000: data <= 32'hbf7f3b6b;
    11'b01001110001: data <= 32'hba7e3cfe;
    11'b01001110010: data <= 32'h2f233e90;
    11'b01001110011: data <= 32'hb0783a4f;
    11'b01001110100: data <= 32'hb64abbf4;
    11'b01001110101: data <= 32'h37c0be41;
    11'b01001110110: data <= 32'h3eb022f9;
    11'b01001110111: data <= 32'h3f423f21;
    11'b01001111000: data <= 32'h3c7c3df9;
    11'b01001111001: data <= 32'h3963b441;
    11'b01001111010: data <= 32'h36dfbc84;
    11'b01001111011: data <= 32'hb69ab7ef;
    11'b01001111100: data <= 32'hbda1af8e;
    11'b01001111101: data <= 32'hbc34bc5a;
    11'b01001111110: data <= 32'h395ec03c;
    11'b01001111111: data <= 32'h3e88be97;
    11'b01010000000: data <= 32'h3702b20e;
    11'b01010000001: data <= 32'hbdb839b3;
    11'b01010000010: data <= 32'hbec13a80;
    11'b01010000011: data <= 32'hb8683b92;
    11'b01010000100: data <= 32'hb1ac3c55;
    11'b01010000101: data <= 32'hbcd335f5;
    11'b01010000110: data <= 32'hbf28bad7;
    11'b01010000111: data <= 32'hb831bb6d;
    11'b01010001000: data <= 32'h3d883915;
    11'b01010001001: data <= 32'h3fdc3fef;
    11'b01010001010: data <= 32'h3cd03dc9;
    11'b01010001011: data <= 32'h380a26b0;
    11'b01010001100: data <= 32'h3500b107;
    11'b01010001101: data <= 32'hac563a89;
    11'b01010001110: data <= 32'hb8a13a5e;
    11'b01010001111: data <= 32'hb1d7bc08;
    11'b01010010000: data <= 32'h3c75c144;
    11'b01010010001: data <= 32'h3eb5c059;
    11'b01010010010: data <= 32'h38b6b693;
    11'b01010010011: data <= 32'hb9f1389c;
    11'b01010010100: data <= 32'hb933357f;
    11'b01010010101: data <= 32'h30d12af0;
    11'b01010010110: data <= 32'hb57330db;
    11'b01010010111: data <= 32'hc02aaf9d;
    11'b01010011000: data <= 32'hc179baad;
    11'b01010011001: data <= 32'hbc4bba9a;
    11'b01010011010: data <= 32'h3c783594;
    11'b01010011011: data <= 32'h3e253d5b;
    11'b01010011100: data <= 32'h36b83c18;
    11'b01010011101: data <= 32'hb514364f;
    11'b01010011110: data <= 32'hab323bb7;
    11'b01010011111: data <= 32'h30db401e;
    11'b01010100000: data <= 32'hb0cf3e38;
    11'b01010100001: data <= 32'haa2cba0b;
    11'b01010100010: data <= 32'h3af4c0dc;
    11'b01010100011: data <= 32'h3e0ebebe;
    11'b01010100100: data <= 32'h3c483113;
    11'b01010100101: data <= 32'h372039d8;
    11'b01010100110: data <= 32'h397ab01c;
    11'b01010100111: data <= 32'h3ba7b9a5;
    11'b01010101000: data <= 32'hb33cb595;
    11'b01010101001: data <= 32'hc079b195;
    11'b01010101010: data <= 32'hc160ba8c;
    11'b01010101011: data <= 32'hbad5bd24;
    11'b01010101100: data <= 32'h3c2fb9cd;
    11'b01010101101: data <= 32'h3af62fe6;
    11'b01010101110: data <= 32'hb8a9357c;
    11'b01010101111: data <= 32'hbc4a3813;
    11'b01010110000: data <= 32'hb43c3e10;
    11'b01010110001: data <= 32'h322c40fb;
    11'b01010110010: data <= 32'hb6c63ed8;
    11'b01010110011: data <= 32'hbad5b815;
    11'b01010110100: data <= 32'had10bed9;
    11'b01010110101: data <= 32'h3c50b8f8;
    11'b01010110110: data <= 32'h3dd63c04;
    11'b01010110111: data <= 32'h3d693b91;
    11'b01010111000: data <= 32'h3e0eb591;
    11'b01010111001: data <= 32'h3da5ba2b;
    11'b01010111010: data <= 32'h2e092ce8;
    11'b01010111011: data <= 32'hbe8a3729;
    11'b01010111100: data <= 32'hbf1db923;
    11'b01010111101: data <= 32'haf05bfa5;
    11'b01010111110: data <= 32'h3c96bf8b;
    11'b01010111111: data <= 32'h3650bb98;
    11'b01011000000: data <= 32'hbc3bb3f6;
    11'b01011000001: data <= 32'hbc4e3412;
    11'b01011000010: data <= 32'h29f73cb5;
    11'b01011000011: data <= 32'h32573fa7;
    11'b01011000100: data <= 32'hbca03cf0;
    11'b01011000101: data <= 32'hc03bb693;
    11'b01011000110: data <= 32'hbce0bbe9;
    11'b01011000111: data <= 32'h384132f5;
    11'b01011001000: data <= 32'h3db13d93;
    11'b01011001001: data <= 32'h3d8d3afc;
    11'b01011001010: data <= 32'h3d71b52d;
    11'b01011001011: data <= 32'h3d1eb00c;
    11'b01011001100: data <= 32'h36a73cfb;
    11'b01011001101: data <= 32'hb9e73dfd;
    11'b01011001110: data <= 32'hb9c5b45e;
    11'b01011001111: data <= 32'h3828c067;
    11'b01011010000: data <= 32'h3cc3c0b5;
    11'b01011010001: data <= 32'h34efbce2;
    11'b01011010010: data <= 32'hb981b6ca;
    11'b01011010011: data <= 32'hb217b307;
    11'b01011010100: data <= 32'h3b0a3360;
    11'b01011010101: data <= 32'h357c3a96;
    11'b01011010110: data <= 32'hbf193889;
    11'b01011010111: data <= 32'hc1fdb6a2;
    11'b01011011000: data <= 32'hbf67b973;
    11'b01011011001: data <= 32'h3170338b;
    11'b01011011010: data <= 32'h3b9b3b4e;
    11'b01011011011: data <= 32'h3874354b;
    11'b01011011100: data <= 32'h36a1b457;
    11'b01011011101: data <= 32'h3a0939b8;
    11'b01011011110: data <= 32'h38c440d4;
    11'b01011011111: data <= 32'hb06240bc;
    11'b01011100000: data <= 32'hb4be302d;
    11'b01011100001: data <= 32'h373cbfa5;
    11'b01011100010: data <= 32'h3b72bf49;
    11'b01011100011: data <= 32'h37a6b882;
    11'b01011100100: data <= 32'h3293b0a5;
    11'b01011100101: data <= 32'h3c41b930;
    11'b01011100110: data <= 32'h3f4bb962;
    11'b01011100111: data <= 32'h39442a6d;
    11'b01011101000: data <= 32'hbf36351d;
    11'b01011101001: data <= 32'hc1ceb549;
    11'b01011101010: data <= 32'hbe56babf;
    11'b01011101011: data <= 32'h31d8b845;
    11'b01011101100: data <= 32'h351ab2cb;
    11'b01011101101: data <= 32'hb888b809;
    11'b01011101110: data <= 32'hb8bcb665;
    11'b01011101111: data <= 32'h35873c6c;
    11'b01011110000: data <= 32'h3963419c;
    11'b01011110001: data <= 32'hb04b410a;
    11'b01011110010: data <= 32'hba583574;
    11'b01011110011: data <= 32'hb641bcd6;
    11'b01011110100: data <= 32'h355bb936;
    11'b01011110101: data <= 32'h38b73813;
    11'b01011110110: data <= 32'h3b5e3455;
    11'b01011110111: data <= 32'h3f6fbb04;
    11'b01011111000: data <= 32'h40a3bbe8;
    11'b01011111001: data <= 32'h3bfd314b;
    11'b01011111010: data <= 32'hbcc43a87;
    11'b01011111011: data <= 32'hbf9c9799;
    11'b01011111100: data <= 32'hb91dbcb0;
    11'b01011111101: data <= 32'h379abde6;
    11'b01011111110: data <= 32'hb0b5bd02;
    11'b01011111111: data <= 32'hbd11bcba;
    11'b01100000000: data <= 32'hbb3cb9dc;
    11'b01100000001: data <= 32'h381339d4;
    11'b01100000010: data <= 32'h3a7f404d;
    11'b01100000011: data <= 32'hb8813f83;
    11'b01100000100: data <= 32'hbf3f3446;
    11'b01100000101: data <= 32'hbdfbb80c;
    11'b01100000110: data <= 32'hb5593644;
    11'b01100000111: data <= 32'h36b53cd1;
    11'b01100001000: data <= 32'h3b1635de;
    11'b01100001001: data <= 32'h3e95bbb1;
    11'b01100001010: data <= 32'h4022b928;
    11'b01100001011: data <= 32'h3cb53c4d;
    11'b01100001100: data <= 32'hb5133f4a;
    11'b01100001101: data <= 32'hb9473821;
    11'b01100001110: data <= 32'h34a0bd1d;
    11'b01100001111: data <= 32'h39a8bf5e;
    11'b01100010000: data <= 32'hb50bbdec;
    11'b01100010001: data <= 32'hbcc3bd26;
    11'b01100010010: data <= 32'hb4a9bc6d;
    11'b01100010011: data <= 32'h3d25b270;
    11'b01100010100: data <= 32'h3c7a3b2b;
    11'b01100010101: data <= 32'hbbad3b60;
    11'b01100010110: data <= 32'hc11f2bbf;
    11'b01100010111: data <= 32'hc032b08e;
    11'b01100011000: data <= 32'hb971398a;
    11'b01100011001: data <= 32'h9d7c3c0b;
    11'b01100011010: data <= 32'h2b6cae5e;
    11'b01100011011: data <= 32'h3870bc4d;
    11'b01100011100: data <= 32'h3d19aab3;
    11'b01100011101: data <= 32'h3c98402e;
    11'b01100011110: data <= 32'h350e415b;
    11'b01100011111: data <= 32'h28a93ba3;
    11'b01100100000: data <= 32'h3834bbda;
    11'b01100100001: data <= 32'h3863bd2b;
    11'b01100100010: data <= 32'hb4e1b99e;
    11'b01100100011: data <= 32'hb886ba32;
    11'b01100100100: data <= 32'h3a4ebd57;
    11'b01100100101: data <= 32'h4072bc7a;
    11'b01100100110: data <= 32'h3e0fb053;
    11'b01100100111: data <= 32'hbb6c35b8;
    11'b01100101000: data <= 32'hc0dd22be;
    11'b01100101001: data <= 32'hbef0b125;
    11'b01100101010: data <= 32'hb79f328f;
    11'b01100101011: data <= 32'hb75c2d4a;
    11'b01100101100: data <= 32'hbc4abb72;
    11'b01100101101: data <= 32'hb98dbd49;
    11'b01100101110: data <= 32'h38523363;
    11'b01100101111: data <= 32'h3c4340d9;
    11'b01100110000: data <= 32'h370c4183;
    11'b01100110001: data <= 32'hb1723c17;
    11'b01100110010: data <= 32'hae19b6c3;
    11'b01100110011: data <= 32'ha893af6a;
    11'b01100110100: data <= 32'hb56a38c7;
    11'b01100110101: data <= 32'h0e5fa879;
    11'b01100110110: data <= 32'h3e0abd85;
    11'b01100110111: data <= 32'h4159be21;
    11'b01100111000: data <= 32'h3f11b502;
    11'b01100111001: data <= 32'hb6b538d6;
    11'b01100111010: data <= 32'hbdae34fb;
    11'b01100111011: data <= 32'hb8a8b545;
    11'b01100111100: data <= 32'h301bb866;
    11'b01100111101: data <= 32'hb9d6baf0;
    11'b01100111110: data <= 32'hbf67be5d;
    11'b01100111111: data <= 32'hbd33be7c;
    11'b01101000000: data <= 32'h36d9ad99;
    11'b01101000001: data <= 32'h3c963f05;
    11'b01101000010: data <= 32'h31963fba;
    11'b01101000011: data <= 32'hbbc93944;
    11'b01101000100: data <= 32'hbc5b2d50;
    11'b01101000101: data <= 32'hb9ac3bed;
    11'b01101000110: data <= 32'hb83e3e57;
    11'b01101000111: data <= 32'ha58a35c9;
    11'b01101001000: data <= 32'h3d1abd81;
    11'b01101001001: data <= 32'h408abd61;
    11'b01101001010: data <= 32'h3ec035ba;
    11'b01101001011: data <= 32'h34433de7;
    11'b01101001100: data <= 32'hafe83ac0;
    11'b01101001101: data <= 32'h3919b5de;
    11'b01101001110: data <= 32'h3973bb12;
    11'b01101001111: data <= 32'hba3dbc46;
    11'b01101010000: data <= 32'hbfadbe53;
    11'b01101010001: data <= 32'hbb8ebf22;
    11'b01101010010: data <= 32'h3c2bbac8;
    11'b01101010011: data <= 32'h3dde373c;
    11'b01101010100: data <= 32'haf9e3989;
    11'b01101010101: data <= 32'hbe982f6e;
    11'b01101010110: data <= 32'hbea234d6;
    11'b01101010111: data <= 32'hbbd43db4;
    11'b01101011000: data <= 32'hba5f3eab;
    11'b01101011001: data <= 32'hb9ab2d9d;
    11'b01101011010: data <= 32'h309ebdf7;
    11'b01101011011: data <= 32'h3cd5bb08;
    11'b01101011100: data <= 32'h3d483d0c;
    11'b01101011101: data <= 32'h39e04093;
    11'b01101011110: data <= 32'h39913cf6;
    11'b01101011111: data <= 32'h3cabb183;
    11'b01101100000: data <= 32'h3a00b70a;
    11'b01101100001: data <= 32'hba05b415;
    11'b01101100010: data <= 32'hbdbdba9a;
    11'b01101100011: data <= 32'h9f87bebc;
    11'b01101100100: data <= 32'h3fb2be5b;
    11'b01101100101: data <= 32'h3f66b989;
    11'b01101100110: data <= 32'hb05ab1da;
    11'b01101100111: data <= 32'hbe59b23f;
    11'b01101101000: data <= 32'hbd0d33b8;
    11'b01101101001: data <= 32'hb8833c59;
    11'b01101101010: data <= 32'hbb963b4b;
    11'b01101101011: data <= 32'hbea5b95e;
    11'b01101101100: data <= 32'hbcd4befc;
    11'b01101101101: data <= 32'h30f0b8c0;
    11'b01101101110: data <= 32'h3b813e84;
    11'b01101101111: data <= 32'h3a4b40ae;
    11'b01101110000: data <= 32'h39233c8c;
    11'b01101110001: data <= 32'h3a032fbc;
    11'b01101110010: data <= 32'h3436388d;
    11'b01101110011: data <= 32'hba723c8e;
    11'b01101110100: data <= 32'hbb423390;
    11'b01101110101: data <= 32'h39b9bd9d;
    11'b01101110110: data <= 32'h40b6bf9a;
    11'b01101110111: data <= 32'h3fe2bc17;
    11'b01101111000: data <= 32'h30d4b193;
    11'b01101111001: data <= 32'hb9cea766;
    11'b01101111010: data <= 32'ha66e2ded;
    11'b01101111011: data <= 32'h35b03679;
    11'b01101111100: data <= 32'hbb0c9f5e;
    11'b01101111101: data <= 32'hc0a2bd45;
    11'b01101111110: data <= 32'hbfdcbfd6;
    11'b01101111111: data <= 32'hb34ab9e8;
    11'b01110000000: data <= 32'h3ac63c5c;
    11'b01110000001: data <= 32'h383a3dc2;
    11'b01110000010: data <= 32'habe93795;
    11'b01110000011: data <= 32'hb1ae34a1;
    11'b01110000100: data <= 32'hb6543e27;
    11'b01110000101: data <= 32'hbb9a408d;
    11'b01110000110: data <= 32'hba6f3b72;
    11'b01110000111: data <= 32'h38b9bcbe;
    11'b01110001000: data <= 32'h3f90becd;
    11'b01110001001: data <= 32'h3e7cb784;
    11'b01110001010: data <= 32'h381638c5;
    11'b01110001011: data <= 32'h36dc37a6;
    11'b01110001100: data <= 32'h3d6028f7;
    11'b01110001101: data <= 32'h3ceb9e27;
    11'b01110001110: data <= 32'hb96cb4bd;
    11'b01110001111: data <= 32'hc0b2bd11;
    11'b01110010000: data <= 32'hbef7bf8c;
    11'b01110010001: data <= 32'h33efbcc8;
    11'b01110010010: data <= 32'h3c7bac72;
    11'b01110010011: data <= 32'h339e2acb;
    11'b01110010100: data <= 32'hba2ab683;
    11'b01110010101: data <= 32'hba793320;
    11'b01110010110: data <= 32'hb9243fac;
    11'b01110010111: data <= 32'hbc1c4102;
    11'b01110011000: data <= 32'hbce23aae;
    11'b01110011001: data <= 32'hb669bce5;
    11'b01110011010: data <= 32'h3987bcfb;
    11'b01110011011: data <= 32'h3b4236e8;
    11'b01110011100: data <= 32'h39583dc6;
    11'b01110011101: data <= 32'h3cb33af0;
    11'b01110011110: data <= 32'h40122dd5;
    11'b01110011111: data <= 32'h3e1332a1;
    11'b01110100000: data <= 32'hb84b3624;
    11'b01110100001: data <= 32'hbf7eb635;
    11'b01110100010: data <= 32'hbab4bdcb;
    11'b01110100011: data <= 32'h3c8cbe72;
    11'b01110100100: data <= 32'h3e03bc81;
    11'b01110100101: data <= 32'h2fbebbf9;
    11'b01110100110: data <= 32'hbb30bbd9;
    11'b01110100111: data <= 32'hb84f1f6d;
    11'b01110101000: data <= 32'hb0153e53;
    11'b01110101001: data <= 32'hbae63f3e;
    11'b01110101010: data <= 32'hbf642e5d;
    11'b01110101011: data <= 32'hbe9ebde9;
    11'b01110101100: data <= 32'hb861bb27;
    11'b01110101101: data <= 32'h33233b95;
    11'b01110101110: data <= 32'h382f3e72;
    11'b01110101111: data <= 32'h3c74397f;
    11'b01110110000: data <= 32'h3ed72e65;
    11'b01110110001: data <= 32'h3c5f3b38;
    11'b01110110010: data <= 32'hb8a43eb1;
    11'b01110110011: data <= 32'hbd3a3ae2;
    11'b01110110100: data <= 32'h98e4bab1;
    11'b01110110101: data <= 32'h3eb2bebf;
    11'b01110110110: data <= 32'h3e4bbdbf;
    11'b01110110111: data <= 32'h312fbc6f;
    11'b01110111000: data <= 32'hb544bb61;
    11'b01110111001: data <= 32'h38bbb187;
    11'b01110111010: data <= 32'h3bcb3b08;
    11'b01110111011: data <= 32'hb7233a83;
    11'b01110111100: data <= 32'hc078b91d;
    11'b01110111101: data <= 32'hc0c1bea8;
    11'b01110111110: data <= 32'hbc50baab;
    11'b01110111111: data <= 32'ha7023969;
    11'b01111000000: data <= 32'h32733a92;
    11'b01111000001: data <= 32'h366bb0ae;
    11'b01111000010: data <= 32'h39e9ad5b;
    11'b01111000011: data <= 32'h35c43e56;
    11'b01111000100: data <= 32'hb9c04189;
    11'b01111000101: data <= 32'hbc293eea;
    11'b01111000110: data <= 32'h2f4bb688;
    11'b01111000111: data <= 32'h3d4abd89;
    11'b01111001000: data <= 32'h3c49bb08;
    11'b01111001001: data <= 32'h31b5b550;
    11'b01111001010: data <= 32'h383bb5e8;
    11'b01111001011: data <= 32'h3fa5b310;
    11'b01111001100: data <= 32'h4016357d;
    11'b01111001101: data <= 32'h230334fb;
    11'b01111001110: data <= 32'hc040b9ac;
    11'b01111001111: data <= 32'hc04dbddf;
    11'b01111010000: data <= 32'hb911bbbb;
    11'b01111010001: data <= 32'h3413b1f0;
    11'b01111010010: data <= 32'had6cb818;
    11'b01111010011: data <= 32'hb669bcf3;
    11'b01111010100: data <= 32'hacecb724;
    11'b01111010101: data <= 32'ha2453f24;
    11'b01111010110: data <= 32'hb9a541fb;
    11'b01111010111: data <= 32'hbca53ece;
    11'b01111011000: data <= 32'hb8abb68d;
    11'b01111011001: data <= 32'h31f0bb59;
    11'b01111011010: data <= 32'h30832dd2;
    11'b01111011011: data <= 32'h20ee3958;
    11'b01111011100: data <= 32'h3c44309c;
    11'b01111011101: data <= 32'h4132b33e;
    11'b01111011110: data <= 32'h40e134be;
    11'b01111011111: data <= 32'h33bb39a8;
    11'b01111100000: data <= 32'hbe772e17;
    11'b01111100001: data <= 32'hbcc7ba8b;
    11'b01111100010: data <= 32'h3605bc27;
    11'b01111100011: data <= 32'h3a04bc09;
    11'b01111100100: data <= 32'hb37abe3c;
    11'b01111100101: data <= 32'hba02bfd7;
    11'b01111100110: data <= 32'hace6ba6a;
    11'b01111100111: data <= 32'h369c3d8d;
    11'b01111101000: data <= 32'hb58a4084;
    11'b01111101001: data <= 32'hbdc23b0c;
    11'b01111101010: data <= 32'hbe57ba15;
    11'b01111101011: data <= 32'hbc33b86b;
    11'b01111101100: data <= 32'hb9d43a5f;
    11'b01111101101: data <= 32'hb5463c5c;
    11'b01111101110: data <= 32'h3b502c6c;
    11'b01111101111: data <= 32'h4080b627;
    11'b01111110000: data <= 32'h3fe13937;
    11'b01111110001: data <= 32'h301f3eee;
    11'b01111110010: data <= 32'hbc2b3d58;
    11'b01111110011: data <= 32'hb25c1f24;
    11'b01111110100: data <= 32'h3c99baf4;
    11'b01111110101: data <= 32'h3b88bcc9;
    11'b01111110110: data <= 32'hb543bea6;
    11'b01111110111: data <= 32'hb805bf9d;
    11'b01111111000: data <= 32'h3a47bb9b;
    11'b01111111001: data <= 32'h3dfe396a;
    11'b01111111010: data <= 32'h34c83c81;
    11'b01111111011: data <= 32'hbe2cacf0;
    11'b01111111100: data <= 32'hc050bc4f;
    11'b01111111101: data <= 32'hbe58b62e;
    11'b01111111110: data <= 32'hbc213a96;
    11'b01111111111: data <= 32'hb9583890;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    