
module memory_rom_57(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3481be35;
    11'b00000000001: data <= 32'h2e22bb86;
    11'b00000000010: data <= 32'hb1733adf;
    11'b00000000011: data <= 32'hbc563e18;
    11'b00000000100: data <= 32'hbedfac1d;
    11'b00000000101: data <= 32'hbd10bfde;
    11'b00000000110: data <= 32'hb836bf44;
    11'b00000000111: data <= 32'hb84ca5e1;
    11'b00000001000: data <= 32'hb9a23c99;
    11'b00000001001: data <= 32'h304d3b85;
    11'b00000001010: data <= 32'h3d62399f;
    11'b00000001011: data <= 32'h3c333d24;
    11'b00000001100: data <= 32'hbab13ec8;
    11'b00000001101: data <= 32'hbfc93be7;
    11'b00000001110: data <= 32'hb94fad98;
    11'b00000001111: data <= 32'h3e0eb6c1;
    11'b00000010000: data <= 32'h4035b5b6;
    11'b00000010001: data <= 32'h3c45ba29;
    11'b00000010010: data <= 32'h369dbca0;
    11'b00000010011: data <= 32'h3b63b57f;
    11'b00000010100: data <= 32'h3cbb3c7e;
    11'b00000010101: data <= 32'h30403cb0;
    11'b00000010110: data <= 32'hbcceb9f1;
    11'b00000010111: data <= 32'hbdb8c0e6;
    11'b00000011000: data <= 32'hbad2bfd4;
    11'b00000011001: data <= 32'hb874b350;
    11'b00000011010: data <= 32'hb7633676;
    11'b00000011011: data <= 32'h3185b4a9;
    11'b00000011100: data <= 32'h3aa2b648;
    11'b00000011101: data <= 32'h30ff3b91;
    11'b00000011110: data <= 32'hbe54404e;
    11'b00000011111: data <= 32'hc0823edb;
    11'b00000100000: data <= 32'hba6e3598;
    11'b00000100001: data <= 32'h3c24b574;
    11'b00000100010: data <= 32'h3cbeb332;
    11'b00000100011: data <= 32'h3344b267;
    11'b00000100100: data <= 32'h34f2b356;
    11'b00000100101: data <= 32'h3ec0375f;
    11'b00000100110: data <= 32'h40943dbc;
    11'b00000100111: data <= 32'h3b5f3c87;
    11'b00000101000: data <= 32'hbb4eb926;
    11'b00000101001: data <= 32'hbd16bfe0;
    11'b00000101010: data <= 32'hb62bbdd1;
    11'b00000101011: data <= 32'h334eb57f;
    11'b00000101100: data <= 32'h32ccb88c;
    11'b00000101101: data <= 32'h3552bea1;
    11'b00000101110: data <= 32'h3840bda5;
    11'b00000101111: data <= 32'hb0af38c3;
    11'b00000110000: data <= 32'hbe35404b;
    11'b00000110001: data <= 32'hc02c3e1b;
    11'b00000110010: data <= 32'hbc45b0b1;
    11'b00000110011: data <= 32'h24c4ba2a;
    11'b00000110100: data <= 32'hb38cb0f9;
    11'b00000110101: data <= 32'hbaca35fd;
    11'b00000110110: data <= 32'h27ea36b8;
    11'b00000110111: data <= 32'h3fdd3a44;
    11'b00000111000: data <= 32'h410b3e00;
    11'b00000111001: data <= 32'h3a893db5;
    11'b00000111010: data <= 32'hbc4633d1;
    11'b00000111011: data <= 32'hbc04b9a9;
    11'b00000111100: data <= 32'h364fb813;
    11'b00000111101: data <= 32'h3c71b3cf;
    11'b00000111110: data <= 32'h39dbbcb8;
    11'b00000111111: data <= 32'h3769c0b4;
    11'b00001000000: data <= 32'h399fbee8;
    11'b00001000001: data <= 32'h37753817;
    11'b00001000010: data <= 32'hb8e23f34;
    11'b00001000011: data <= 32'hbda839a5;
    11'b00001000100: data <= 32'hbcd7bc64;
    11'b00001000101: data <= 32'hbb28bd4e;
    11'b00001000110: data <= 32'hbd42b1f6;
    11'b00001000111: data <= 32'hbe0e379d;
    11'b00001001000: data <= 32'hb28f3221;
    11'b00001001001: data <= 32'h3ec63359;
    11'b00001001010: data <= 32'h3f793c90;
    11'b00001001011: data <= 32'h9d7a3f34;
    11'b00001001100: data <= 32'hbe163d75;
    11'b00001001101: data <= 32'hbab638c3;
    11'b00001001110: data <= 32'h3ac73571;
    11'b00001001111: data <= 32'h3d43203b;
    11'b00001010000: data <= 32'h3873bc7c;
    11'b00001010001: data <= 32'h358fc015;
    11'b00001010010: data <= 32'h3ccdbcd8;
    11'b00001010011: data <= 32'h3e993a0b;
    11'b00001010100: data <= 32'h39dd3db5;
    11'b00001010101: data <= 32'hb89dac13;
    11'b00001010110: data <= 32'hbc65bec4;
    11'b00001010111: data <= 32'hbc9dbdd5;
    11'b00001011000: data <= 32'hbdc3b1e0;
    11'b00001011001: data <= 32'hbd96282e;
    11'b00001011010: data <= 32'hb2e4bafa;
    11'b00001011011: data <= 32'h3caabbe1;
    11'b00001011100: data <= 32'h3b58377e;
    11'b00001011101: data <= 32'hbabc3fce;
    11'b00001011110: data <= 32'hbf574001;
    11'b00001011111: data <= 32'hba7f3ca0;
    11'b00001100000: data <= 32'h391a38c2;
    11'b00001100001: data <= 32'h38793344;
    11'b00001100010: data <= 32'hb642b857;
    11'b00001100011: data <= 32'hada8bc5d;
    11'b00001100100: data <= 32'h3e8db575;
    11'b00001100101: data <= 32'h414d3c56;
    11'b00001100110: data <= 32'h3ea53d0a;
    11'b00001100111: data <= 32'hac43b269;
    11'b00001101000: data <= 32'hba79bd7a;
    11'b00001101001: data <= 32'hb960baed;
    11'b00001101010: data <= 32'hb9502508;
    11'b00001101011: data <= 32'hb981b8dc;
    11'b00001101100: data <= 32'ha83fc03e;
    11'b00001101101: data <= 32'h3a36c04f;
    11'b00001101110: data <= 32'h36a0b0ae;
    11'b00001101111: data <= 32'hbbbb3f10;
    11'b00001110000: data <= 32'hbe683f28;
    11'b00001110001: data <= 32'hba3e3999;
    11'b00001110010: data <= 32'haa7e317c;
    11'b00001110011: data <= 32'hb9ee348a;
    11'b00001110100: data <= 32'hbe822e15;
    11'b00001110101: data <= 32'hb953b469;
    11'b00001110110: data <= 32'h3ec93031;
    11'b00001110111: data <= 32'h41b13c73;
    11'b00001111000: data <= 32'h3e813d2a;
    11'b00001111001: data <= 32'hb16435ee;
    11'b00001111010: data <= 32'hb840b38b;
    11'b00001111011: data <= 32'h30da33bc;
    11'b00001111100: data <= 32'h359b3718;
    11'b00001111101: data <= 32'ha76cbbbc;
    11'b00001111110: data <= 32'h2d82c189;
    11'b00001111111: data <= 32'h39c9c124;
    11'b00010000000: data <= 32'h39d0b55b;
    11'b00010000001: data <= 32'hb11e3d84;
    11'b00010000010: data <= 32'hba323b79;
    11'b00010000011: data <= 32'hb8aeb596;
    11'b00010000100: data <= 32'hb97bb80e;
    11'b00010000101: data <= 32'hbf0e33cc;
    11'b00010000110: data <= 32'hc0d8361a;
    11'b00010000111: data <= 32'hbc3bb33c;
    11'b00010001000: data <= 32'h3d62b472;
    11'b00010001001: data <= 32'h405338ef;
    11'b00010001010: data <= 32'h39e93d4f;
    11'b00010001011: data <= 32'hb9c03cc7;
    11'b00010001100: data <= 32'hb62d3c05;
    11'b00010001101: data <= 32'h3a083cff;
    11'b00010001110: data <= 32'h3a773b3d;
    11'b00010001111: data <= 32'haa93ba52;
    11'b00010010000: data <= 32'hb071c0dd;
    11'b00010010001: data <= 32'h3b2cc00d;
    11'b00010010010: data <= 32'h3e6ca6c9;
    11'b00010010011: data <= 32'h3c733c19;
    11'b00010010100: data <= 32'h33be297f;
    11'b00010010101: data <= 32'hb2f3bcb0;
    11'b00010010110: data <= 32'hba4eba62;
    11'b00010010111: data <= 32'hbf753533;
    11'b00010011000: data <= 32'hc0a23399;
    11'b00010011001: data <= 32'hbc30bbe0;
    11'b00010011010: data <= 32'h3a9fbda4;
    11'b00010011011: data <= 32'h3c73b3d1;
    11'b00010011100: data <= 32'hb4d63cbc;
    11'b00010011101: data <= 32'hbcc63e90;
    11'b00010011110: data <= 32'hb4f23e2c;
    11'b00010011111: data <= 32'h3a853e3d;
    11'b00010100000: data <= 32'h35a43c9c;
    11'b00010100001: data <= 32'hbb3db270;
    11'b00010100010: data <= 32'hba15bd99;
    11'b00010100011: data <= 32'h3c11bbd3;
    11'b00010100100: data <= 32'h40c53761;
    11'b00010100101: data <= 32'h40093aa9;
    11'b00010100110: data <= 32'h3ad0b55c;
    11'b00010100111: data <= 32'h311bbc92;
    11'b00010101000: data <= 32'hb44db506;
    11'b00010101001: data <= 32'hbc19399d;
    11'b00010101010: data <= 32'hbddbacd6;
    11'b00010101011: data <= 32'hb9bfbff7;
    11'b00010101100: data <= 32'h36f0c11d;
    11'b00010101101: data <= 32'h3652bbfa;
    11'b00010101110: data <= 32'hb9b43ad5;
    11'b00010101111: data <= 32'hbc593d6c;
    11'b00010110000: data <= 32'haff63c26;
    11'b00010110001: data <= 32'h373e3c22;
    11'b00010110010: data <= 32'hb9853c5a;
    11'b00010110011: data <= 32'hc03b36df;
    11'b00010110100: data <= 32'hbe07b65d;
    11'b00010110101: data <= 32'h3b0bb34d;
    11'b00010110110: data <= 32'h40f33916;
    11'b00010110111: data <= 32'h3fca39e7;
    11'b00010111000: data <= 32'h398ead37;
    11'b00010111001: data <= 32'h35a8b473;
    11'b00010111010: data <= 32'h38633a19;
    11'b00010111011: data <= 32'h30d43d44;
    11'b00010111100: data <= 32'hb854b24e;
    11'b00010111101: data <= 32'hb6f6c101;
    11'b00010111110: data <= 32'h348fc1e6;
    11'b00010111111: data <= 32'h3677bcb7;
    11'b00011000000: data <= 32'hb1f13804;
    11'b00011000001: data <= 32'hb4dd37f2;
    11'b00011000010: data <= 32'h345bb0cb;
    11'b00011000011: data <= 32'h2db02f3c;
    11'b00011000100: data <= 32'hbe393b01;
    11'b00011000101: data <= 32'hc1cd3a3f;
    11'b00011000110: data <= 32'hbfc6ac0f;
    11'b00011000111: data <= 32'h381bb592;
    11'b00011001000: data <= 32'h3f14328c;
    11'b00011001001: data <= 32'h3b8a3897;
    11'b00011001010: data <= 32'hac73372c;
    11'b00011001011: data <= 32'h354a3a46;
    11'b00011001100: data <= 32'h3cc53f19;
    11'b00011001101: data <= 32'h3afb3f7c;
    11'b00011001110: data <= 32'hb4472a5a;
    11'b00011001111: data <= 32'hb88dc03f;
    11'b00011010000: data <= 32'h345ec09e;
    11'b00011010001: data <= 32'h3bcdb98d;
    11'b00011010010: data <= 32'h3b1a34d0;
    11'b00011010011: data <= 32'h39cbb6c2;
    11'b00011010100: data <= 32'h3a3abcde;
    11'b00011010101: data <= 32'h2ee3b7a2;
    11'b00011010110: data <= 32'hbe613ab6;
    11'b00011010111: data <= 32'hc1733a66;
    11'b00011011000: data <= 32'hbf32b814;
    11'b00011011001: data <= 32'h2fbfbd0c;
    11'b00011011010: data <= 32'h3993b954;
    11'b00011011011: data <= 32'hb5323420;
    11'b00011011100: data <= 32'hbabe39cb;
    11'b00011011101: data <= 32'h34423cf8;
    11'b00011011110: data <= 32'h3d8f4016;
    11'b00011011111: data <= 32'h39cf4014;
    11'b00011100000: data <= 32'hbb0f3861;
    11'b00011100001: data <= 32'hbcc1bc48;
    11'b00011100010: data <= 32'h326abc38;
    11'b00011100011: data <= 32'h3e2e2d6b;
    11'b00011100100: data <= 32'h3ec63446;
    11'b00011100101: data <= 32'h3d48bb4e;
    11'b00011100110: data <= 32'h3c88bdf8;
    11'b00011100111: data <= 32'h38a4b403;
    11'b00011101000: data <= 32'hb9d53cc7;
    11'b00011101001: data <= 32'hbec3397d;
    11'b00011101010: data <= 32'hbcc9bd1b;
    11'b00011101011: data <= 32'haec7c094;
    11'b00011101100: data <= 32'haf42bdb6;
    11'b00011101101: data <= 32'hbc24aed3;
    11'b00011101110: data <= 32'hbc0d36ff;
    11'b00011101111: data <= 32'h367c39a2;
    11'b00011110000: data <= 32'h3ce63d75;
    11'b00011110001: data <= 32'hab0f3eeb;
    11'b00011110010: data <= 32'hbfd23c0d;
    11'b00011110011: data <= 32'hbfd71fce;
    11'b00011110100: data <= 32'ha59ca1c4;
    11'b00011110101: data <= 32'h3e543872;
    11'b00011110110: data <= 32'h3e5333e4;
    11'b00011110111: data <= 32'h3c2dbac6;
    11'b00011111000: data <= 32'h3c80bb3d;
    11'b00011111001: data <= 32'h3cfd3959;
    11'b00011111010: data <= 32'h38143f5e;
    11'b00011111011: data <= 32'hb7bc3987;
    11'b00011111100: data <= 32'hb8cfbec5;
    11'b00011111101: data <= 32'hb0d5c143;
    11'b00011111110: data <= 32'hb46ebe1d;
    11'b00011111111: data <= 32'hba66b4ed;
    11'b00100000000: data <= 32'hb693b4c9;
    11'b00100000001: data <= 32'h3aaab850;
    11'b00100000010: data <= 32'h3c11319e;
    11'b00100000011: data <= 32'hba4b3ccc;
    11'b00100000100: data <= 32'hc15e3cf0;
    11'b00100000101: data <= 32'hc0b337f6;
    11'b00100000110: data <= 32'hb4b5318e;
    11'b00100000111: data <= 32'h3bb8355b;
    11'b00100001000: data <= 32'h38332c0e;
    11'b00100001001: data <= 32'h287fb7e9;
    11'b00100001010: data <= 32'h3a56a0b9;
    11'b00100001011: data <= 32'h3efb3e75;
    11'b00100001100: data <= 32'h3d7b40c5;
    11'b00100001101: data <= 32'h2eba3b30;
    11'b00100001110: data <= 32'hb7e1bd75;
    11'b00100001111: data <= 32'hb11abfc5;
    11'b00100010000: data <= 32'h2ec0ba9a;
    11'b00100010001: data <= 32'h2cdfb30b;
    11'b00100010010: data <= 32'h3852bc45;
    11'b00100010011: data <= 32'h3d6dbeec;
    11'b00100010100: data <= 32'h3c33b9e0;
    11'b00100010101: data <= 32'hbab73b1e;
    11'b00100010110: data <= 32'hc0ed3ce2;
    11'b00100010111: data <= 32'hc00c33bc;
    11'b00100011000: data <= 32'hb6dcb81c;
    11'b00100011001: data <= 32'h28bab709;
    11'b00100011010: data <= 32'hbadcb4a5;
    11'b00100011011: data <= 32'hbc3db481;
    11'b00100011100: data <= 32'h36e036cf;
    11'b00100011101: data <= 32'h3f863f62;
    11'b00100011110: data <= 32'h3da440d3;
    11'b00100011111: data <= 32'hb41e3cb8;
    11'b00100100000: data <= 32'hbbeab70d;
    11'b00100100001: data <= 32'hb46cb8a4;
    11'b00100100010: data <= 32'h38933453;
    11'b00100100011: data <= 32'h3a972bbd;
    11'b00100100100: data <= 32'h3c6abde3;
    11'b00100100101: data <= 32'h3e78c05f;
    11'b00100100110: data <= 32'h3d6dba47;
    11'b00100100111: data <= 32'had683c5c;
    11'b00100101000: data <= 32'hbd533c95;
    11'b00100101001: data <= 32'hbc77b649;
    11'b00100101010: data <= 32'hb55cbdcc;
    11'b00100101011: data <= 32'hb959bcaf;
    11'b00100101100: data <= 32'hbefab8d7;
    11'b00100101101: data <= 32'hbe1eb74e;
    11'b00100101110: data <= 32'h360ba670;
    11'b00100101111: data <= 32'h3ef43c56;
    11'b00100110000: data <= 32'h3a3e3f4a;
    11'b00100110001: data <= 32'hbcd33d53;
    11'b00100110010: data <= 32'hbee5382b;
    11'b00100110011: data <= 32'hb7c93917;
    11'b00100110100: data <= 32'h39583c41;
    11'b00100110101: data <= 32'h3a2b3445;
    11'b00100110110: data <= 32'h3a19bda2;
    11'b00100110111: data <= 32'h3d75bf0f;
    11'b00100111000: data <= 32'h3eeaa590;
    11'b00100111001: data <= 32'h3c223ec0;
    11'b00100111010: data <= 32'h29a53ca9;
    11'b00100111011: data <= 32'hb1c5ba8e;
    11'b00100111100: data <= 32'haf8bbf4b;
    11'b00100111101: data <= 32'hba83bce2;
    11'b00100111110: data <= 32'hbebfb8da;
    11'b00100111111: data <= 32'hbc78bb72;
    11'b00101000000: data <= 32'h39e5bc99;
    11'b00101000001: data <= 32'h3e40b436;
    11'b00101000010: data <= 32'h2d073b8c;
    11'b00101000011: data <= 32'hbfc33d0b;
    11'b00101000100: data <= 32'hc0293bc4;
    11'b00101000101: data <= 32'hb8d83c0b;
    11'b00101000110: data <= 32'h34563c47;
    11'b00101000111: data <= 32'hb1a831cd;
    11'b00101001000: data <= 32'hb648bc61;
    11'b00101001001: data <= 32'h3980bb78;
    11'b00101001010: data <= 32'h3fab3b3e;
    11'b00101001011: data <= 32'h3f56406b;
    11'b00101001100: data <= 32'h3aa43d10;
    11'b00101001101: data <= 32'h323ab955;
    11'b00101001110: data <= 32'h2033bceb;
    11'b00101001111: data <= 32'hb77bb63c;
    11'b00101010000: data <= 32'hbb40b222;
    11'b00101010001: data <= 32'hb2d1bd8b;
    11'b00101010010: data <= 32'h3cfec089;
    11'b00101010011: data <= 32'h3e1fbd82;
    11'b00101010100: data <= 32'haec9354b;
    11'b00101010101: data <= 32'hbf353c49;
    11'b00101010110: data <= 32'hbe9539ed;
    11'b00101010111: data <= 32'hb70f3723;
    11'b00101011000: data <= 32'hb5ab3606;
    11'b00101011001: data <= 32'hbdeab113;
    11'b00101011010: data <= 32'hbec6bad4;
    11'b00101011011: data <= 32'h9e1bb68b;
    11'b00101011100: data <= 32'h3f593cd5;
    11'b00101011101: data <= 32'h3f89404f;
    11'b00101011110: data <= 32'h38ed3d24;
    11'b00101011111: data <= 32'hb1caa6ee;
    11'b00101100000: data <= 32'had322a73;
    11'b00101100001: data <= 32'h91573b4a;
    11'b00101100010: data <= 32'haf013709;
    11'b00101100011: data <= 32'h368fbe2b;
    11'b00101100100: data <= 32'h3dd1c170;
    11'b00101100101: data <= 32'h3e79be64;
    11'b00101100110: data <= 32'h364035db;
    11'b00101100111: data <= 32'hba063b8c;
    11'b00101101000: data <= 32'hb8512fcf;
    11'b00101101001: data <= 32'h2266b7ff;
    11'b00101101010: data <= 32'hba4eb657;
    11'b00101101011: data <= 32'hc0b3b71e;
    11'b00101101100: data <= 32'hc0b6badd;
    11'b00101101101: data <= 32'hb44ab90f;
    11'b00101101110: data <= 32'h3e6e383f;
    11'b00101101111: data <= 32'h3d1b3d88;
    11'b00101110000: data <= 32'hb4ee3c50;
    11'b00101110001: data <= 32'hbb773933;
    11'b00101110010: data <= 32'hb4793cfa;
    11'b00101110011: data <= 32'h33093fac;
    11'b00101110100: data <= 32'h27d43b36;
    11'b00101110101: data <= 32'h30f4bd6d;
    11'b00101110110: data <= 32'h3c2ec0a4;
    11'b00101110111: data <= 32'h3e99bb22;
    11'b00101111000: data <= 32'h3ce03b9d;
    11'b00101111001: data <= 32'h38bd3ba7;
    11'b00101111010: data <= 32'h3904b63d;
    11'b00101111011: data <= 32'h3836bc20;
    11'b00101111100: data <= 32'hba33b846;
    11'b00101111101: data <= 32'hc0a1b525;
    11'b00101111110: data <= 32'hc011bc16;
    11'b00101111111: data <= 32'h2971bde4;
    11'b00110000000: data <= 32'h3db0ba3b;
    11'b00110000001: data <= 32'h38273436;
    11'b00110000010: data <= 32'hbcaa396b;
    11'b00110000011: data <= 32'hbd803b40;
    11'b00110000100: data <= 32'hb4eb3e8e;
    11'b00110000101: data <= 32'h2e0c401b;
    11'b00110000110: data <= 32'hb92c3b43;
    11'b00110000111: data <= 32'hbba2bc13;
    11'b00110001000: data <= 32'h3025bdd3;
    11'b00110001001: data <= 32'h3df1300f;
    11'b00110001010: data <= 32'h3f303e37;
    11'b00110001011: data <= 32'h3d983bf7;
    11'b00110001100: data <= 32'h3cadb77e;
    11'b00110001101: data <= 32'h3a5db982;
    11'b00110001110: data <= 32'hb61c33c5;
    11'b00110001111: data <= 32'hbe143518;
    11'b00110010000: data <= 32'hbc4abc77;
    11'b00110010001: data <= 32'h38fbc0b2;
    11'b00110010010: data <= 32'h3d6abfa4;
    11'b00110010011: data <= 32'h3090b868;
    11'b00110010100: data <= 32'hbd0934a9;
    11'b00110010101: data <= 32'hbc0538cc;
    11'b00110010110: data <= 32'h2bbd3c4d;
    11'b00110010111: data <= 32'hb1a83d5b;
    11'b00110011000: data <= 32'hbec83827;
    11'b00110011001: data <= 32'hc08aba12;
    11'b00110011010: data <= 32'hba5aba35;
    11'b00110011011: data <= 32'h3ca23920;
    11'b00110011100: data <= 32'h3ef33e4e;
    11'b00110011101: data <= 32'h3cc93ab8;
    11'b00110011110: data <= 32'h3a89b14a;
    11'b00110011111: data <= 32'h3983355b;
    11'b00110100000: data <= 32'h2e2b3e37;
    11'b00110100001: data <= 32'hb8cd3ccc;
    11'b00110100010: data <= 32'hb424bbe2;
    11'b00110100011: data <= 32'h3b5ac151;
    11'b00110100100: data <= 32'h3d33c04e;
    11'b00110100101: data <= 32'h3539b8b0;
    11'b00110100110: data <= 32'hb7733060;
    11'b00110100111: data <= 32'h2eada870;
    11'b00110101000: data <= 32'h3a3128c3;
    11'b00110101001: data <= 32'hb4b1366e;
    11'b00110101010: data <= 32'hc0cd3046;
    11'b00110101011: data <= 32'hc1edb941;
    11'b00110101100: data <= 32'hbcb1b9b9;
    11'b00110101101: data <= 32'h3ad332f9;
    11'b00110101110: data <= 32'h3c653a81;
    11'b00110101111: data <= 32'h328f3600;
    11'b00110110000: data <= 32'hac653196;
    11'b00110110001: data <= 32'h36463d5f;
    11'b00110110010: data <= 32'h36414135;
    11'b00110110011: data <= 32'hb2a93f4b;
    11'b00110110100: data <= 32'hb437b95f;
    11'b00110110101: data <= 32'h3850c06a;
    11'b00110110110: data <= 32'h3c58bd9b;
    11'b00110110111: data <= 32'h3a792e24;
    11'b00110111000: data <= 32'h396f338e;
    11'b00110111001: data <= 32'h3d4ab8c8;
    11'b00110111010: data <= 32'h3df7b9b7;
    11'b00110111011: data <= 32'hae7c2519;
    11'b00110111100: data <= 32'hc0953289;
    11'b00110111101: data <= 32'hc13db8d0;
    11'b00110111110: data <= 32'hba78bcda;
    11'b00110111111: data <= 32'h39d4bb08;
    11'b00111000000: data <= 32'h34dbb5c6;
    11'b00111000001: data <= 32'hbabfb43b;
    11'b00111000010: data <= 32'hb9f4329a;
    11'b00111000011: data <= 32'h34a43e95;
    11'b00111000100: data <= 32'h373f417a;
    11'b00111000101: data <= 32'hb86f3f4c;
    11'b00111000110: data <= 32'hbc98b5ca;
    11'b00111000111: data <= 32'hb6cdbd3d;
    11'b00111001000: data <= 32'h3948b303;
    11'b00111001001: data <= 32'h3c7d3b56;
    11'b00111001010: data <= 32'h3d7f35db;
    11'b00111001011: data <= 32'h3f91baa5;
    11'b00111001100: data <= 32'h3f3db97b;
    11'b00111001101: data <= 32'h34df3883;
    11'b00111001110: data <= 32'hbdd73b06;
    11'b00111001111: data <= 32'hbe13b6d6;
    11'b00111010000: data <= 32'ha78abf2d;
    11'b00111010001: data <= 32'h3a16bf86;
    11'b00111010010: data <= 32'hb25cbce7;
    11'b00111010011: data <= 32'hbcecba0d;
    11'b00111010100: data <= 32'hb8eab128;
    11'b00111010101: data <= 32'h395e3c28;
    11'b00111010110: data <= 32'h371e3fac;
    11'b00111010111: data <= 32'hbd2a3d0f;
    11'b00111011000: data <= 32'hc0a3b27c;
    11'b00111011001: data <= 32'hbdabb837;
    11'b00111011010: data <= 32'h319d3891;
    11'b00111011011: data <= 32'h3b9d3cbf;
    11'b00111011100: data <= 32'h3c7b3319;
    11'b00111011101: data <= 32'h3ddcba34;
    11'b00111011110: data <= 32'h3e4b24d5;
    11'b00111011111: data <= 32'h398b3edd;
    11'b00111100000: data <= 32'hb7553f5a;
    11'b00111100001: data <= 32'hb72cae0b;
    11'b00111100010: data <= 32'h382cbfc8;
    11'b00111100011: data <= 32'h39f6c01f;
    11'b00111100100: data <= 32'hb3c2bce3;
    11'b00111100101: data <= 32'hba12baa7;
    11'b00111100110: data <= 32'h3526b9d6;
    11'b00111100111: data <= 32'h3ddcac59;
    11'b00111101000: data <= 32'h387d39f6;
    11'b00111101001: data <= 32'hbf3138fe;
    11'b00111101010: data <= 32'hc1e1b149;
    11'b00111101011: data <= 32'hbf2cb436;
    11'b00111101100: data <= 32'haee13786;
    11'b00111101101: data <= 32'h358438eb;
    11'b00111101110: data <= 32'h2c4eb514;
    11'b00111101111: data <= 32'h35f1b981;
    11'b00111110000: data <= 32'h3c1e3a62;
    11'b00111110001: data <= 32'h3b39415e;
    11'b00111110010: data <= 32'h2f2340fc;
    11'b00111110011: data <= 32'hb0413413;
    11'b00111110100: data <= 32'h35a6bdf1;
    11'b00111110101: data <= 32'h3797bd01;
    11'b00111110110: data <= 32'ha58fb5d2;
    11'b00111110111: data <= 32'h3034b80f;
    11'b00111111000: data <= 32'h3dcebccb;
    11'b00111111001: data <= 32'h407dbbc9;
    11'b00111111010: data <= 32'h3ac02a3e;
    11'b00111111011: data <= 32'hbe8e375f;
    11'b00111111100: data <= 32'hc113ad02;
    11'b00111111101: data <= 32'hbd26b7ff;
    11'b00111111110: data <= 32'ha93eb5a0;
    11'b00111111111: data <= 32'hb5c5b757;
    11'b01000000000: data <= 32'hbc76bc2b;
    11'b01000000001: data <= 32'hb8dfba62;
    11'b01000000010: data <= 32'h39663c0b;
    11'b01000000011: data <= 32'h3bbb4188;
    11'b01000000100: data <= 32'h240340c9;
    11'b01000000101: data <= 32'hb9cd36aa;
    11'b01000000110: data <= 32'hb7e3b94e;
    11'b01000000111: data <= 32'haa7b2acf;
    11'b01000001000: data <= 32'h2ee439fd;
    11'b01000001001: data <= 32'h399baf50;
    11'b01000001010: data <= 32'h3fe1bd9e;
    11'b01000001011: data <= 32'h4103bcb7;
    11'b01000001100: data <= 32'h3c9b3498;
    11'b01000001101: data <= 32'hbae53bf1;
    11'b01000001110: data <= 32'hbd4f323a;
    11'b01000001111: data <= 32'hb382baeb;
    11'b01000010000: data <= 32'h341cbcc7;
    11'b01000010001: data <= 32'hba83bd1c;
    11'b01000010010: data <= 32'hbee3be1b;
    11'b01000010011: data <= 32'hba5dbc7f;
    11'b01000010100: data <= 32'h3b1936f1;
    11'b01000010101: data <= 32'h3c2d3f63;
    11'b01000010110: data <= 32'hb7c63e57;
    11'b01000010111: data <= 32'hbed33515;
    11'b01000011000: data <= 32'hbdc02b3c;
    11'b01000011001: data <= 32'hb88f3c32;
    11'b01000011010: data <= 32'had293d60;
    11'b01000011011: data <= 32'h3723abe7;
    11'b01000011100: data <= 32'h3dd9bdaa;
    11'b01000011101: data <= 32'h401eb9c0;
    11'b01000011110: data <= 32'h3d363ce5;
    11'b01000011111: data <= 32'h2c8e3f97;
    11'b01000100000: data <= 32'hac0b38c3;
    11'b01000100001: data <= 32'h3931bb8f;
    11'b01000100010: data <= 32'h3772bd5e;
    11'b01000100011: data <= 32'hbb36bcd6;
    11'b01000100100: data <= 32'hbdfdbdbd;
    11'b01000100101: data <= 32'hae42bdf4;
    11'b01000100110: data <= 32'h3e74b8da;
    11'b01000100111: data <= 32'h3d0037e8;
    11'b01000101000: data <= 32'hbb0038e0;
    11'b01000101001: data <= 32'hc0872ed7;
    11'b01000101010: data <= 32'hbf0d356f;
    11'b01000101011: data <= 32'hb9e63cc8;
    11'b01000101100: data <= 32'hb83b3c23;
    11'b01000101101: data <= 32'hb866b81b;
    11'b01000101110: data <= 32'h328bbdb6;
    11'b01000101111: data <= 32'h3cc1adf8;
    11'b01000110000: data <= 32'h3cfe4034;
    11'b01000110001: data <= 32'h39194108;
    11'b01000110010: data <= 32'h37ff3b09;
    11'b01000110011: data <= 32'h3a29b8bc;
    11'b01000110100: data <= 32'h34f5b894;
    11'b01000110101: data <= 32'hba3fb28e;
    11'b01000110110: data <= 32'hba50ba71;
    11'b01000110111: data <= 32'h3b53bec2;
    11'b01000111000: data <= 32'h40bbbdf5;
    11'b01000111001: data <= 32'h3e0fb727;
    11'b01000111010: data <= 32'hba2c302c;
    11'b01000111011: data <= 32'hbf8929b8;
    11'b01000111100: data <= 32'hbc88323b;
    11'b01000111101: data <= 32'hb65838a2;
    11'b01000111110: data <= 32'hbbd22ea2;
    11'b01000111111: data <= 32'hbeccbcde;
    11'b01001000000: data <= 32'hbc0fbe40;
    11'b01001000001: data <= 32'h37f23011;
    11'b01001000010: data <= 32'h3c814060;
    11'b01001000011: data <= 32'h38ef40a1;
    11'b01001000100: data <= 32'h30353a76;
    11'b01001000101: data <= 32'h2e3e99ee;
    11'b01001000110: data <= 32'hb20e3990;
    11'b01001000111: data <= 32'hb9ad3c8e;
    11'b01001001000: data <= 32'hb420abe4;
    11'b01001001001: data <= 32'h3db1beb8;
    11'b01001001010: data <= 32'h411cbf00;
    11'b01001001011: data <= 32'h3e8cb728;
    11'b01001001100: data <= 32'hb2443745;
    11'b01001001101: data <= 32'hb9a83466;
    11'b01001001110: data <= 32'h3081adb6;
    11'b01001001111: data <= 32'h3412b1e2;
    11'b01001010000: data <= 32'hbcc5b97e;
    11'b01001010001: data <= 32'hc0b0be9e;
    11'b01001010010: data <= 32'hbdcebf05;
    11'b01001010011: data <= 32'h376eb497;
    11'b01001010100: data <= 32'h3c8a3d31;
    11'b01001010101: data <= 32'h329b3d35;
    11'b01001010110: data <= 32'hb9de35cf;
    11'b01001010111: data <= 32'hba62377b;
    11'b01001011000: data <= 32'hb97b3edd;
    11'b01001011001: data <= 32'hba893ffb;
    11'b01001011010: data <= 32'hb6403453;
    11'b01001011011: data <= 32'h3b89be5b;
    11'b01001011100: data <= 32'h3fb4bd87;
    11'b01001011101: data <= 32'h3dd9357e;
    11'b01001011110: data <= 32'h37c93d23;
    11'b01001011111: data <= 32'h38963953;
    11'b01001100000: data <= 32'h3d2db272;
    11'b01001100001: data <= 32'h3a33b68f;
    11'b01001100010: data <= 32'hbc94b921;
    11'b01001100011: data <= 32'hc069bda8;
    11'b01001100100: data <= 32'hbb6cbf4e;
    11'b01001100101: data <= 32'h3c57bc57;
    11'b01001100110: data <= 32'h3d54ac16;
    11'b01001100111: data <= 32'hb1a12a98;
    11'b01001101000: data <= 32'hbd50b202;
    11'b01001101001: data <= 32'hbc9138ab;
    11'b01001101010: data <= 32'hb9eb3fc6;
    11'b01001101011: data <= 32'hbc103f8b;
    11'b01001101100: data <= 32'hbca7a92a;
    11'b01001101101: data <= 32'hb519be57;
    11'b01001101110: data <= 32'h3a45ba55;
    11'b01001101111: data <= 32'h3c313ce1;
    11'b01001110000: data <= 32'h3add3fa5;
    11'b01001110001: data <= 32'h3cd83af9;
    11'b01001110010: data <= 32'h3e94aa1c;
    11'b01001110011: data <= 32'h3a683137;
    11'b01001110100: data <= 32'hbbed35c2;
    11'b01001110101: data <= 32'hbe35b838;
    11'b01001110110: data <= 32'h2a7ebea7;
    11'b01001110111: data <= 32'h3f5abf03;
    11'b01001111000: data <= 32'h3e32bc4b;
    11'b01001111001: data <= 32'hb31db979;
    11'b01001111010: data <= 32'hbc74b79d;
    11'b01001111011: data <= 32'hb8283619;
    11'b01001111100: data <= 32'hb1503d96;
    11'b01001111101: data <= 32'hbc723c19;
    11'b01001111110: data <= 32'hc02cb9d4;
    11'b01001111111: data <= 32'hbe66bec7;
    11'b01010000000: data <= 32'hb201b77a;
    11'b01010000001: data <= 32'h393f3dc3;
    11'b01010000010: data <= 32'h39ff3ee7;
    11'b01010000011: data <= 32'h3b6038c8;
    11'b01010000100: data <= 32'h3c5032c7;
    11'b01010000101: data <= 32'h35763cd3;
    11'b01010000110: data <= 32'hbb473f0a;
    11'b01010000111: data <= 32'hbba93816;
    11'b01010001000: data <= 32'h3950bd5f;
    11'b01010001001: data <= 32'h4019bf94;
    11'b01010001010: data <= 32'h3e05bca3;
    11'b01010001011: data <= 32'h2b3fb80f;
    11'b01010001100: data <= 32'hb0e3b520;
    11'b01010001101: data <= 32'h3a702dd2;
    11'b01010001110: data <= 32'h3a4938d8;
    11'b01010001111: data <= 32'hbbec310a;
    11'b01010010000: data <= 32'hc12bbcc9;
    11'b01010010001: data <= 32'hc041bf09;
    11'b01010010010: data <= 32'hb682b8fa;
    11'b01010010011: data <= 32'h385e3a0a;
    11'b01010010100: data <= 32'h3531395e;
    11'b01010010101: data <= 32'h2ba9b099;
    11'b01010010110: data <= 32'h3074354a;
    11'b01010010111: data <= 32'hb203401e;
    11'b01010011000: data <= 32'hbb6e416b;
    11'b01010011001: data <= 32'hbafb3c46;
    11'b01010011010: data <= 32'h35f9bc59;
    11'b01010011011: data <= 32'h3d90bdf9;
    11'b01010011100: data <= 32'h3c30b653;
    11'b01010011101: data <= 32'h36253548;
    11'b01010011110: data <= 32'h3b972e26;
    11'b01010011111: data <= 32'h401dacf4;
    11'b01010100000: data <= 32'h3e44328e;
    11'b01010100001: data <= 32'hb9d62724;
    11'b01010100010: data <= 32'hc0c8bb92;
    11'b01010100011: data <= 32'hbe98be4c;
    11'b01010100100: data <= 32'h31cfbc4b;
    11'b01010100101: data <= 32'h3a01b6bb;
    11'b01010100110: data <= 32'hade6b975;
    11'b01010100111: data <= 32'hb95bbbe2;
    11'b01010101000: data <= 32'hb5c93220;
    11'b01010101001: data <= 32'hb40b406b;
    11'b01010101010: data <= 32'hbb444155;
    11'b01010101011: data <= 32'hbd443aaa;
    11'b01010101100: data <= 32'hb993bc3f;
    11'b01010101101: data <= 32'h30c7bb07;
    11'b01010101110: data <= 32'h352638a5;
    11'b01010101111: data <= 32'h376b3c60;
    11'b01010110000: data <= 32'h3df63548;
    11'b01010110001: data <= 32'h40fcae97;
    11'b01010110010: data <= 32'h3edc37a4;
    11'b01010110011: data <= 32'hb8243ab3;
    11'b01010110100: data <= 32'hbedc2797;
    11'b01010110101: data <= 32'hb8d0bc5d;
    11'b01010110110: data <= 32'h3c2fbdb0;
    11'b01010110111: data <= 32'h3c06bd44;
    11'b01010111000: data <= 32'hb477be17;
    11'b01010111001: data <= 32'hb9c8bdc9;
    11'b01010111010: data <= 32'h2c7faf2f;
    11'b01010111011: data <= 32'h36463e8c;
    11'b01010111100: data <= 32'hb9863f0f;
    11'b01010111101: data <= 32'hbfa02bcc;
    11'b01010111110: data <= 32'hbf66bcd9;
    11'b01010111111: data <= 32'hbb8db724;
    11'b01011000000: data <= 32'hb4ae3c25;
    11'b01011000001: data <= 32'h329f3c60;
    11'b01011000010: data <= 32'h3caa1f38;
    11'b01011000011: data <= 32'h3facb05b;
    11'b01011000100: data <= 32'h3cd43cbc;
    11'b01011000101: data <= 32'hb78e4032;
    11'b01011000110: data <= 32'hbc273ccd;
    11'b01011000111: data <= 32'h32fcb80f;
    11'b01011001000: data <= 32'h3dc3bd79;
    11'b01011001001: data <= 32'h3b7fbd6d;
    11'b01011001010: data <= 32'hb43ebd7b;
    11'b01011001011: data <= 32'hadd5bd27;
    11'b01011001100: data <= 32'h3cfdb624;
    11'b01011001101: data <= 32'h3dea3a46;
    11'b01011001110: data <= 32'hb46339c4;
    11'b01011001111: data <= 32'hc055b8ae;
    11'b01011010000: data <= 32'hc0a2bd1d;
    11'b01011010001: data <= 32'hbce2b5e4;
    11'b01011010010: data <= 32'hb7413958;
    11'b01011010011: data <= 32'hb356323c;
    11'b01011010100: data <= 32'h3414baeb;
    11'b01011010101: data <= 32'h3aa9b549;
    11'b01011010110: data <= 32'h38163f16;
    11'b01011010111: data <= 32'hb81e41f5;
    11'b01011011000: data <= 32'hba093f62;
    11'b01011011001: data <= 32'h3352b098;
    11'b01011011010: data <= 32'h3b93bb55;
    11'b01011011011: data <= 32'h35cab865;
    11'b01011011100: data <= 32'hb41bb6bf;
    11'b01011011101: data <= 32'h39c8b9ce;
    11'b01011011110: data <= 32'h40d8b81b;
    11'b01011011111: data <= 32'h40c132f4;
    11'b01011100000: data <= 32'h30c234e7;
    11'b01011100001: data <= 32'hbf87b818;
    11'b01011100010: data <= 32'hbf30bbfc;
    11'b01011100011: data <= 32'hb876b80c;
    11'b01011100100: data <= 32'hb053b2a3;
    11'b01011100101: data <= 32'hb8d5bc4b;
    11'b01011100110: data <= 32'hb8e2bf64;
    11'b01011100111: data <= 32'h2c4eb972;
    11'b01011101000: data <= 32'h341d3f28;
    11'b01011101001: data <= 32'hb6d941c8;
    11'b01011101010: data <= 32'hbb353e4c;
    11'b01011101011: data <= 32'hb843b214;
    11'b01011101100: data <= 32'hb266b559;
    11'b01011101101: data <= 32'hb82a3852;
    11'b01011101110: data <= 32'hb6e238ab;
    11'b01011101111: data <= 32'h3c61b4ba;
    11'b01011110000: data <= 32'h41a2b897;
    11'b01011110001: data <= 32'h410f32ea;
    11'b01011110010: data <= 32'h35673a6f;
    11'b01011110011: data <= 32'hbcdf35ad;
    11'b01011110100: data <= 32'hb939b5a6;
    11'b01011110101: data <= 32'h3830b88e;
    11'b01011110110: data <= 32'h350cbb38;
    11'b01011110111: data <= 32'hba64bf83;
    11'b01011111000: data <= 32'hbb47c0b7;
    11'b01011111001: data <= 32'h320ebc10;
    11'b01011111010: data <= 32'h3a313ccd;
    11'b01011111011: data <= 32'hab633fa0;
    11'b01011111100: data <= 32'hbcbf38ea;
    11'b01011111101: data <= 32'hbdd5b835;
    11'b01011111110: data <= 32'hbd082d8e;
    11'b01011111111: data <= 32'hbce93cdd;
    11'b01100000000: data <= 32'hba363b1e;
    11'b01100000001: data <= 32'h39d0b785;
    11'b01100000010: data <= 32'h4058b9ec;
    11'b01100000011: data <= 32'h3f7b38e8;
    11'b01100000100: data <= 32'h32f93f42;
    11'b01100000101: data <= 32'hb8813df2;
    11'b01100000110: data <= 32'h35d535c2;
    11'b01100000111: data <= 32'h3cdfb5e9;
    11'b01100001000: data <= 32'h36a5baeb;
    11'b01100001001: data <= 32'hbb24beae;
    11'b01100001010: data <= 32'hb8a9c02e;
    11'b01100001011: data <= 32'h3c66bc9e;
    11'b01100001100: data <= 32'h3f4135f1;
    11'b01100001101: data <= 32'h381b397a;
    11'b01100001110: data <= 32'hbd02b52f;
    11'b01100001111: data <= 32'hbf43ba3a;
    11'b01100010000: data <= 32'hbdfb33da;
    11'b01100010001: data <= 32'hbd523c91;
    11'b01100010010: data <= 32'hbc7d344c;
    11'b01100010011: data <= 32'hb15ebd20;
    11'b01100010100: data <= 32'h3b6fbc68;
    11'b01100010101: data <= 32'h3b273bbe;
    11'b01100010110: data <= 32'ha654411c;
    11'b01100010111: data <= 32'hb3334036;
    11'b01100011000: data <= 32'h394139bf;
    11'b01100011001: data <= 32'h3c0f29bc;
    11'b01100011010: data <= 32'had31ab94;
    11'b01100011011: data <= 32'hbc36b8af;
    11'b01100011100: data <= 32'ha719bd16;
    11'b01100011101: data <= 32'h4039bc51;
    11'b01100011110: data <= 32'h4164b337;
    11'b01100011111: data <= 32'h3bd8188a;
    11'b01100100000: data <= 32'hbb95b871;
    11'b01100100001: data <= 32'hbd1ab8d0;
    11'b01100100010: data <= 32'hb9bd344d;
    11'b01100100011: data <= 32'hba503858;
    11'b01100100100: data <= 32'hbd36ba87;
    11'b01100100101: data <= 32'hbc2fc083;
    11'b01100100110: data <= 32'hadb4be2a;
    11'b01100100111: data <= 32'h35303b4e;
    11'b01100101000: data <= 32'hac8c40db;
    11'b01100101001: data <= 32'hb3433ef8;
    11'b01100101010: data <= 32'h31dd37df;
    11'b01100101011: data <= 32'h2cb2374d;
    11'b01100101100: data <= 32'hbba93c23;
    11'b01100101101: data <= 32'hbd68393f;
    11'b01100101110: data <= 32'h332fb828;
    11'b01100101111: data <= 32'h40e3bbd3;
    11'b01100110000: data <= 32'h4190b591;
    11'b01100110001: data <= 32'h3c273296;
    11'b01100110010: data <= 32'hb6b72d47;
    11'b01100110011: data <= 32'hb010276a;
    11'b01100110100: data <= 32'h38a935ba;
    11'b01100110101: data <= 32'ha5572117;
    11'b01100110110: data <= 32'hbd41be29;
    11'b01100110111: data <= 32'hbdc4c174;
    11'b01100111000: data <= 32'hb432bf32;
    11'b01100111001: data <= 32'h38b036b5;
    11'b01100111010: data <= 32'h34433dba;
    11'b01100111011: data <= 32'hb58938aa;
    11'b01100111100: data <= 32'hb859b0c4;
    11'b01100111101: data <= 32'hbb173975;
    11'b01100111110: data <= 32'hbe9a3f25;
    11'b01100111111: data <= 32'hbeb53d05;
    11'b01101000000: data <= 32'hae18b6a2;
    11'b01101000001: data <= 32'h3f21bc56;
    11'b01101000010: data <= 32'h3fc9af96;
    11'b01101000011: data <= 32'h39183beb;
    11'b01101000100: data <= 32'h29143c61;
    11'b01101000101: data <= 32'h3b9c39fb;
    11'b01101000110: data <= 32'h3e4538b9;
    11'b01101000111: data <= 32'h361a29e9;
    11'b01101001000: data <= 32'hbd44bd3c;
    11'b01101001001: data <= 32'hbd18c0a1;
    11'b01101001010: data <= 32'h3667bec1;
    11'b01101001011: data <= 32'h3deeb333;
    11'b01101001100: data <= 32'h3ad13119;
    11'b01101001101: data <= 32'hb553b922;
    11'b01101001110: data <= 32'hbad9b9c7;
    11'b01101001111: data <= 32'hbc5e39c4;
    11'b01101010000: data <= 32'hbe943f6e;
    11'b01101010001: data <= 32'hbf493b31;
    11'b01101010010: data <= 32'hba99bc39;
    11'b01101010011: data <= 32'h37efbdd5;
    11'b01101010100: data <= 32'h39892fd9;
    11'b01101010101: data <= 32'h2bc13e92;
    11'b01101010110: data <= 32'h33683eb3;
    11'b01101010111: data <= 32'h3d823c24;
    11'b01101011000: data <= 32'h3e943adb;
    11'b01101011001: data <= 32'h2d6439bc;
    11'b01101011010: data <= 32'hbdeab1f2;
    11'b01101011011: data <= 32'hbad5bcee;
    11'b01101011100: data <= 32'h3d26bd1d;
    11'b01101011101: data <= 32'h40a1b93e;
    11'b01101011110: data <= 32'h3d22b929;
    11'b01101011111: data <= 32'hafa0bcad;
    11'b01101100000: data <= 32'hb6a0ba3a;
    11'b01101100001: data <= 32'hb47f39ce;
    11'b01101100010: data <= 32'hbaf03da1;
    11'b01101100011: data <= 32'hbeb6a7c8;
    11'b01101100100: data <= 32'hbe1abfdf;
    11'b01101100101: data <= 32'hb910bf8e;
    11'b01101100110: data <= 32'hb2062ebc;
    11'b01101100111: data <= 32'hb4103e4b;
    11'b01101101000: data <= 32'h31ee3d1f;
    11'b01101101001: data <= 32'h3c3c38d9;
    11'b01101101010: data <= 32'h3b1a3bc7;
    11'b01101101011: data <= 32'hb9b23e88;
    11'b01101101100: data <= 32'hbf283c9f;
    11'b01101101101: data <= 32'hb8e5b133;
    11'b01101101110: data <= 32'h3e92bb02;
    11'b01101101111: data <= 32'h40bfb9a0;
    11'b01101110000: data <= 32'h3cb4b8ca;
    11'b01101110001: data <= 32'h30d8b9fa;
    11'b01101110010: data <= 32'h388cb40b;
    11'b01101110011: data <= 32'h3c703ab3;
    11'b01101110100: data <= 32'h330b3b66;
    11'b01101110101: data <= 32'hbd73b9f1;
    11'b01101110110: data <= 32'hbf45c0d5;
    11'b01101110111: data <= 32'hbbb1c00c;
    11'b01101111000: data <= 32'hb189b1a6;
    11'b01101111001: data <= 32'hab1939cd;
    11'b01101111010: data <= 32'h2d9f28f8;
    11'b01101111011: data <= 32'h36a8b585;
    11'b01101111100: data <= 32'ha71f3ae3;
    11'b01101111101: data <= 32'hbd8c4084;
    11'b01101111110: data <= 32'hc0113fa0;
    11'b01101111111: data <= 32'hba253301;
    11'b01110000000: data <= 32'h3c6cba6d;
    11'b01110000001: data <= 32'h3ddcb7b9;
    11'b01110000010: data <= 32'h37b52cd8;
    11'b01110000011: data <= 32'h34673200;
    11'b01110000100: data <= 32'h3e073723;
    11'b01110000101: data <= 32'h407c3c1d;
    11'b01110000110: data <= 32'h3b653ac9;
    11'b01110000111: data <= 32'hbc95b8e9;
    11'b01110001000: data <= 32'hbe8cbfc8;
    11'b01110001001: data <= 32'hb6d1be98;
    11'b01110001010: data <= 32'h38e0b7f8;
    11'b01110001011: data <= 32'h37fbb674;
    11'b01110001100: data <= 32'h2dcbbd55;
    11'b01110001101: data <= 32'h2913bcf8;
    11'b01110001110: data <= 32'hb4ff3922;
    11'b01110001111: data <= 32'hbd5c4096;
    11'b01110010000: data <= 32'hbfcd3ec2;
    11'b01110010001: data <= 32'hbcccb45b;
    11'b01110010010: data <= 32'ha8b2bc7f;
    11'b01110010011: data <= 32'h2c4bb400;
    11'b01110010100: data <= 32'hb6ee39fe;
    11'b01110010101: data <= 32'h31aa3a8e;
    11'b01110010110: data <= 32'h3f8039b0;
    11'b01110010111: data <= 32'h40f13c74;
    11'b01110011000: data <= 32'h3a873d05;
    11'b01110011001: data <= 32'hbce535e9;
    11'b01110011010: data <= 32'hbcedb9d4;
    11'b01110011011: data <= 32'h3721bb27;
    11'b01110011100: data <= 32'h3dddb8eb;
    11'b01110011101: data <= 32'h3b5dbc86;
    11'b01110011110: data <= 32'h316dc00d;
    11'b01110011111: data <= 32'h3425be1b;
    11'b01110100000: data <= 32'h35e13836;
    11'b01110100001: data <= 32'hb7193f6d;
    11'b01110100010: data <= 32'hbde23a73;
    11'b01110100011: data <= 32'hbe4bbcb8;
    11'b01110100100: data <= 32'hbc4cbe35;
    11'b01110100101: data <= 32'hbbeab199;
    11'b01110100110: data <= 32'hbc123ade;
    11'b01110100111: data <= 32'ha7a9385e;
    11'b01110101000: data <= 32'h3e3f31e1;
    11'b01110101001: data <= 32'h3f273b53;
    11'b01110101010: data <= 32'h2b143f61;
    11'b01110101011: data <= 32'hbe1f3e6f;
    11'b01110101100: data <= 32'hbb753834;
    11'b01110101101: data <= 32'h3b80b1e3;
    11'b01110101110: data <= 32'h3e89b75a;
    11'b01110101111: data <= 32'h39ebbc50;
    11'b01110110000: data <= 32'h3126bed1;
    11'b01110110001: data <= 32'h3b70bc4c;
    11'b01110110010: data <= 32'h3e9938fd;
    11'b01110110011: data <= 32'h3aa13d5e;
    11'b01110110100: data <= 32'hba909e5c;
    11'b01110110101: data <= 32'hbe7dbee5;
    11'b01110110110: data <= 32'hbd87be8c;
    11'b01110110111: data <= 32'hbc69b2f2;
    11'b01110111000: data <= 32'hbb8134c9;
    11'b01110111001: data <= 32'hb13bb8b0;
    11'b01110111010: data <= 32'h3b40bb94;
    11'b01110111011: data <= 32'h3a763742;
    11'b01110111100: data <= 32'hb99e4064;
    11'b01110111101: data <= 32'hbeff40a6;
    11'b01110111110: data <= 32'hbb203c3f;
    11'b01110111111: data <= 32'h394d2b72;
    11'b01111000000: data <= 32'h3aafb172;
    11'b01111000001: data <= 32'hafd9b66e;
    11'b01111000010: data <= 32'hac59b9ec;
    11'b01111000011: data <= 32'h3e4eb500;
    11'b01111000100: data <= 32'h41793a79;
    11'b01111000101: data <= 32'h3ed83c70;
    11'b01111000110: data <= 32'hb624af1b;
    11'b01111000111: data <= 32'hbd55bd77;
    11'b01111001000: data <= 32'hbac7bc74;
    11'b01111001001: data <= 32'hb53db246;
    11'b01111001010: data <= 32'hb595b83c;
    11'b01111001011: data <= 32'hb0fbbf9f;
    11'b01111001100: data <= 32'h369cc015;
    11'b01111001101: data <= 32'h351ca7db;
    11'b01111001110: data <= 32'hba30402a;
    11'b01111001111: data <= 32'hbe2e4036;
    11'b01111010000: data <= 32'hbc0038e9;
    11'b01111010001: data <= 32'hb1c2b427;
    11'b01111010010: data <= 32'hb80a2baa;
    11'b01111010011: data <= 32'hbcff35b1;
    11'b01111010100: data <= 32'hb7802c1a;
    11'b01111010101: data <= 32'h3f092caa;
    11'b01111010110: data <= 32'h41ed3a73;
    11'b01111010111: data <= 32'h3eba3ce6;
    11'b01111011000: data <= 32'hb69e38a2;
    11'b01111011001: data <= 32'hbb55b2df;
    11'b01111011010: data <= 32'h2d5eb08b;
    11'b01111011011: data <= 32'h395924d4;
    11'b01111011100: data <= 32'h3218bc2b;
    11'b01111011101: data <= 32'hb03bc12f;
    11'b01111011110: data <= 32'h360fc0e3;
    11'b01111011111: data <= 32'h39bdb3cb;
    11'b01111100000: data <= 32'h2a033e70;
    11'b01111100001: data <= 32'hbad73cb8;
    11'b01111100010: data <= 32'hbc19b666;
    11'b01111100011: data <= 32'hbbd2ba5b;
    11'b01111100100: data <= 32'hbe3b3144;
    11'b01111100101: data <= 32'hbff53971;
    11'b01111100110: data <= 32'hba9d2b30;
    11'b01111100111: data <= 32'h3d86b5d2;
    11'b01111101000: data <= 32'h407f36a7;
    11'b01111101001: data <= 32'h3acc3ddb;
    11'b01111101010: data <= 32'hba773e3e;
    11'b01111101011: data <= 32'hb8d43c23;
    11'b01111101100: data <= 32'h3a0d3a13;
    11'b01111101101: data <= 32'h3c55360e;
    11'b01111101110: data <= 32'h2f4ebb24;
    11'b01111101111: data <= 32'hb4e5c082;
    11'b01111110000: data <= 32'h39acbfd6;
    11'b01111110001: data <= 32'h3eedad8c;
    11'b01111110010: data <= 32'h3d3d3c5b;
    11'b01111110011: data <= 32'h22ba32ec;
    11'b01111110100: data <= 32'hba92bcb0;
    11'b01111110101: data <= 32'hbca1bbf9;
    11'b01111110110: data <= 32'hbeaa3419;
    11'b01111110111: data <= 32'hbfb2370d;
    11'b01111111000: data <= 32'hbb83ba6e;
    11'b01111111001: data <= 32'h39bcbde7;
    11'b01111111010: data <= 32'h3c92b473;
    11'b01111111011: data <= 32'haf753e18;
    11'b01111111100: data <= 32'hbc9d403c;
    11'b01111111101: data <= 32'hb75a3e50;
    11'b01111111110: data <= 32'h3a373c43;
    11'b01111111111: data <= 32'h3875398f;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    