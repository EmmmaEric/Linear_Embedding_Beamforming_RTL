
module memory_rom_26(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3be7bcf5;
    11'b00000000001: data <= 32'h380bb9ac;
    11'b00000000010: data <= 32'hb91439c2;
    11'b00000000011: data <= 32'hbedf39ff;
    11'b00000000100: data <= 32'hbdaabbf3;
    11'b00000000101: data <= 32'had43c0b7;
    11'b00000000110: data <= 32'h369bbf19;
    11'b00000000111: data <= 32'hb81fb2cd;
    11'b00000001000: data <= 32'hbcb13970;
    11'b00000001001: data <= 32'hb45c3b2c;
    11'b00000001010: data <= 32'h3ad63d30;
    11'b00000001011: data <= 32'h32c23e89;
    11'b00000001100: data <= 32'hbe8d3c11;
    11'b00000001101: data <= 32'hc04bb04e;
    11'b00000001110: data <= 32'hb6c2b614;
    11'b00000001111: data <= 32'h3e62369a;
    11'b00000010000: data <= 32'h3ff73997;
    11'b00000010001: data <= 32'h3d17b292;
    11'b00000010010: data <= 32'h3b67ba67;
    11'b00000010011: data <= 32'h3bbf3361;
    11'b00000010100: data <= 32'h37073e5f;
    11'b00000010101: data <= 32'hb7e43c01;
    11'b00000010110: data <= 32'hb958bd6b;
    11'b00000010111: data <= 32'ha4ccc1b5;
    11'b00000011000: data <= 32'h325ac017;
    11'b00000011001: data <= 32'hb682b687;
    11'b00000011010: data <= 32'hb8a22fcd;
    11'b00000011011: data <= 32'h3591b1c3;
    11'b00000011100: data <= 32'h3b382e40;
    11'b00000011101: data <= 32'hb6e03b7d;
    11'b00000011110: data <= 32'hc1053c59;
    11'b00000011111: data <= 32'hc18135ad;
    11'b00000100000: data <= 32'hba06ada6;
    11'b00000100001: data <= 32'h3c7b3357;
    11'b00000100010: data <= 32'h3c6d35f5;
    11'b00000100011: data <= 32'h344cad88;
    11'b00000100100: data <= 32'h36b0a2fe;
    11'b00000100101: data <= 32'h3d1f3d38;
    11'b00000100110: data <= 32'h3d0d40c3;
    11'b00000100111: data <= 32'h32393d57;
    11'b00000101000: data <= 32'hb7d2bc7b;
    11'b00000101001: data <= 32'haf6fc0af;
    11'b00000101010: data <= 32'h362bbd87;
    11'b00000101011: data <= 32'h35c6b112;
    11'b00000101100: data <= 32'h37c2b6fd;
    11'b00000101101: data <= 32'h3c84bd3a;
    11'b00000101110: data <= 32'h3c75bb52;
    11'b00000101111: data <= 32'hb836381b;
    11'b00000110000: data <= 32'hc0ef3c6b;
    11'b00000110001: data <= 32'hc1063412;
    11'b00000110010: data <= 32'hba21b964;
    11'b00000110011: data <= 32'h3681b927;
    11'b00000110100: data <= 32'hb1dbb391;
    11'b00000110101: data <= 32'hbb6ead24;
    11'b00000110110: data <= 32'haea636d7;
    11'b00000110111: data <= 32'h3d8a3ed9;
    11'b00000111000: data <= 32'h3db04116;
    11'b00000111001: data <= 32'hac1a3e39;
    11'b00000111010: data <= 32'hbc40b641;
    11'b00000111011: data <= 32'hb79bbc62;
    11'b00000111100: data <= 32'h3917b24f;
    11'b00000111101: data <= 32'h3c623510;
    11'b00000111110: data <= 32'h3ce8b9f8;
    11'b00000111111: data <= 32'h3e45bf5f;
    11'b00001000000: data <= 32'h3dafbc55;
    11'b00001000001: data <= 32'h2c853a00;
    11'b00001000010: data <= 32'hbdd93cfa;
    11'b00001000011: data <= 32'hbe2cb141;
    11'b00001000100: data <= 32'hb783be5a;
    11'b00001000101: data <= 32'hb0ecbe41;
    11'b00001000110: data <= 32'hbc70ba27;
    11'b00001000111: data <= 32'hbe21b4f8;
    11'b00001001000: data <= 32'hb1b42e63;
    11'b00001001001: data <= 32'h3da23c56;
    11'b00001001010: data <= 32'h3bff3fb3;
    11'b00001001011: data <= 32'hbbd73e14;
    11'b00001001100: data <= 32'hbff8366e;
    11'b00001001101: data <= 32'hbb86300a;
    11'b00001001110: data <= 32'h390c39e6;
    11'b00001001111: data <= 32'h3c9338db;
    11'b00001010000: data <= 32'h3c21ba40;
    11'b00001010001: data <= 32'h3d4cbe6d;
    11'b00001010010: data <= 32'h3e8cb5f4;
    11'b00001010011: data <= 32'h3c123e1f;
    11'b00001010100: data <= 32'hae973e2d;
    11'b00001010101: data <= 32'hb770b72c;
    11'b00001010110: data <= 32'haf99c019;
    11'b00001010111: data <= 32'hb540bf29;
    11'b00001011000: data <= 32'hbcd1baa3;
    11'b00001011001: data <= 32'hbcc6b952;
    11'b00001011010: data <= 32'h353bbae7;
    11'b00001011011: data <= 32'h3e0bb395;
    11'b00001011100: data <= 32'h378c3b3b;
    11'b00001011101: data <= 32'hbf223d22;
    11'b00001011110: data <= 32'hc11e3a9b;
    11'b00001011111: data <= 32'hbcba38f2;
    11'b00001100000: data <= 32'h34ed3aaf;
    11'b00001100001: data <= 32'h35a236d1;
    11'b00001100010: data <= 32'had1eb9ba;
    11'b00001100011: data <= 32'h3815bbb3;
    11'b00001100100: data <= 32'h3e8d38d7;
    11'b00001100101: data <= 32'h3f064092;
    11'b00001100110: data <= 32'h3a3e3f53;
    11'b00001100111: data <= 32'h25a2b504;
    11'b00001101000: data <= 32'ha863be6c;
    11'b00001101001: data <= 32'hb1d5bc20;
    11'b00001101010: data <= 32'hb8cfb4cc;
    11'b00001101011: data <= 32'hb41bbb60;
    11'b00001101100: data <= 32'h3c4dbf91;
    11'b00001101101: data <= 32'h3eddbdc2;
    11'b00001101110: data <= 32'h353930d8;
    11'b00001101111: data <= 32'hbf253c53;
    11'b00001110000: data <= 32'hc07b39f9;
    11'b00001110001: data <= 32'hbb9b32df;
    11'b00001110010: data <= 32'hb00e2fe0;
    11'b00001110011: data <= 32'hbab4b07b;
    11'b00001110100: data <= 32'hbdd8b9de;
    11'b00001110101: data <= 32'hb5b2b828;
    11'b00001110110: data <= 32'h3df33c22;
    11'b00001110111: data <= 32'h3fa640c7;
    11'b00001111000: data <= 32'h39bb3f67;
    11'b00001111001: data <= 32'hb5ad315e;
    11'b00001111010: data <= 32'hb548b740;
    11'b00001111011: data <= 32'h26433543;
    11'b00001111100: data <= 32'h2dec3834;
    11'b00001111101: data <= 32'h37c0bb9e;
    11'b00001111110: data <= 32'h3de7c0cf;
    11'b00001111111: data <= 32'h3f7bbf3e;
    11'b00010000000: data <= 32'h39b630ed;
    11'b00010000001: data <= 32'hbaf33c82;
    11'b00010000010: data <= 32'hbc6d360e;
    11'b00010000011: data <= 32'hb4e8b8f8;
    11'b00010000100: data <= 32'hb649ba27;
    11'b00010000101: data <= 32'hbee7b936;
    11'b00010000110: data <= 32'hc08dbae3;
    11'b00010000111: data <= 32'hb99ab973;
    11'b00010001000: data <= 32'h3d8637c5;
    11'b00010001001: data <= 32'h3e263e80;
    11'b00010001010: data <= 32'hadd83dee;
    11'b00010001011: data <= 32'hbce9394c;
    11'b00010001100: data <= 32'hba4139c1;
    11'b00010001101: data <= 32'h2ce43df0;
    11'b00010001110: data <= 32'h342b3c7c;
    11'b00010001111: data <= 32'h35c5ba8f;
    11'b00010010000: data <= 32'h3c73c069;
    11'b00010010001: data <= 32'h3f22bcef;
    11'b00010010010: data <= 32'h3d7b3ac3;
    11'b00010010011: data <= 32'h36f23da4;
    11'b00010010100: data <= 32'h325b2cb0;
    11'b00010010101: data <= 32'h3610bca2;
    11'b00010010110: data <= 32'hb5d2bc38;
    11'b00010010111: data <= 32'hbf63b8f8;
    11'b00010011000: data <= 32'hc031bba2;
    11'b00010011001: data <= 32'hb522bd7c;
    11'b00010011010: data <= 32'h3dd2ba30;
    11'b00010011011: data <= 32'h3c0e360f;
    11'b00010011100: data <= 32'hbb753b1e;
    11'b00010011101: data <= 32'hbf5b3acd;
    11'b00010011110: data <= 32'hbbb03ce9;
    11'b00010011111: data <= 32'ha8203f12;
    11'b00010100000: data <= 32'hb4963c6e;
    11'b00010100001: data <= 32'hb980b9a3;
    11'b00010100010: data <= 32'h2d62be55;
    11'b00010100011: data <= 32'h3dacb414;
    11'b00010100100: data <= 32'h3f643e85;
    11'b00010100101: data <= 32'h3d4b3ea4;
    11'b00010100110: data <= 32'h3b2b2930;
    11'b00010100111: data <= 32'h396dbb69;
    11'b00010101000: data <= 32'hb073b5c9;
    11'b00010101001: data <= 32'hbd1b2e9a;
    11'b00010101010: data <= 32'hbcc5bad2;
    11'b00010101011: data <= 32'h3700c040;
    11'b00010101100: data <= 32'h3e91bfe4;
    11'b00010101101: data <= 32'h39f5b8d9;
    11'b00010101110: data <= 32'hbc7436cd;
    11'b00010101111: data <= 32'hbe593940;
    11'b00010110000: data <= 32'hb87b3ae4;
    11'b00010110001: data <= 32'hb01d3c7e;
    11'b00010110010: data <= 32'hbcce3878;
    11'b00010110011: data <= 32'hc01eb9b7;
    11'b00010110100: data <= 32'hbc1ebc39;
    11'b00010110101: data <= 32'h3bb83524;
    11'b00010110110: data <= 32'h3f683f36;
    11'b00010110111: data <= 32'h3d303e29;
    11'b00010111000: data <= 32'h390232d2;
    11'b00010111001: data <= 32'h3700a94c;
    11'b00010111010: data <= 32'h2ceb3bdf;
    11'b00010111011: data <= 32'hb8413cbc;
    11'b00010111100: data <= 32'hb55fb863;
    11'b00010111101: data <= 32'h3b47c0e8;
    11'b00010111110: data <= 32'h3ec4c0c2;
    11'b00010111111: data <= 32'h3adfb9fb;
    11'b00011000000: data <= 32'hb73435eb;
    11'b00011000001: data <= 32'hb798343d;
    11'b00011000010: data <= 32'h356813ca;
    11'b00011000011: data <= 32'ha94830ca;
    11'b00011000100: data <= 32'hbf84a5b1;
    11'b00011000101: data <= 32'hc1d1ba2d;
    11'b00011000110: data <= 32'hbe38bbe1;
    11'b00011000111: data <= 32'h39a8223b;
    11'b00011001000: data <= 32'h3db73c48;
    11'b00011001001: data <= 32'h37be3b6f;
    11'b00011001010: data <= 32'hb4ac358c;
    11'b00011001011: data <= 32'haca33b3d;
    11'b00011001100: data <= 32'h3174405a;
    11'b00011001101: data <= 32'hb18a3ffa;
    11'b00011001110: data <= 32'hb3a2b2e5;
    11'b00011001111: data <= 32'h38bfc05c;
    11'b00011010000: data <= 32'h3d89bf3f;
    11'b00011010001: data <= 32'h3ca3aa65;
    11'b00011010010: data <= 32'h38ec3984;
    11'b00011010011: data <= 32'h3af2ac18;
    11'b00011010100: data <= 32'h3d13b97f;
    11'b00011010101: data <= 32'h338bb55e;
    11'b00011010110: data <= 32'hbf97aafa;
    11'b00011010111: data <= 32'hc180b96b;
    11'b00011011000: data <= 32'hbcd6bd58;
    11'b00011011001: data <= 32'h3a4bbc04;
    11'b00011011010: data <= 32'h3b1ab2b9;
    11'b00011011011: data <= 32'hb79a2c5e;
    11'b00011011100: data <= 32'hbc5233da;
    11'b00011011101: data <= 32'hb53a3d22;
    11'b00011011110: data <= 32'h32d040fe;
    11'b00011011111: data <= 32'hb687401f;
    11'b00011100000: data <= 32'hbc2cac32;
    11'b00011100001: data <= 32'hb75abe24;
    11'b00011100010: data <= 32'h39eeb9f0;
    11'b00011100011: data <= 32'h3d433b17;
    11'b00011100100: data <= 32'h3d673c16;
    11'b00011100101: data <= 32'h3e77b2cf;
    11'b00011100110: data <= 32'h3ecbb9e3;
    11'b00011100111: data <= 32'h38562f87;
    11'b00011101000: data <= 32'hbd2e396e;
    11'b00011101001: data <= 32'hbf20b4d6;
    11'b00011101010: data <= 32'hb53fbf00;
    11'b00011101011: data <= 32'h3c38c00f;
    11'b00011101100: data <= 32'h3842bd08;
    11'b00011101101: data <= 32'hbb3fb899;
    11'b00011101110: data <= 32'hbc40ad3c;
    11'b00011101111: data <= 32'h2c183af5;
    11'b00011110000: data <= 32'h35f83f40;
    11'b00011110001: data <= 32'hbbd23db2;
    11'b00011110010: data <= 32'hc073b0c1;
    11'b00011110011: data <= 32'hbe93bb90;
    11'b00011110100: data <= 32'h2c472af6;
    11'b00011110101: data <= 32'h3c893d27;
    11'b00011110110: data <= 32'h3d083b76;
    11'b00011110111: data <= 32'h3d56b459;
    11'b00011111000: data <= 32'h3da8b21f;
    11'b00011111001: data <= 32'h39a43d0f;
    11'b00011111010: data <= 32'hb8063f54;
    11'b00011111011: data <= 32'hb9dc3415;
    11'b00011111100: data <= 32'h35ddbf63;
    11'b00011111101: data <= 32'h3ca2c0b3;
    11'b00011111110: data <= 32'h371dbda8;
    11'b00011111111: data <= 32'hb892b91d;
    11'b00100000000: data <= 32'hb105b743;
    11'b00100000001: data <= 32'h3c1fa796;
    11'b00100000010: data <= 32'h39de3968;
    11'b00100000011: data <= 32'hbd8e3910;
    11'b00100000100: data <= 32'hc1f1b47a;
    11'b00100000101: data <= 32'hc06bb9a2;
    11'b00100000110: data <= 32'hb4182b99;
    11'b00100000111: data <= 32'h39803a2d;
    11'b00100001000: data <= 32'h367d3440;
    11'b00100001001: data <= 32'h348ab6b7;
    11'b00100001010: data <= 32'h39b93767;
    11'b00100001011: data <= 32'h39b340ad;
    11'b00100001100: data <= 32'h9eab4169;
    11'b00100001101: data <= 32'hb56b39a8;
    11'b00100001110: data <= 32'h346fbe02;
    11'b00100001111: data <= 32'h3a85bef2;
    11'b00100010000: data <= 32'h3776b8ed;
    11'b00100010001: data <= 32'h31eab13a;
    11'b00100010010: data <= 32'h3c39b992;
    11'b00100010011: data <= 32'h4017baa1;
    11'b00100010100: data <= 32'h3cb8ad85;
    11'b00100010101: data <= 32'hbd2735d1;
    11'b00100010110: data <= 32'hc185b1ab;
    11'b00100010111: data <= 32'hbf2eba53;
    11'b00100011000: data <= 32'habd2b91a;
    11'b00100011001: data <= 32'h330ab5db;
    11'b00100011010: data <= 32'hb929b98f;
    11'b00100011011: data <= 32'hba13b9e0;
    11'b00100011100: data <= 32'h33013972;
    11'b00100011101: data <= 32'h39dd4132;
    11'b00100011110: data <= 32'h8958417b;
    11'b00100011111: data <= 32'hba903a52;
    11'b00100100000: data <= 32'hb8efbb42;
    11'b00100100001: data <= 32'h2c79b8b1;
    11'b00100100010: data <= 32'h35ff386b;
    11'b00100100011: data <= 32'h39c6368d;
    11'b00100100100: data <= 32'h3ef6ba62;
    11'b00100100101: data <= 32'h40f7bc5e;
    11'b00100100110: data <= 32'h3de529c2;
    11'b00100100111: data <= 32'hb9a43b5a;
    11'b00100101000: data <= 32'hbedf34a8;
    11'b00100101001: data <= 32'hb9a8bb80;
    11'b00100101010: data <= 32'h3702bdba;
    11'b00100101011: data <= 32'hac8bbd60;
    11'b00100101100: data <= 32'hbd0fbd89;
    11'b00100101101: data <= 32'hbc3cbc6f;
    11'b00100101110: data <= 32'h369533fe;
    11'b00100101111: data <= 32'h3bbe3f66;
    11'b00100110000: data <= 32'hb4b83fb6;
    11'b00100110001: data <= 32'hbefb37ee;
    11'b00100110010: data <= 32'hbee3b63c;
    11'b00100110011: data <= 32'hb977360d;
    11'b00100110100: data <= 32'h2da73d11;
    11'b00100110101: data <= 32'h3893384f;
    11'b00100110110: data <= 32'h3d99bb41;
    11'b00100110111: data <= 32'h401fba8b;
    11'b00100111000: data <= 32'h3dd43b55;
    11'b00100111001: data <= 32'h23223fec;
    11'b00100111010: data <= 32'hb8263b9a;
    11'b00100111011: data <= 32'h34adbb05;
    11'b00100111100: data <= 32'h3a38be9f;
    11'b00100111101: data <= 32'hb1cebdcc;
    11'b00100111110: data <= 32'hbcc4bd6e;
    11'b00100111111: data <= 32'hb712bd60;
    11'b00101000000: data <= 32'h3d16b8b2;
    11'b00101000001: data <= 32'h3dc438a2;
    11'b00101000010: data <= 32'hb8133abf;
    11'b00101000011: data <= 32'hc0b82f58;
    11'b00101000100: data <= 32'hc07bb0e6;
    11'b00101000101: data <= 32'hbbb4390e;
    11'b00101000110: data <= 32'hb4683c35;
    11'b00101000111: data <= 32'hb39e99c3;
    11'b00101001000: data <= 32'h336cbcad;
    11'b00101001001: data <= 32'h3c5bb63a;
    11'b00101001010: data <= 32'h3cd73f51;
    11'b00101001011: data <= 32'h37b841a0;
    11'b00101001100: data <= 32'h2f133d9f;
    11'b00101001101: data <= 32'h3827b875;
    11'b00101001110: data <= 32'h38b0bc39;
    11'b00101001111: data <= 32'hb440b861;
    11'b00101010000: data <= 32'hb970b919;
    11'b00101010001: data <= 32'h38abbd5e;
    11'b00101010010: data <= 32'h407ebd5d;
    11'b00101010011: data <= 32'h3fbab672;
    11'b00101010100: data <= 32'hb60f33e1;
    11'b00101010101: data <= 32'hc044287c;
    11'b00101010110: data <= 32'hbef6b0db;
    11'b00101010111: data <= 32'hb8813223;
    11'b00101011000: data <= 32'hb82d300b;
    11'b00101011001: data <= 32'hbcf3bb5d;
    11'b00101011010: data <= 32'hbc10be40;
    11'b00101011011: data <= 32'h3425b40a;
    11'b00101011100: data <= 32'h3c134017;
    11'b00101011101: data <= 32'h386a418d;
    11'b00101011110: data <= 32'haef63d4f;
    11'b00101011111: data <= 32'hb05eb0c2;
    11'b00101100000: data <= 32'haeb929d9;
    11'b00101100001: data <= 32'hb7643a7d;
    11'b00101100010: data <= 32'hb4503447;
    11'b00101100011: data <= 32'h3ccdbcd5;
    11'b00101100100: data <= 32'h4143be90;
    11'b00101100101: data <= 32'h403bb845;
    11'b00101100110: data <= 32'h2bda384b;
    11'b00101100111: data <= 32'hbc8336d8;
    11'b00101101000: data <= 32'hb79cb1c9;
    11'b00101101001: data <= 32'h3422b6fd;
    11'b00101101010: data <= 32'hb885ba14;
    11'b00101101011: data <= 32'hbf7dbe4f;
    11'b00101101100: data <= 32'hbe4cbf84;
    11'b00101101101: data <= 32'h312ab8b4;
    11'b00101101110: data <= 32'h3c983d4a;
    11'b00101101111: data <= 32'h35fb3f3a;
    11'b00101110000: data <= 32'hbab539d6;
    11'b00101110001: data <= 32'hbc7f2fa2;
    11'b00101110010: data <= 32'hbab83c0a;
    11'b00101110011: data <= 32'hb9f03f20;
    11'b00101110100: data <= 32'hb60039ad;
    11'b00101110101: data <= 32'h3afabcb8;
    11'b00101110110: data <= 32'h4027bde5;
    11'b00101110111: data <= 32'h3f4d2fbf;
    11'b00101111000: data <= 32'h38523dd0;
    11'b00101111001: data <= 32'h2be43c4a;
    11'b00101111010: data <= 32'h3a38ad4e;
    11'b00101111011: data <= 32'h3b73b93c;
    11'b00101111100: data <= 32'hb80dbae4;
    11'b00101111101: data <= 32'hbf8fbdc9;
    11'b00101111110: data <= 32'hbcc3bf8a;
    11'b00101111111: data <= 32'h3ac6bcd2;
    11'b00110000000: data <= 32'h3e682c43;
    11'b00110000001: data <= 32'h335d3794;
    11'b00110000010: data <= 32'hbd9a0e6f;
    11'b00110000011: data <= 32'hbe7d310d;
    11'b00110000100: data <= 32'hbc2e3d5c;
    11'b00110000101: data <= 32'hbb6c3f43;
    11'b00110000110: data <= 32'hbbfb35fd;
    11'b00110000111: data <= 32'hb47bbda1;
    11'b00110001000: data <= 32'h3af7bc8b;
    11'b00110001001: data <= 32'h3ce63b8a;
    11'b00110001010: data <= 32'h3a4d407e;
    11'b00110001011: data <= 32'h3a043dec;
    11'b00110001100: data <= 32'h3d122f47;
    11'b00110001101: data <= 32'h3bd9b27e;
    11'b00110001110: data <= 32'hb844267d;
    11'b00110001111: data <= 32'hbdecb819;
    11'b00110010000: data <= 32'hb4a0be27;
    11'b00110010001: data <= 32'h3f12bee6;
    11'b00110010010: data <= 32'h4023bbb4;
    11'b00110010011: data <= 32'h349fb666;
    11'b00110010100: data <= 32'hbd1db5b9;
    11'b00110010101: data <= 32'hbc882c9e;
    11'b00110010110: data <= 32'hb7553c07;
    11'b00110010111: data <= 32'hbad43c2c;
    11'b00110011000: data <= 32'hbf0cb777;
    11'b00110011001: data <= 32'hbe42bf2c;
    11'b00110011010: data <= 32'hb3d6bbca;
    11'b00110011011: data <= 32'h39c33ce6;
    11'b00110011100: data <= 32'h39e34070;
    11'b00110011101: data <= 32'h391a3cfe;
    11'b00110011110: data <= 32'h3a5f3397;
    11'b00110011111: data <= 32'h36513967;
    11'b00110100000: data <= 32'hb9d33da7;
    11'b00110100001: data <= 32'hbc56396f;
    11'b00110100010: data <= 32'h35b0bc42;
    11'b00110100011: data <= 32'h4051bf7b;
    11'b00110100100: data <= 32'h4043bcc5;
    11'b00110100101: data <= 32'h37cab530;
    11'b00110100110: data <= 32'hb7a6aed2;
    11'b00110100111: data <= 32'h30fd28ad;
    11'b00110101000: data <= 32'h392836c8;
    11'b00110101001: data <= 32'hb8553151;
    11'b00110101010: data <= 32'hc06ebc82;
    11'b00110101011: data <= 32'hc06ec00d;
    11'b00110101100: data <= 32'hb8afbc75;
    11'b00110101101: data <= 32'h39543970;
    11'b00110101110: data <= 32'h38453ceb;
    11'b00110101111: data <= 32'ha5ce361c;
    11'b00110110000: data <= 32'hb0a730b9;
    11'b00110110001: data <= 32'hb5613dc5;
    11'b00110110010: data <= 32'hbbaf40f0;
    11'b00110110011: data <= 32'hbc2e3d8f;
    11'b00110110100: data <= 32'h31b8ba77;
    11'b00110110101: data <= 32'h3e5fbe9c;
    11'b00110110110: data <= 32'h3e63b8f9;
    11'b00110110111: data <= 32'h38f13814;
    11'b00110111000: data <= 32'h380f3824;
    11'b00110111001: data <= 32'h3df92f3b;
    11'b00110111010: data <= 32'h3e6e2f0d;
    11'b00110111011: data <= 32'hb2dcab8a;
    11'b00110111100: data <= 32'hc04fbbfa;
    11'b00110111101: data <= 32'hbfb2bf47;
    11'b00110111110: data <= 32'ha4cabd9f;
    11'b00110111111: data <= 32'h3c4bb5f1;
    11'b00111000000: data <= 32'h3620b1e3;
    11'b00111000001: data <= 32'hb91ab93e;
    11'b00111000010: data <= 32'hb9e6af90;
    11'b00111000011: data <= 32'hb86e3eab;
    11'b00111000100: data <= 32'hbbca4135;
    11'b00111000101: data <= 32'hbd7f3cd8;
    11'b00111000110: data <= 32'hba30bba6;
    11'b00111000111: data <= 32'h34febd3e;
    11'b00111001000: data <= 32'h397132f7;
    11'b00111001001: data <= 32'h38423d77;
    11'b00111001010: data <= 32'h3c463b92;
    11'b00111001011: data <= 32'h402f31c0;
    11'b00111001100: data <= 32'h3f6a34f4;
    11'b00111001101: data <= 32'hafce391d;
    11'b00111001110: data <= 32'hbef096ef;
    11'b00111001111: data <= 32'hbc20bca6;
    11'b00111010000: data <= 32'h3b78be4d;
    11'b00111010001: data <= 32'h3e3ebd03;
    11'b00111010010: data <= 32'h3598bcb2;
    11'b00111010011: data <= 32'hb9ccbd00;
    11'b00111010100: data <= 32'hb6bfb5e3;
    11'b00111010101: data <= 32'h2d063d3c;
    11'b00111010110: data <= 32'hb8dd3f77;
    11'b00111010111: data <= 32'hbf2535ef;
    11'b00111011000: data <= 32'hbf95bd6e;
    11'b00111011001: data <= 32'hbb67bc59;
    11'b00111011010: data <= 32'hae683956;
    11'b00111011011: data <= 32'h344f3dfc;
    11'b00111011100: data <= 32'h3b4c397d;
    11'b00111011101: data <= 32'h3eb62936;
    11'b00111011110: data <= 32'h3d3a3ac8;
    11'b00111011111: data <= 32'hb5173f6e;
    11'b00111100000: data <= 32'hbd333d40;
    11'b00111100001: data <= 32'hb41cb623;
    11'b00111100010: data <= 32'h3dddbddc;
    11'b00111100011: data <= 32'h3e77bdad;
    11'b00111100100: data <= 32'h3522bcb8;
    11'b00111100101: data <= 32'hb3c3bc56;
    11'b00111100110: data <= 32'h3991b6d9;
    11'b00111100111: data <= 32'h3d33399f;
    11'b00111101000: data <= 32'h26e23b26;
    11'b00111101001: data <= 32'hbfccb6a1;
    11'b00111101010: data <= 32'hc0edbe69;
    11'b00111101011: data <= 32'hbd79bc28;
    11'b00111101100: data <= 32'hb4a536a2;
    11'b00111101101: data <= 32'h1e07396a;
    11'b00111101110: data <= 32'h337ab4a2;
    11'b00111101111: data <= 32'h3967b607;
    11'b00111110000: data <= 32'h37923d34;
    11'b00111110001: data <= 32'hb89e41a1;
    11'b00111110010: data <= 32'hbc72404a;
    11'b00111110011: data <= 32'hb1732b91;
    11'b00111110100: data <= 32'h3c49bc91;
    11'b00111110101: data <= 32'h3be7ba9d;
    11'b00111110110: data <= 32'h302bb515;
    11'b00111110111: data <= 32'h36adb633;
    11'b00111111000: data <= 32'h3fb1b517;
    11'b00111111001: data <= 32'h40cd346d;
    11'b00111111010: data <= 32'h38b236fa;
    11'b00111111011: data <= 32'hbef3b74a;
    11'b00111111100: data <= 32'hc048bd4e;
    11'b00111111101: data <= 32'hba71bc1b;
    11'b00111111110: data <= 32'h30d4b4ee;
    11'b00111111111: data <= 32'haf8eb8f3;
    11'b01000000000: data <= 32'hb76dbdea;
    11'b01000000001: data <= 32'haf82bb53;
    11'b01000000010: data <= 32'h2d6f3d53;
    11'b01000000011: data <= 32'hb86641d1;
    11'b01000000100: data <= 32'hbca84000;
    11'b01000000101: data <= 32'hba64acf3;
    11'b01000000110: data <= 32'had56ba75;
    11'b01000000111: data <= 32'had862cda;
    11'b01000001000: data <= 32'hb42939a9;
    11'b01000001001: data <= 32'h39fc328f;
    11'b01000001010: data <= 32'h40f2b438;
    11'b01000001011: data <= 32'h416f338a;
    11'b01000001100: data <= 32'h39ee3a93;
    11'b01000001101: data <= 32'hbd2f3671;
    11'b01000001110: data <= 32'hbccab81f;
    11'b01000001111: data <= 32'h348cbaf9;
    11'b01000010000: data <= 32'h3a52bb6e;
    11'b01000010001: data <= 32'hb085be39;
    11'b01000010010: data <= 32'hba0ac05b;
    11'b01000010011: data <= 32'hae2ebd20;
    11'b01000010100: data <= 32'h388c3b58;
    11'b01000010101: data <= 32'haa144040;
    11'b01000010110: data <= 32'hbcfc3c39;
    11'b01000010111: data <= 32'hbe8db8e1;
    11'b01000011000: data <= 32'hbd0bb8db;
    11'b01000011001: data <= 32'hbc033992;
    11'b01000011010: data <= 32'hb9903c73;
    11'b01000011011: data <= 32'h37fa2eba;
    11'b01000011100: data <= 32'h400bb81e;
    11'b01000011101: data <= 32'h40343738;
    11'b01000011110: data <= 32'h37183efa;
    11'b01000011111: data <= 32'hbb1a3e98;
    11'b01000100000: data <= 32'hb47536cc;
    11'b01000100001: data <= 32'h3c4bb84d;
    11'b01000100010: data <= 32'h3c10bbb5;
    11'b01000100011: data <= 32'hb40fbe1d;
    11'b01000100100: data <= 32'hb89dbff1;
    11'b01000100101: data <= 32'h39c2bd1e;
    11'b01000100110: data <= 32'h3ed83553;
    11'b01000100111: data <= 32'h3a193c21;
    11'b01000101000: data <= 32'hbc922856;
    11'b01000101001: data <= 32'hc012bc22;
    11'b01000101010: data <= 32'hbeb3b809;
    11'b01000101011: data <= 32'hbcda39cc;
    11'b01000101100: data <= 32'hbb9438c3;
    11'b01000101101: data <= 32'hb19cba3c;
    11'b01000101110: data <= 32'h3b58bc70;
    11'b01000101111: data <= 32'h3c3738e3;
    11'b01000110000: data <= 32'h1af54100;
    11'b01000110001: data <= 32'hb96040e8;
    11'b01000110010: data <= 32'h2c1c3b77;
    11'b01000110011: data <= 32'h3bd6b162;
    11'b01000110100: data <= 32'h37e9b598;
    11'b01000110101: data <= 32'hb8ebb8aa;
    11'b01000110110: data <= 32'hb340bc6d;
    11'b01000110111: data <= 32'h3ee4bbfa;
    11'b01000111000: data <= 32'h4194ae4d;
    11'b01000111001: data <= 32'h3db8357f;
    11'b01000111010: data <= 32'hba9fb4ec;
    11'b01000111011: data <= 32'hbea5bb13;
    11'b01000111100: data <= 32'hbc2eb569;
    11'b01000111101: data <= 32'hb90a3513;
    11'b01000111110: data <= 32'hbb5bb758;
    11'b01000111111: data <= 32'hbaebbfc7;
    11'b01001000000: data <= 32'had28bf2b;
    11'b01001000001: data <= 32'h35e937c2;
    11'b01001000010: data <= 32'hafbb4105;
    11'b01001000011: data <= 32'hb8c64084;
    11'b01001000100: data <= 32'hb4043999;
    11'b01001000101: data <= 32'h2d3c2a47;
    11'b01001000110: data <= 32'hb86a3856;
    11'b01001000111: data <= 32'hbcb338ff;
    11'b01001001000: data <= 32'hae3db345;
    11'b01001001001: data <= 32'h4053ba2a;
    11'b01001001010: data <= 32'h4222b39f;
    11'b01001001011: data <= 32'h3e2536cd;
    11'b01001001100: data <= 32'hb75a3474;
    11'b01001001101: data <= 32'hb9c3af4f;
    11'b01001001110: data <= 32'h32971b20;
    11'b01001001111: data <= 32'h347cac14;
    11'b01001010000: data <= 32'hba11bd0c;
    11'b01001010001: data <= 32'hbce6c140;
    11'b01001010010: data <= 32'hb59ac053;
    11'b01001010011: data <= 32'h38872e1f;
    11'b01001010100: data <= 32'h351f3ede;
    11'b01001010101: data <= 32'hb7d33cb0;
    11'b01001010110: data <= 32'hba92ad24;
    11'b01001010111: data <= 32'hbb832c16;
    11'b01001011000: data <= 32'hbddd3cd6;
    11'b01001011001: data <= 32'hbeab3d37;
    11'b01001011010: data <= 32'hb602a75f;
    11'b01001011011: data <= 32'h3ebbbb76;
    11'b01001011100: data <= 32'h40aab270;
    11'b01001011101: data <= 32'h3c173c3d;
    11'b01001011110: data <= 32'hb3463d61;
    11'b01001011111: data <= 32'h335d3aab;
    11'b01001100000: data <= 32'h3d043714;
    11'b01001100001: data <= 32'h3a81a444;
    11'b01001100010: data <= 32'hba08bcc1;
    11'b01001100011: data <= 32'hbcd3c0af;
    11'b01001100100: data <= 32'h3171bff2;
    11'b01001100101: data <= 32'h3e08b55c;
    11'b01001100110: data <= 32'h3c8d38cb;
    11'b01001100111: data <= 32'hb3c7ae19;
    11'b01001101000: data <= 32'hbc59ba86;
    11'b01001101001: data <= 32'hbd282620;
    11'b01001101010: data <= 32'hbe763d80;
    11'b01001101011: data <= 32'hbf303c58;
    11'b01001101100: data <= 32'hbb69b985;
    11'b01001101101: data <= 32'h3877be1b;
    11'b01001101110: data <= 32'h3c3bb2b4;
    11'b01001101111: data <= 32'h34583e93;
    11'b01001110000: data <= 32'hb1964023;
    11'b01001110001: data <= 32'h39843d3e;
    11'b01001110010: data <= 32'h3dd939fb;
    11'b01001110011: data <= 32'h384c381f;
    11'b01001110100: data <= 32'hbc63b319;
    11'b01001110101: data <= 32'hbc25bd07;
    11'b01001110110: data <= 32'h3bbebd9d;
    11'b01001110111: data <= 32'h40f8b8b7;
    11'b01001111000: data <= 32'h3f32b1f8;
    11'b01001111001: data <= 32'h2c37b9ea;
    11'b01001111010: data <= 32'hb9fcbb80;
    11'b01001111011: data <= 32'hb91030c5;
    11'b01001111100: data <= 32'hbad73c9a;
    11'b01001111101: data <= 32'hbdfa3433;
    11'b01001111110: data <= 32'hbdbfbef4;
    11'b01001111111: data <= 32'hb829c071;
    11'b01010000000: data <= 32'h2c8fb617;
    11'b01010000001: data <= 32'hb0bf3e90;
    11'b01010000010: data <= 32'hb16e3f5c;
    11'b01010000011: data <= 32'h386a3b77;
    11'b01010000100: data <= 32'h3a8839d2;
    11'b01010000101: data <= 32'hb5f63cf4;
    11'b01010000110: data <= 32'hbebb3c36;
    11'b01010000111: data <= 32'hbbf8ad35;
    11'b01010001000: data <= 32'h3d68bae2;
    11'b01010001001: data <= 32'h4173b904;
    11'b01010001010: data <= 32'h3f31b45a;
    11'b01010001011: data <= 32'h33d2b6d1;
    11'b01010001100: data <= 32'h2a19b544;
    11'b01010001101: data <= 32'h396b3825;
    11'b01010001110: data <= 32'h356e3b26;
    11'b01010001111: data <= 32'hbc06b721;
    11'b01010010000: data <= 32'hbeabc0c0;
    11'b01010010001: data <= 32'hbb8bc10b;
    11'b01010010010: data <= 32'ha5d7b910;
    11'b01010010011: data <= 32'h2e533bb2;
    11'b01010010100: data <= 32'ha9a53997;
    11'b01010010101: data <= 32'h3036af3d;
    11'b01010010110: data <= 32'hacc236ac;
    11'b01010010111: data <= 32'hbcf33f07;
    11'b01010011000: data <= 32'hc0493f7c;
    11'b01010011001: data <= 32'hbcc436c3;
    11'b01010011010: data <= 32'h3ba1ba59;
    11'b01010011011: data <= 32'h3fc3b8b3;
    11'b01010011100: data <= 32'h3c2b3250;
    11'b01010011101: data <= 32'h314737a5;
    11'b01010011110: data <= 32'h3abb3878;
    11'b01010011111: data <= 32'h3f6a3ba9;
    11'b01010100000: data <= 32'h3cc13b4e;
    11'b01010100001: data <= 32'hb9e9b6bb;
    11'b01010100010: data <= 32'hbe78c019;
    11'b01010100011: data <= 32'hb8c0c046;
    11'b01010100100: data <= 32'h39cbba37;
    11'b01010100101: data <= 32'h3ab59459;
    11'b01010100110: data <= 32'h3332b983;
    11'b01010100111: data <= 32'haf2cbcb1;
    11'b01010101000: data <= 32'hb7032d74;
    11'b01010101001: data <= 32'hbd6a3f75;
    11'b01010101010: data <= 32'hc0363f4c;
    11'b01010101011: data <= 32'hbdf8a3c3;
    11'b01010101100: data <= 32'ha68bbd22;
    11'b01010101101: data <= 32'h386bb906;
    11'b01010101110: data <= 32'ha89039bb;
    11'b01010101111: data <= 32'hae303cb8;
    11'b01010110000: data <= 32'h3cde3c0a;
    11'b01010110001: data <= 32'h40763c91;
    11'b01010110010: data <= 32'h3ca93cf7;
    11'b01010110011: data <= 32'hbb9136a7;
    11'b01010110100: data <= 32'hbde9bae6;
    11'b01010110101: data <= 32'h2edebcf0;
    11'b01010110110: data <= 32'h3e96b9a1;
    11'b01010110111: data <= 32'h3de9b977;
    11'b01010111000: data <= 32'h3754be04;
    11'b01010111001: data <= 32'h2cdebe4e;
    11'b01010111010: data <= 32'h2eef28e6;
    11'b01010111011: data <= 32'hb80b3ea2;
    11'b01010111100: data <= 32'hbe023c7c;
    11'b01010111101: data <= 32'hbeb3bbd0;
    11'b01010111110: data <= 32'hbbe4bfd1;
    11'b01010111111: data <= 32'hb8d8ba19;
    11'b01011000000: data <= 32'hba203a81;
    11'b01011000001: data <= 32'hb4d93c25;
    11'b01011000010: data <= 32'h3c543880;
    11'b01011000011: data <= 32'h3ee73ad6;
    11'b01011000100: data <= 32'h35fd3e9b;
    11'b01011000101: data <= 32'hbdfe3e43;
    11'b01011000110: data <= 32'hbdb837b5;
    11'b01011000111: data <= 32'h385bb5b9;
    11'b01011001000: data <= 32'h3fcbb7dd;
    11'b01011001001: data <= 32'h3db2ba03;
    11'b01011001010: data <= 32'h368fbd63;
    11'b01011001011: data <= 32'h38afbc7e;
    11'b01011001100: data <= 32'h3d2c35b5;
    11'b01011001101: data <= 32'h3acd3da9;
    11'b01011001110: data <= 32'hb9543668;
    11'b01011001111: data <= 32'hbe7cbe9d;
    11'b01011010000: data <= 32'hbd7ac070;
    11'b01011010001: data <= 32'hbaf6baa8;
    11'b01011010010: data <= 32'hb9b73627;
    11'b01011010011: data <= 32'hb419235d;
    11'b01011010100: data <= 32'h397eb913;
    11'b01011010101: data <= 32'h3add323c;
    11'b01011010110: data <= 32'hb80f3f74;
    11'b01011010111: data <= 32'hbfc240a6;
    11'b01011011000: data <= 32'hbdf53cad;
    11'b01011011001: data <= 32'h35b7aab3;
    11'b01011011010: data <= 32'h3d18b55d;
    11'b01011011011: data <= 32'h3842b4ea;
    11'b01011011100: data <= 32'h9ff8b801;
    11'b01011011101: data <= 32'h3c42b3d9;
    11'b01011011110: data <= 32'h40cb3a51;
    11'b01011011111: data <= 32'h3f923d5e;
    11'b01011100000: data <= 32'hafb23415;
    11'b01011100001: data <= 32'hbda7bdb6;
    11'b01011100010: data <= 32'hbc26bee0;
    11'b01011100011: data <= 32'hb2c2b947;
    11'b01011100100: data <= 32'ha4deb444;
    11'b01011100101: data <= 32'h2017bd2d;
    11'b01011100110: data <= 32'h3638bf95;
    11'b01011100111: data <= 32'h35d5b734;
    11'b01011101000: data <= 32'hb9be3f16;
    11'b01011101001: data <= 32'hbf404090;
    11'b01011101010: data <= 32'hbe063ac6;
    11'b01011101011: data <= 32'hb52ab754;
    11'b01011101100: data <= 32'ha7e0b5c2;
    11'b01011101101: data <= 32'hba013390;
    11'b01011101110: data <= 32'hb8df34aa;
    11'b01011101111: data <= 32'h3cd334a8;
    11'b01011110000: data <= 32'h41893b50;
    11'b01011110001: data <= 32'h40053db5;
    11'b01011110010: data <= 32'hb25d3a7f;
    11'b01011110011: data <= 32'hbcf0b545;
    11'b01011110100: data <= 32'hb547b8ec;
    11'b01011110101: data <= 32'h3a1cb361;
    11'b01011110110: data <= 32'h3986b981;
    11'b01011110111: data <= 32'h32adc02f;
    11'b01011111000: data <= 32'h3610c0ef;
    11'b01011111001: data <= 32'h3944b962;
    11'b01011111010: data <= 32'h28ce3dfc;
    11'b01011111011: data <= 32'hbc173e53;
    11'b01011111100: data <= 32'hbd4fb03f;
    11'b01011111101: data <= 32'hbc03bcb6;
    11'b01011111110: data <= 32'hbca9b7b0;
    11'b01011111111: data <= 32'hbeb437ca;
    11'b01100000000: data <= 32'hbc2835ef;
    11'b01100000001: data <= 32'h3bbdab93;
    11'b01100000010: data <= 32'h4089376c;
    11'b01100000011: data <= 32'h3cf13df3;
    11'b01100000100: data <= 32'hba313eaf;
    11'b01100000101: data <= 32'hbcbb3be1;
    11'b01100000110: data <= 32'h332037ad;
    11'b01100000111: data <= 32'h3d06340d;
    11'b01100001000: data <= 32'h39e6b8eb;
    11'b01100001001: data <= 32'h270fbfc8;
    11'b01100001010: data <= 32'h3884c022;
    11'b01100001011: data <= 32'h3e37b5d9;
    11'b01100001100: data <= 32'h3d6c3cfe;
    11'b01100001101: data <= 32'h29bc3a35;
    11'b01100001110: data <= 32'hbbb4bbc3;
    11'b01100001111: data <= 32'hbcd6be2f;
    11'b01100010000: data <= 32'hbdc5b732;
    11'b01100010001: data <= 32'hbedf3595;
    11'b01100010010: data <= 32'hbc30b5f0;
    11'b01100010011: data <= 32'h3874bcd7;
    11'b01100010100: data <= 32'h3d5eb6e1;
    11'b01100010101: data <= 32'h33193d72;
    11'b01100010110: data <= 32'hbd444072;
    11'b01100010111: data <= 32'hbcb03ebd;
    11'b01100011000: data <= 32'h34a43b5c;
    11'b01100011001: data <= 32'h3ac9381f;
    11'b01100011010: data <= 32'hae52b059;
    11'b01100011011: data <= 32'hb8eebc3e;
    11'b01100011100: data <= 32'h3989bc5b;
    11'b01100011101: data <= 32'h40da3131;
    11'b01100011110: data <= 32'h40d23c86;
    11'b01100011111: data <= 32'h3a1e3696;
    11'b01100100000: data <= 32'hb8c1bbfd;
    11'b01100100001: data <= 32'hba83bc74;
    11'b01100100010: data <= 32'hba19ac65;
    11'b01100100011: data <= 32'hbbb02a53;
    11'b01100100100: data <= 32'hb9a3bdbc;
    11'b01100100101: data <= 32'h3391c0f7;
    11'b01100100110: data <= 32'h3950bd20;
    11'b01100100111: data <= 32'hb3403c39;
    11'b01100101000: data <= 32'hbd19402b;
    11'b01100101001: data <= 32'hbc053d6c;
    11'b01100101010: data <= 32'haa1f37f0;
    11'b01100101011: data <= 32'hb2823712;
    11'b01100101100: data <= 32'hbd9136b8;
    11'b01100101101: data <= 32'hbdccaf7d;
    11'b01100101110: data <= 32'h389bb54d;
    11'b01100101111: data <= 32'h41573634;
    11'b01100110000: data <= 32'h41113c43;
    11'b01100110001: data <= 32'h39b73928;
    11'b01100110010: data <= 32'hb6c5b102;
    11'b01100110011: data <= 32'hade49d30;
    11'b01100110100: data <= 32'h355c38df;
    11'b01100110101: data <= 32'haab0ad03;
    11'b01100110110: data <= 32'hb642c02a;
    11'b01100110111: data <= 32'h2f1cc225;
    11'b01100111000: data <= 32'h3943be53;
    11'b01100111001: data <= 32'h344a39ed;
    11'b01100111010: data <= 32'hb7e43d6e;
    11'b01100111011: data <= 32'hb8993476;
    11'b01100111100: data <= 32'hb68bb652;
    11'b01100111101: data <= 32'hbcab3294;
    11'b01100111110: data <= 32'hc0b33a09;
    11'b01100111111: data <= 32'hc003337d;
    11'b01101000000: data <= 32'h33dfb6b8;
    11'b01101000001: data <= 32'h4041a83b;
    11'b01101000010: data <= 32'h3ebd3b12;
    11'b01101000011: data <= 32'h169b3cae;
    11'b01101000100: data <= 32'hb7a93bc1;
    11'b01101000101: data <= 32'h382a3c8a;
    11'b01101000110: data <= 32'h3c483d0f;
    11'b01101000111: data <= 32'h34113062;
    11'b01101001000: data <= 32'hb825bf7e;
    11'b01101001001: data <= 32'h2cd5c13f;
    11'b01101001010: data <= 32'h3cddbcb4;
    11'b01101001011: data <= 32'h3d8738a5;
    11'b01101001100: data <= 32'h38ff380c;
    11'b01101001101: data <= 32'h1913ba37;
    11'b01101001110: data <= 32'hb6c5bc12;
    11'b01101001111: data <= 32'hbd75311a;
    11'b01101010000: data <= 32'hc0bd3a79;
    11'b01101010001: data <= 32'hbfdbb1a9;
    11'b01101010010: data <= 32'haec8bd6a;
    11'b01101010011: data <= 32'h3ca6bbc8;
    11'b01101010100: data <= 32'h379f3823;
    11'b01101010101: data <= 32'hba4c3df1;
    11'b01101010110: data <= 32'hb8833e48;
    11'b01101010111: data <= 32'h3a043e53;
    11'b01101011000: data <= 32'h3bdc3e22;
    11'b01101011001: data <= 32'hb5a238c5;
    11'b01101011010: data <= 32'hbcc8bb9a;
    11'b01101011011: data <= 32'haa64bde7;
    11'b01101011100: data <= 32'h3f48b6ac;
    11'b01101011101: data <= 32'h40a43898;
    11'b01101011110: data <= 32'h3d811d62;
    11'b01101011111: data <= 32'h36f9bc72;
    11'b01101100000: data <= 32'h9524ba9d;
    11'b01101100001: data <= 32'hb9233871;
    11'b01101100010: data <= 32'hbde43a1a;
    11'b01101100011: data <= 32'hbda8bb99;
    11'b01101100100: data <= 32'hb4f8c0fd;
    11'b01101100101: data <= 32'h35f4bf83;
    11'b01101100110: data <= 32'hb4402def;
    11'b01101100111: data <= 32'hbbff3d15;
    11'b01101101000: data <= 32'hb6833cc4;
    11'b01101101001: data <= 32'h39433c35;
    11'b01101101010: data <= 32'h337b3d29;
    11'b01101101011: data <= 32'hbdff3c2c;
    11'b01101101100: data <= 32'hc0312d7a;
    11'b01101101101: data <= 32'hb54fb709;
    11'b01101101110: data <= 32'h3fc42cd6;
    11'b01101101111: data <= 32'h40c5385e;
    11'b01101110000: data <= 32'h3d07211b;
    11'b01101110001: data <= 32'h37c5b8a7;
    11'b01101110010: data <= 32'h390f2fae;
    11'b01101110011: data <= 32'h38433d3a;
    11'b01101110100: data <= 32'hb4e13ab2;
    11'b01101110101: data <= 32'hba9fbdbd;
    11'b01101110110: data <= 32'hb5ebc209;
    11'b01101110111: data <= 32'h3112c04a;
    11'b01101111000: data <= 32'hadb7b0fd;
    11'b01101111001: data <= 32'hb66838ce;
    11'b01101111010: data <= 32'h2e0f29d3;
    11'b01101111011: data <= 32'h3832acd3;
    11'b01101111100: data <= 32'hb8423a48;
    11'b01101111101: data <= 32'hc0c63d28;
    11'b01101111110: data <= 32'hc15038f7;
    11'b01101111111: data <= 32'hb938b29e;
    11'b01110000000: data <= 32'h3dadb071;
    11'b01110000001: data <= 32'h3de234ee;
    11'b01110000010: data <= 32'h356334ad;
    11'b01110000011: data <= 32'h31ae3513;
    11'b01110000100: data <= 32'h3c943cba;
    11'b01110000101: data <= 32'h3db94001;
    11'b01110000110: data <= 32'h35293c66;
    11'b01110000111: data <= 32'hb9c8bcd4;
    11'b01110001000: data <= 32'hb6ffc103;
    11'b01110001001: data <= 32'h3785be43;
    11'b01110001010: data <= 32'h3a2eadd9;
    11'b01110001011: data <= 32'h3907b0cb;
    11'b01110001100: data <= 32'h39eabca0;
    11'b01110001101: data <= 32'h38e3bc0f;
    11'b01110001110: data <= 32'hb96337c1;
    11'b01110001111: data <= 32'hc0b33d63;
    11'b01110010000: data <= 32'hc0f63735;
    11'b01110010001: data <= 32'hba8abaef;
    11'b01110010010: data <= 32'h3859bbc6;
    11'b01110010011: data <= 32'h3023b093;
    11'b01110010100: data <= 32'hba1a375f;
    11'b01110010101: data <= 32'hb1b63a9c;
    11'b01110010110: data <= 32'h3d673e52;
    11'b01110010111: data <= 32'h3e4b405e;
    11'b01110011000: data <= 32'h1f4a3dae;
    11'b01110011001: data <= 32'hbd14b5ba;
    11'b01110011010: data <= 32'hb934bcf4;
    11'b01110011011: data <= 32'h3b21b811;
    11'b01110011100: data <= 32'h3e5631d1;
    11'b01110011101: data <= 32'h3d5ab8d2;
    11'b01110011110: data <= 32'h3c89bed7;
    11'b01110011111: data <= 32'h3b98bc86;
    11'b01110100000: data <= 32'h9a0639c8;
    11'b01110100001: data <= 32'hbd633d84;
    11'b01110100010: data <= 32'hbea0af74;
    11'b01110100011: data <= 32'hb9f5bf66;
    11'b01110100100: data <= 32'hb1d6bf57;
    11'b01110100101: data <= 32'hba95b895;
    11'b01110100110: data <= 32'hbd30345b;
    11'b01110100111: data <= 32'hb2b3378b;
    11'b01110101000: data <= 32'h3d473baf;
    11'b01110101001: data <= 32'h3c2d3eca;
    11'b01110101010: data <= 32'hbba43e6a;
    11'b01110101011: data <= 32'hc03f38d5;
    11'b01110101100: data <= 32'hbbc9939b;
    11'b01110101101: data <= 32'h3be03520;
    11'b01110101110: data <= 32'h3e9335f7;
    11'b01110101111: data <= 32'h3c94b921;
    11'b01110110000: data <= 32'h3bdfbda3;
    11'b01110110001: data <= 32'h3d65b654;
    11'b01110110010: data <= 32'h3c633dab;
    11'b01110110011: data <= 32'h21b43e15;
    11'b01110110100: data <= 32'hb9cdb835;
    11'b01110110101: data <= 32'hb871c0ae;
    11'b01110110110: data <= 32'hb6a7c017;
    11'b01110110111: data <= 32'hbb0fb95e;
    11'b01110111000: data <= 32'hbb81b291;
    11'b01110111001: data <= 32'h32edb8db;
    11'b01110111010: data <= 32'h3d13b578;
    11'b01110111011: data <= 32'h36453acf;
    11'b01110111100: data <= 32'hbf223e52;
    11'b01110111101: data <= 32'hc14a3c8b;
    11'b01110111110: data <= 32'hbcc6378c;
    11'b01110111111: data <= 32'h38dc360a;
    11'b01111000000: data <= 32'h3a4533a0;
    11'b01111000001: data <= 32'h2c3bb723;
    11'b01111000010: data <= 32'h3599b940;
    11'b01111000011: data <= 32'h3e5638aa;
    11'b01111000100: data <= 32'h3fe4402c;
    11'b01111000101: data <= 32'h3b093eec;
    11'b01111000110: data <= 32'hb515b655;
    11'b01111000111: data <= 32'hb7bfbf78;
    11'b01111001000: data <= 32'hb1f5bd4f;
    11'b01111001001: data <= 32'hb236b4e6;
    11'b01111001010: data <= 32'ha515b979;
    11'b01111001011: data <= 32'h3abfbf19;
    11'b01111001100: data <= 32'h3d64be15;
    11'b01111001101: data <= 32'h326e3318;
    11'b01111001110: data <= 32'hbf183dd9;
    11'b01111001111: data <= 32'hc0b53c22;
    11'b01111010000: data <= 32'hbc602043;
    11'b01111010001: data <= 32'ha2efb4ff;
    11'b01111010010: data <= 32'hb829b228;
    11'b01111010011: data <= 32'hbd14b4ec;
    11'b01111010100: data <= 32'hb5aab092;
    11'b01111010101: data <= 32'h3e523bf5;
    11'b01111010110: data <= 32'h4055405d;
    11'b01111010111: data <= 32'h3a3c3f53;
    11'b01111011000: data <= 32'hb97b3333;
    11'b01111011001: data <= 32'hb94cb91a;
    11'b01111011010: data <= 32'h31bfa91c;
    11'b01111011011: data <= 32'h38a43533;
    11'b01111011100: data <= 32'h397fbb39;
    11'b01111011101: data <= 32'h3cbac0bb;
    11'b01111011110: data <= 32'h3e12bf79;
    11'b01111011111: data <= 32'h396933bc;
    11'b01111100000: data <= 32'hba743dbd;
    11'b01111100001: data <= 32'hbd3f3849;
    11'b01111100010: data <= 32'hb94ebb32;
    11'b01111100011: data <= 32'hb7d2bc9d;
    11'b01111100100: data <= 32'hbdfeb8bc;
    11'b01111100101: data <= 32'hc01ab614;
    11'b01111100110: data <= 32'hb922b573;
    11'b01111100111: data <= 32'h3dd63697;
    11'b01111101000: data <= 32'h3ed83e02;
    11'b01111101001: data <= 32'hacda3eaf;
    11'b01111101010: data <= 32'hbdf93b6f;
    11'b01111101011: data <= 32'hbbc338ee;
    11'b01111101100: data <= 32'h35723c35;
    11'b01111101101: data <= 32'h3a0b3a7d;
    11'b01111101110: data <= 32'h383fba8a;
    11'b01111101111: data <= 32'h3af4c046;
    11'b01111110000: data <= 32'h3e67bd15;
    11'b01111110001: data <= 32'h3e163ae5;
    11'b01111110010: data <= 32'h387b3e44;
    11'b01111110011: data <= 32'haee42e4b;
    11'b01111110100: data <= 32'hb0a5bdde;
    11'b01111110101: data <= 32'hb884bd97;
    11'b01111110110: data <= 32'hbe83b87e;
    11'b01111110111: data <= 32'hbf73b8a6;
    11'b01111111000: data <= 32'hb532bcb7;
    11'b01111111001: data <= 32'h3d94bb24;
    11'b01111111010: data <= 32'h3c3e361b;
    11'b01111111011: data <= 32'hbb903d2c;
    11'b01111111100: data <= 32'hc0163d17;
    11'b01111111101: data <= 32'hbc633ca0;
    11'b01111111110: data <= 32'h32363d3f;
    11'b01111111111: data <= 32'h2f413a9e;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    