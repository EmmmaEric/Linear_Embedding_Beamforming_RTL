
module memory_rom_63(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbdb4b95b;
    11'b00000000001: data <= 32'hbb32b55a;
    11'b00000000010: data <= 32'h3a3135f5;
    11'b00000000011: data <= 32'h3cd33db4;
    11'b00000000100: data <= 32'hb79e3e9a;
    11'b00000000101: data <= 32'hc06e39e5;
    11'b00000000110: data <= 32'hbf9d2a6e;
    11'b00000000111: data <= 32'hb194380d;
    11'b00000001000: data <= 32'h3b703bca;
    11'b00000001001: data <= 32'h3b8f2fc5;
    11'b00000001010: data <= 32'h3c11bc79;
    11'b00000001011: data <= 32'h3e06b9a4;
    11'b00000001100: data <= 32'h3dbd3ce1;
    11'b00000001101: data <= 32'h37934046;
    11'b00000001110: data <= 32'hb4023923;
    11'b00000001111: data <= 32'ha78ebe39;
    11'b00000010000: data <= 32'h3210c043;
    11'b00000010001: data <= 32'hb775bcf3;
    11'b00000010010: data <= 32'hbc0fb98b;
    11'b00000010011: data <= 32'haf42bbd2;
    11'b00000010100: data <= 32'h3d82baed;
    11'b00000010101: data <= 32'h3cb93106;
    11'b00000010110: data <= 32'hbbfe3bc6;
    11'b00000010111: data <= 32'hc1733a26;
    11'b00000011000: data <= 32'hc040354c;
    11'b00000011001: data <= 32'hb60337a5;
    11'b00000011010: data <= 32'h3468386b;
    11'b00000011011: data <= 32'hb379b362;
    11'b00000011100: data <= 32'hb1a9bb37;
    11'b00000011101: data <= 32'h3b8b2c89;
    11'b00000011110: data <= 32'h3ebb401e;
    11'b00000011111: data <= 32'h3c64413e;
    11'b00000100000: data <= 32'h30823b1b;
    11'b00000100001: data <= 32'hac6cbc4e;
    11'b00000100010: data <= 32'h2d4bbcd8;
    11'b00000100011: data <= 32'hb042b46e;
    11'b00000100100: data <= 32'hb0bcb596;
    11'b00000100101: data <= 32'h3ae1be06;
    11'b00000100110: data <= 32'h3fd9bf6d;
    11'b00000100111: data <= 32'h3d61b8f7;
    11'b00000101000: data <= 32'hbaa939b4;
    11'b00000101001: data <= 32'hc07239e7;
    11'b00000101010: data <= 32'hbe122193;
    11'b00000101011: data <= 32'hb47eb4eb;
    11'b00000101100: data <= 32'hb7cab590;
    11'b00000101101: data <= 32'hbe0db9e4;
    11'b00000101110: data <= 32'hbcf8bb01;
    11'b00000101111: data <= 32'h382b3469;
    11'b00000110000: data <= 32'h3eba4010;
    11'b00000110001: data <= 32'h3bb240d2;
    11'b00000110010: data <= 32'hb6713c0c;
    11'b00000110011: data <= 32'hb9f3b2b0;
    11'b00000110100: data <= 32'hb2e431c0;
    11'b00000110101: data <= 32'h30a83b51;
    11'b00000110110: data <= 32'h368c2de7;
    11'b00000110111: data <= 32'h3cfbbec2;
    11'b00000111000: data <= 32'h402cc022;
    11'b00000111001: data <= 32'h3e66b72c;
    11'b00000111010: data <= 32'ha4df3c5b;
    11'b00000111011: data <= 32'hbb813a6c;
    11'b00000111100: data <= 32'hb66bb7fd;
    11'b00000111101: data <= 32'h2a13bc8a;
    11'b00000111110: data <= 32'hbb8abc08;
    11'b00000111111: data <= 32'hc04ebc2a;
    11'b00001000000: data <= 32'hbe0abc7a;
    11'b00001000001: data <= 32'h38c0b556;
    11'b00001000010: data <= 32'h3e5c3c24;
    11'b00001000011: data <= 32'h357d3e32;
    11'b00001000100: data <= 32'hbd6e3b34;
    11'b00001000101: data <= 32'hbe113838;
    11'b00001000110: data <= 32'hb82e3cdd;
    11'b00001000111: data <= 32'h2cd13e5b;
    11'b00001001000: data <= 32'h30393440;
    11'b00001001001: data <= 32'h3924be47;
    11'b00001001010: data <= 32'h3e47be20;
    11'b00001001011: data <= 32'h3efb370c;
    11'b00001001100: data <= 32'h3b8d3f42;
    11'b00001001101: data <= 32'h35d63bd4;
    11'b00001001110: data <= 32'h3854b9c4;
    11'b00001001111: data <= 32'h3593bd16;
    11'b00001010000: data <= 32'hbb6fba9c;
    11'b00001010001: data <= 32'hbf8cbaca;
    11'b00001010010: data <= 32'hbb18bdda;
    11'b00001010011: data <= 32'h3c88bda5;
    11'b00001010100: data <= 32'h3e4cb5c0;
    11'b00001010101: data <= 32'hb1f7384c;
    11'b00001010110: data <= 32'hbfa03916;
    11'b00001010111: data <= 32'hbeda39f1;
    11'b00001011000: data <= 32'hb8683d5e;
    11'b00001011001: data <= 32'hb5163d77;
    11'b00001011010: data <= 32'hbb281c6d;
    11'b00001011011: data <= 32'hb955bd7d;
    11'b00001011100: data <= 32'h395fba49;
    11'b00001011101: data <= 32'h3eaf3d29;
    11'b00001011110: data <= 32'h3dea4091;
    11'b00001011111: data <= 32'h3b563c62;
    11'b00001100000: data <= 32'h39e7b752;
    11'b00001100001: data <= 32'h35e4b7d7;
    11'b00001100010: data <= 32'hb8ea339a;
    11'b00001100011: data <= 32'hbc53b1bd;
    11'b00001100100: data <= 32'h2c56bea2;
    11'b00001100101: data <= 32'h3ed7c096;
    11'b00001100110: data <= 32'h3e9abd35;
    11'b00001100111: data <= 32'hb2201d0f;
    11'b00001101000: data <= 32'hbe1a36f8;
    11'b00001101001: data <= 32'hbc1236e2;
    11'b00001101010: data <= 32'hb0d93929;
    11'b00001101011: data <= 32'hb9ff3824;
    11'b00001101100: data <= 32'hc01bb7e6;
    11'b00001101101: data <= 32'hbf99bd2f;
    11'b00001101110: data <= 32'hab38b741;
    11'b00001101111: data <= 32'h3dd43d78;
    11'b00001110000: data <= 32'h3d544003;
    11'b00001110001: data <= 32'h37c73b90;
    11'b00001110010: data <= 32'h30e92df6;
    11'b00001110011: data <= 32'h2db33a38;
    11'b00001110100: data <= 32'hb50c3e64;
    11'b00001110101: data <= 32'hb70638be;
    11'b00001110110: data <= 32'h3857be5c;
    11'b00001110111: data <= 32'h3f28c0f2;
    11'b00001111000: data <= 32'h3eaebd0d;
    11'b00001111001: data <= 32'h354233ee;
    11'b00001111010: data <= 32'hb5d13756;
    11'b00001111011: data <= 32'h343bad35;
    11'b00001111100: data <= 32'h382fb348;
    11'b00001111101: data <= 32'hbb63b2dd;
    11'b00001111110: data <= 32'hc14bba36;
    11'b00001111111: data <= 32'hc0a3bd65;
    11'b00010000000: data <= 32'hb129ba64;
    11'b00010000001: data <= 32'h3d2837e4;
    11'b00010000010: data <= 32'h39c13be6;
    11'b00010000011: data <= 32'hb7a737b9;
    11'b00010000100: data <= 32'hb9563838;
    11'b00010000101: data <= 32'hb2d73f05;
    11'b00010000110: data <= 32'hb3b740e3;
    11'b00010000111: data <= 32'hb7cb3bea;
    11'b00010001000: data <= 32'h2bf9bd6c;
    11'b00010001001: data <= 32'h3c8bbfc5;
    11'b00010001010: data <= 32'h3de4b65b;
    11'b00010001011: data <= 32'h3bd43bf0;
    11'b00010001100: data <= 32'h3af8391a;
    11'b00010001101: data <= 32'h3d95b681;
    11'b00010001110: data <= 32'h3c5db873;
    11'b00010001111: data <= 32'hba0db0dd;
    11'b00010010000: data <= 32'hc0c3b794;
    11'b00010010001: data <= 32'hbf00bd7e;
    11'b00010010010: data <= 32'h35ccbe41;
    11'b00010010011: data <= 32'h3d1aba99;
    11'b00010010100: data <= 32'h2f97b33a;
    11'b00010010101: data <= 32'hbcbbadab;
    11'b00010010110: data <= 32'hbbd53866;
    11'b00010010111: data <= 32'hb12e3f80;
    11'b00010011000: data <= 32'hb596409d;
    11'b00010011001: data <= 32'hbcd83a46;
    11'b00010011010: data <= 32'hbca6bc95;
    11'b00010011011: data <= 32'h2823bc98;
    11'b00010011100: data <= 32'h3c40389a;
    11'b00010011101: data <= 32'h3d233e48;
    11'b00010011110: data <= 32'h3da6399f;
    11'b00010011111: data <= 32'h3edcb63a;
    11'b00010100000: data <= 32'h3cddab75;
    11'b00010100001: data <= 32'hb6833a90;
    11'b00010100010: data <= 32'hbe2e364c;
    11'b00010100011: data <= 32'hb9a3bcdd;
    11'b00010100100: data <= 32'h3c26c060;
    11'b00010100101: data <= 32'h3d4cbf00;
    11'b00010100110: data <= 32'hadf6bb52;
    11'b00010100111: data <= 32'hbc42b72a;
    11'b00010101000: data <= 32'hb6203182;
    11'b00010101001: data <= 32'h36b43ca4;
    11'b00010101010: data <= 32'hb6da3d9c;
    11'b00010101011: data <= 32'hc0313298;
    11'b00010101100: data <= 32'hc0bebc3f;
    11'b00010101101: data <= 32'hbb0fb92d;
    11'b00010101110: data <= 32'h39173b25;
    11'b00010101111: data <= 32'h3c253d99;
    11'b00010110000: data <= 32'h3bc6364f;
    11'b00010110001: data <= 32'h3c74b1bc;
    11'b00010110010: data <= 32'h3b133b6c;
    11'b00010110011: data <= 32'haf03404d;
    11'b00010110100: data <= 32'hba213d80;
    11'b00010110101: data <= 32'ha16abb1c;
    11'b00010110110: data <= 32'h3cefc075;
    11'b00010110111: data <= 32'h3cdcbed4;
    11'b00010111000: data <= 32'h2ed0b997;
    11'b00010111001: data <= 32'hb1e9b699;
    11'b00010111010: data <= 32'h3aecb572;
    11'b00010111011: data <= 32'h3d4431cd;
    11'b00010111100: data <= 32'hb4e1379c;
    11'b00010111101: data <= 32'hc109b280;
    11'b00010111110: data <= 32'hc195bc13;
    11'b00010111111: data <= 32'hbc3bb996;
    11'b00011000000: data <= 32'h36e934cb;
    11'b00011000001: data <= 32'h368936cc;
    11'b00011000010: data <= 32'hacbfb4bd;
    11'b00011000011: data <= 32'h3013ac60;
    11'b00011000100: data <= 32'h37413ed4;
    11'b00011000101: data <= 32'h27294201;
    11'b00011000110: data <= 32'hb8693f8b;
    11'b00011000111: data <= 32'hb2deb883;
    11'b00011001000: data <= 32'h391ebea4;
    11'b00011001001: data <= 32'h3a60ba3b;
    11'b00011001010: data <= 32'h36af31ae;
    11'b00011001011: data <= 32'h3aa9af51;
    11'b00011001100: data <= 32'h4004b99f;
    11'b00011001101: data <= 32'h4015b60a;
    11'b00011001110: data <= 32'h1d52344b;
    11'b00011001111: data <= 32'hc05f2508;
    11'b00011010000: data <= 32'hc05bbabc;
    11'b00011010001: data <= 32'hb70ebc7b;
    11'b00011010010: data <= 32'h3820ba48;
    11'b00011010011: data <= 32'hb2dfba70;
    11'b00011010100: data <= 32'hbbd4bc3f;
    11'b00011010101: data <= 32'hb71ab3b0;
    11'b00011010110: data <= 32'h36783ef2;
    11'b00011010111: data <= 32'h2dec41ae;
    11'b00011011000: data <= 32'hbb863e86;
    11'b00011011001: data <= 32'hbcc6b6c0;
    11'b00011011010: data <= 32'hb79fbacb;
    11'b00011011011: data <= 32'h313d35df;
    11'b00011011100: data <= 32'h37bc3c01;
    11'b00011011101: data <= 32'h3d082c6f;
    11'b00011011110: data <= 32'h40a5ba9b;
    11'b00011011111: data <= 32'h4055b25a;
    11'b00011100000: data <= 32'h353b3be1;
    11'b00011100001: data <= 32'hbd513b1b;
    11'b00011100010: data <= 32'hbbdcb728;
    11'b00011100011: data <= 32'h3765bddf;
    11'b00011100100: data <= 32'h398ebe4a;
    11'b00011100101: data <= 32'hb84bbe08;
    11'b00011100110: data <= 32'hbca3bde8;
    11'b00011100111: data <= 32'haf09b91b;
    11'b00011101000: data <= 32'h3bc03bf2;
    11'b00011101001: data <= 32'h34053f3e;
    11'b00011101010: data <= 32'hbe183aca;
    11'b00011101011: data <= 32'hc07db786;
    11'b00011101100: data <= 32'hbdb0b430;
    11'b00011101101: data <= 32'hb5f63bb9;
    11'b00011101110: data <= 32'h31313c65;
    11'b00011101111: data <= 32'h3a35b26b;
    11'b00011110000: data <= 32'h3e7fbabe;
    11'b00011110001: data <= 32'h3ea93790;
    11'b00011110010: data <= 32'h37f94047;
    11'b00011110011: data <= 32'hb7c63fa4;
    11'b00011110100: data <= 32'ha6c228c4;
    11'b00011110101: data <= 32'h3b78bd89;
    11'b00011110110: data <= 32'h3930bde1;
    11'b00011110111: data <= 32'hb85dbce6;
    11'b00011111000: data <= 32'hb8cbbd44;
    11'b00011111001: data <= 32'h3b92bc2d;
    11'b00011111010: data <= 32'h3fa6a8c7;
    11'b00011111011: data <= 32'h388b3922;
    11'b00011111100: data <= 32'hbf16312a;
    11'b00011111101: data <= 32'hc12db825;
    11'b00011111110: data <= 32'hbe3fb013;
    11'b00011111111: data <= 32'hb80b3989;
    11'b00100000000: data <= 32'hb6463550;
    11'b00100000001: data <= 32'hb508bb76;
    11'b00100000010: data <= 32'h36b5bb9a;
    11'b00100000011: data <= 32'h3bb03c2b;
    11'b00100000100: data <= 32'h382f41cd;
    11'b00100000101: data <= 32'haf1a40d5;
    11'b00100000110: data <= 32'h2da3358f;
    11'b00100000111: data <= 32'h3888bac5;
    11'b00100001000: data <= 32'h3274b7f7;
    11'b00100001001: data <= 32'hb77ab10a;
    11'b00100001010: data <= 32'h31abba15;
    11'b00100001011: data <= 32'h3ff4bd1e;
    11'b00100001100: data <= 32'h4151b9d9;
    11'b00100001101: data <= 32'h3b5c2fbb;
    11'b00100001110: data <= 32'hbdb73052;
    11'b00100001111: data <= 32'hbfb3b559;
    11'b00100010000: data <= 32'hba44b505;
    11'b00100010001: data <= 32'hb224b018;
    11'b00100010010: data <= 32'hbb19ba43;
    11'b00100010011: data <= 32'hbd55befc;
    11'b00100010100: data <= 32'hb751bcde;
    11'b00100010101: data <= 32'h39233c0e;
    11'b00100010110: data <= 32'h3884415f;
    11'b00100010111: data <= 32'hb4584011;
    11'b00100011000: data <= 32'hb8d934c3;
    11'b00100011001: data <= 32'hb6adb0da;
    11'b00100011010: data <= 32'hb7ee39fb;
    11'b00100011011: data <= 32'hb85a3bae;
    11'b00100011100: data <= 32'h3809b4b1;
    11'b00100011101: data <= 32'h407fbd66;
    11'b00100011110: data <= 32'h4165ba20;
    11'b00100011111: data <= 32'h3c63384e;
    11'b00100100000: data <= 32'hb9563aca;
    11'b00100100001: data <= 32'hb91f301c;
    11'b00100100010: data <= 32'h3664b7b4;
    11'b00100100011: data <= 32'h346dba39;
    11'b00100100100: data <= 32'hbc86bdbb;
    11'b00100100101: data <= 32'hbed7c03b;
    11'b00100100110: data <= 32'hb6eebe19;
    11'b00100100111: data <= 32'h3c1a356e;
    11'b00100101000: data <= 32'h3a433e4c;
    11'b00100101001: data <= 32'hb9323bef;
    11'b00100101010: data <= 32'hbdf0a8de;
    11'b00100101011: data <= 32'hbd38356f;
    11'b00100101100: data <= 32'hbc1d3e1b;
    11'b00100101101: data <= 32'hbaaa3d81;
    11'b00100101110: data <= 32'h2b7eb5ab;
    11'b00100101111: data <= 32'h3de9bda1;
    11'b00100110000: data <= 32'h3fdbb4fd;
    11'b00100110001: data <= 32'h3bf53df7;
    11'b00100110010: data <= 32'h2c863f39;
    11'b00100110011: data <= 32'h37be3928;
    11'b00100110100: data <= 32'h3ccab5f0;
    11'b00100110101: data <= 32'h377db969;
    11'b00100110110: data <= 32'hbca1bc5a;
    11'b00100110111: data <= 32'hbd7cbf0d;
    11'b00100111000: data <= 32'h3657bebc;
    11'b00100111001: data <= 32'h3f8fb8ac;
    11'b00100111010: data <= 32'h3c9f33ff;
    11'b00100111011: data <= 32'hba92a6f8;
    11'b00100111100: data <= 32'hbf2cb597;
    11'b00100111101: data <= 32'hbd933776;
    11'b00100111110: data <= 32'hbc0e3de6;
    11'b00100111111: data <= 32'hbcba3ae1;
    11'b00101000000: data <= 32'hbb77bbe8;
    11'b00101000001: data <= 32'h3026be56;
    11'b00101000010: data <= 32'h3b70307b;
    11'b00101000011: data <= 32'h39df405e;
    11'b00101000100: data <= 32'h36994089;
    11'b00101000101: data <= 32'h3a8c3ad7;
    11'b00101000110: data <= 32'h3c6d2154;
    11'b00101000111: data <= 32'h30a132d9;
    11'b00101001000: data <= 32'hbc9b2ef6;
    11'b00101001001: data <= 32'hb9f3bb20;
    11'b00101001010: data <= 32'h3d5dbe7f;
    11'b00101001011: data <= 32'h4134bce3;
    11'b00101001100: data <= 32'h3dd1b7cd;
    11'b00101001101: data <= 32'hb8a5b5b2;
    11'b00101001110: data <= 32'hbcc3b528;
    11'b00101001111: data <= 32'hb8033588;
    11'b00101010000: data <= 32'hb68c3aa3;
    11'b00101010001: data <= 32'hbd8ab021;
    11'b00101010010: data <= 32'hbf86bf15;
    11'b00101010011: data <= 32'hbba9bf5d;
    11'b00101010100: data <= 32'h3490313b;
    11'b00101010101: data <= 32'h38a84003;
    11'b00101010110: data <= 32'h34d53f29;
    11'b00101010111: data <= 32'h35183863;
    11'b00101011000: data <= 32'h347436e7;
    11'b00101011001: data <= 32'hb8243d88;
    11'b00101011010: data <= 32'hbd033db8;
    11'b00101011011: data <= 32'hb69ead25;
    11'b00101011100: data <= 32'h3e76bddc;
    11'b00101011101: data <= 32'h4120bd24;
    11'b00101011110: data <= 32'h3daab475;
    11'b00101011111: data <= 32'hac1b315e;
    11'b00101100000: data <= 32'h252d2ddd;
    11'b00101100001: data <= 32'h3b043354;
    11'b00101100010: data <= 32'h36943316;
    11'b00101100011: data <= 32'hbd7cba2f;
    11'b00101100100: data <= 32'hc087c02c;
    11'b00101100101: data <= 32'hbc9cbfec;
    11'b00101100110: data <= 32'h3715b4d9;
    11'b00101100111: data <= 32'h39cf3bb5;
    11'b00101101000: data <= 32'ha1c4387e;
    11'b00101101001: data <= 32'hb7a9b068;
    11'b00101101010: data <= 32'hb8a5392e;
    11'b00101101011: data <= 32'hbc14404d;
    11'b00101101100: data <= 32'hbdb54026;
    11'b00101101101: data <= 32'hb98b2fb4;
    11'b00101101110: data <= 32'h3b41bdaa;
    11'b00101101111: data <= 32'h3ea5bb2f;
    11'b00101110000: data <= 32'h3bcc387b;
    11'b00101110001: data <= 32'h36443c46;
    11'b00101110010: data <= 32'h3c7d38ba;
    11'b00101110011: data <= 32'h3fa53460;
    11'b00101110100: data <= 32'h3b303270;
    11'b00101110101: data <= 32'hbd06b7ba;
    11'b00101110110: data <= 32'hbff1be5c;
    11'b00101110111: data <= 32'hb770bf4e;
    11'b00101111000: data <= 32'h3ce2bb95;
    11'b00101111001: data <= 32'h3c57b54d;
    11'b00101111010: data <= 32'hb2a0b99a;
    11'b00101111011: data <= 32'hbae9ba36;
    11'b00101111100: data <= 32'hb9b738c5;
    11'b00101111101: data <= 32'hbb22404d;
    11'b00101111110: data <= 32'hbdff3ee6;
    11'b00101111111: data <= 32'hbdafb64d;
    11'b00110000000: data <= 32'hb679be4a;
    11'b00110000001: data <= 32'h3621b741;
    11'b00110000010: data <= 32'h35ca3d27;
    11'b00110000011: data <= 32'h382e3e43;
    11'b00110000100: data <= 32'h3dfd39c2;
    11'b00110000101: data <= 32'h400636d0;
    11'b00110000110: data <= 32'h39de3ad1;
    11'b00110000111: data <= 32'hbcdb3962;
    11'b00110001000: data <= 32'hbd8cb7b6;
    11'b00110001001: data <= 32'h37a6bd9a;
    11'b00110001010: data <= 32'h3fd0bd65;
    11'b00110001011: data <= 32'h3d53bc67;
    11'b00110001100: data <= 32'hb0b1bcfe;
    11'b00110001101: data <= 32'hb77fbb9e;
    11'b00110001110: data <= 32'h304a36a6;
    11'b00110001111: data <= 32'hac573e30;
    11'b00110010000: data <= 32'hbd5b3a2b;
    11'b00110010001: data <= 32'hc03abcb9;
    11'b00110010010: data <= 32'hbe0fbf32;
    11'b00110010011: data <= 32'hb809b4be;
    11'b00110010100: data <= 32'ha9063d23;
    11'b00110010101: data <= 32'h35203c88;
    11'b00110010110: data <= 32'h3c323300;
    11'b00110010111: data <= 32'h3d053800;
    11'b00110011000: data <= 32'h2dac3f0b;
    11'b00110011001: data <= 32'hbd344005;
    11'b00110011010: data <= 32'hbbb938b7;
    11'b00110011011: data <= 32'h3b2abb98;
    11'b00110011100: data <= 32'h3fdbbd23;
    11'b00110011101: data <= 32'h3c84bb94;
    11'b00110011110: data <= 32'h2a80baa9;
    11'b00110011111: data <= 32'h37cdb8b3;
    11'b00110100000: data <= 32'h3e1734a6;
    11'b00110100001: data <= 32'h3c183b14;
    11'b00110100010: data <= 32'hbbfe240b;
    11'b00110100011: data <= 32'hc0acbe34;
    11'b00110100100: data <= 32'hbf10bf3d;
    11'b00110100101: data <= 32'hb7e7b7a9;
    11'b00110100110: data <= 32'h230937bd;
    11'b00110100111: data <= 32'h9fdaae66;
    11'b00110101000: data <= 32'h3352b9ec;
    11'b00110101001: data <= 32'h351535df;
    11'b00110101010: data <= 32'hb77c40af;
    11'b00110101011: data <= 32'hbd87416b;
    11'b00110101100: data <= 32'hbc003bcc;
    11'b00110101101: data <= 32'h36a0ba16;
    11'b00110101110: data <= 32'h3c43bae8;
    11'b00110101111: data <= 32'h36c3aefe;
    11'b00110110000: data <= 32'h30b12f29;
    11'b00110110001: data <= 32'h3d88a90b;
    11'b00110110010: data <= 32'h413b3469;
    11'b00110110011: data <= 32'h3eec394d;
    11'b00110110100: data <= 32'hb98e2e1a;
    11'b00110110101: data <= 32'hbfffbc49;
    11'b00110110110: data <= 32'hbc62bda3;
    11'b00110110111: data <= 32'h34a1ba1e;
    11'b00110111000: data <= 32'h367cb8bf;
    11'b00110111001: data <= 32'hb3a2bdb0;
    11'b00110111010: data <= 32'hb50fbe86;
    11'b00110111011: data <= 32'h9f6f2d21;
    11'b00110111100: data <= 32'hb5ff4082;
    11'b00110111101: data <= 32'hbcf440c9;
    11'b00110111110: data <= 32'hbd8737ed;
    11'b00110111111: data <= 32'hb963bb63;
    11'b00111000000: data <= 32'hb45ab658;
    11'b00111000001: data <= 32'hb77e39ef;
    11'b00111000010: data <= 32'h000f3a38;
    11'b00111000011: data <= 32'h3e98307b;
    11'b00111000100: data <= 32'h418733fa;
    11'b00111000101: data <= 32'h3e943bf0;
    11'b00111000110: data <= 32'hb8fb3c19;
    11'b00111000111: data <= 32'hbd842dc0;
    11'b00111001000: data <= 32'habd8b986;
    11'b00111001001: data <= 32'h3cabbad3;
    11'b00111001010: data <= 32'h39b3bceb;
    11'b00111001011: data <= 32'hb51ac011;
    11'b00111001100: data <= 32'hb2c6bfbc;
    11'b00111001101: data <= 32'h38f0b189;
    11'b00111001110: data <= 32'h37cf3e81;
    11'b00111001111: data <= 32'hba473d7f;
    11'b00111010000: data <= 32'hbef5b68d;
    11'b00111010001: data <= 32'hbe86bcdc;
    11'b00111010010: data <= 32'hbcf4b03f;
    11'b00111010011: data <= 32'hbc2f3bf6;
    11'b00111010100: data <= 32'hb52b3882;
    11'b00111010101: data <= 32'h3ca5b61a;
    11'b00111010110: data <= 32'h3fe02988;
    11'b00111010111: data <= 32'h3b503e39;
    11'b00111011000: data <= 32'hba2d4063;
    11'b00111011001: data <= 32'hbb063d01;
    11'b00111011010: data <= 32'h38a8a417;
    11'b00111011011: data <= 32'h3d90b8ef;
    11'b00111011100: data <= 32'h3816bc17;
    11'b00111011101: data <= 32'hb60dbe70;
    11'b00111011110: data <= 32'h366fbe19;
    11'b00111011111: data <= 32'h3f4fb403;
    11'b00111100000: data <= 32'h3eb23b3c;
    11'b00111100001: data <= 32'hb1ec36c1;
    11'b00111100010: data <= 32'hbef8bbe4;
    11'b00111100011: data <= 32'hbf3ebcff;
    11'b00111100100: data <= 32'hbcfead90;
    11'b00111100101: data <= 32'hbbfc3836;
    11'b00111100110: data <= 32'hb90cb7b8;
    11'b00111100111: data <= 32'h34bbbdbc;
    11'b00111101000: data <= 32'h3ae8b5fa;
    11'b00111101001: data <= 32'h311e3f83;
    11'b00111101010: data <= 32'hbb2f419c;
    11'b00111101011: data <= 32'hb9bd3ebc;
    11'b00111101100: data <= 32'h36b1336f;
    11'b00111101101: data <= 32'h397fb1b4;
    11'b00111101110: data <= 32'hb47cb09c;
    11'b00111101111: data <= 32'hb8a0b83a;
    11'b00111110000: data <= 32'h3c0cba5d;
    11'b00111110001: data <= 32'h41a2b27b;
    11'b00111110010: data <= 32'h40e83829;
    11'b00111110011: data <= 32'h33853271;
    11'b00111110100: data <= 32'hbd5eb9b0;
    11'b00111110101: data <= 32'hbc64ba3f;
    11'b00111110110: data <= 32'hb5c7ace1;
    11'b00111110111: data <= 32'hb742b3e1;
    11'b00111111000: data <= 32'hba56bec5;
    11'b00111111001: data <= 32'hb617c0d8;
    11'b00111111010: data <= 32'h3420ba9f;
    11'b00111111011: data <= 32'h28cc3ebc;
    11'b00111111100: data <= 32'hb9b340e1;
    11'b00111111101: data <= 32'hba813c8a;
    11'b00111111110: data <= 32'hb5a7a9c7;
    11'b00111111111: data <= 32'hb83b3337;
    11'b01000000000: data <= 32'hbd253a83;
    11'b01000000001: data <= 32'hbb833653;
    11'b01000000010: data <= 32'h3c81b649;
    11'b01000000011: data <= 32'h41d3b3ba;
    11'b01000000100: data <= 32'h40ab38ab;
    11'b01000000101: data <= 32'h339b3a7a;
    11'b01000000110: data <= 32'hba233505;
    11'b01000000111: data <= 32'h27162bf5;
    11'b01000001000: data <= 32'h3a032d97;
    11'b01000001001: data <= 32'h2cf9b98c;
    11'b01000001010: data <= 32'hbad9c07f;
    11'b01000001011: data <= 32'hb81ec176;
    11'b01000001100: data <= 32'h387dbc42;
    11'b01000001101: data <= 32'h39fa3c49;
    11'b01000001110: data <= 32'hb0693d5d;
    11'b01000001111: data <= 32'hbb23254a;
    11'b01000010000: data <= 32'hbc5bb86f;
    11'b01000010001: data <= 32'hbdbf373a;
    11'b01000010010: data <= 32'hbfa53d1d;
    11'b01000010011: data <= 32'hbd3637f9;
    11'b01000010100: data <= 32'h38ffb9ef;
    11'b01000010101: data <= 32'h4018b86d;
    11'b01000010110: data <= 32'h3db33add;
    11'b01000010111: data <= 32'haf453eea;
    11'b01000011000: data <= 32'hb5103da5;
    11'b01000011001: data <= 32'h3adf3a92;
    11'b01000011010: data <= 32'h3d2436c5;
    11'b01000011011: data <= 32'h2c5cb6f7;
    11'b01000011100: data <= 32'hbbfcbf0c;
    11'b01000011101: data <= 32'hb214c05b;
    11'b01000011110: data <= 32'h3e02bbbb;
    11'b01000011111: data <= 32'h3f71367a;
    11'b01000100000: data <= 32'h38993313;
    11'b01000100001: data <= 32'hb9eebae0;
    11'b01000100010: data <= 32'hbcb7ba64;
    11'b01000100011: data <= 32'hbd93386d;
    11'b01000100100: data <= 32'hbf103c5c;
    11'b01000100101: data <= 32'hbde5b43b;
    11'b01000100110: data <= 32'hb225bed6;
    11'b01000100111: data <= 32'h3a55bc66;
    11'b01000101000: data <= 32'h36083bda;
    11'b01000101001: data <= 32'hb774406e;
    11'b01000101010: data <= 32'hb0133f33;
    11'b01000101011: data <= 32'h3bb43c15;
    11'b01000101100: data <= 32'h3b043a33;
    11'b01000101101: data <= 32'hb8f7368a;
    11'b01000101110: data <= 32'hbd56b866;
    11'b01000101111: data <= 32'h3208bcb1;
    11'b01000110000: data <= 32'h40acb978;
    11'b01000110001: data <= 32'h4135246e;
    11'b01000110010: data <= 32'h3bf6b410;
    11'b01000110011: data <= 32'hb5f1bb24;
    11'b01000110100: data <= 32'hb7a4b748;
    11'b01000110101: data <= 32'hb64b3990;
    11'b01000110110: data <= 32'hbbc63891;
    11'b01000110111: data <= 32'hbd9dbd2c;
    11'b01000111000: data <= 32'hbacfc154;
    11'b01000111001: data <= 32'haad4be65;
    11'b01000111010: data <= 32'hac303a15;
    11'b01000111011: data <= 32'hb6ec3f56;
    11'b01000111100: data <= 32'haeb73c9e;
    11'b01000111101: data <= 32'h3757383f;
    11'b01000111110: data <= 32'hb04f3bb9;
    11'b01000111111: data <= 32'hbe623d5a;
    11'b01001000000: data <= 32'hbf1d38c7;
    11'b01001000001: data <= 32'h332bb712;
    11'b01001000010: data <= 32'h40c7b852;
    11'b01001000011: data <= 32'h40d0a39d;
    11'b01001000100: data <= 32'h3aa22d0f;
    11'b01001000101: data <= 32'h2578ae1d;
    11'b01001000110: data <= 32'h38f035a1;
    11'b01001000111: data <= 32'h3b693bc9;
    11'b01001001000: data <= 32'haf1f33fa;
    11'b01001001001: data <= 32'hbd09bf22;
    11'b01001001010: data <= 32'hbc38c1d4;
    11'b01001001011: data <= 32'ha6e1bede;
    11'b01001001100: data <= 32'h364034a5;
    11'b01001001101: data <= 32'h2dc43a12;
    11'b01001001110: data <= 32'haa89b0d1;
    11'b01001001111: data <= 32'haf0cb4cb;
    11'b01001010000: data <= 32'hbba23bbb;
    11'b01001010001: data <= 32'hc05f3f64;
    11'b01001010010: data <= 32'hc0273bcc;
    11'b01001010011: data <= 32'hb1ceb818;
    11'b01001010100: data <= 32'h3e24ba32;
    11'b01001010101: data <= 32'h3d4a2fb6;
    11'b01001010110: data <= 32'h318b3a63;
    11'b01001010111: data <= 32'h33ba3b1e;
    11'b01001011000: data <= 32'h3de73c60;
    11'b01001011001: data <= 32'h3eec3d30;
    11'b01001011010: data <= 32'h31cc375f;
    11'b01001011011: data <= 32'hbd2cbd31;
    11'b01001011100: data <= 32'hbae6c06d;
    11'b01001011101: data <= 32'h3983bd5d;
    11'b01001011110: data <= 32'h3d77b0d9;
    11'b01001011111: data <= 32'h3a5fb609;
    11'b01001100000: data <= 32'h3060bd31;
    11'b01001100001: data <= 32'hb24abaef;
    11'b01001100010: data <= 32'hbb343b6d;
    11'b01001100011: data <= 32'hbfad3f1d;
    11'b01001100100: data <= 32'hc0043745;
    11'b01001100101: data <= 32'hba50bd41;
    11'b01001100110: data <= 32'h3458bd42;
    11'b01001100111: data <= 32'h22463163;
    11'b01001101000: data <= 32'hb8243cee;
    11'b01001101001: data <= 32'h34303d04;
    11'b01001101010: data <= 32'h3ebc3cd3;
    11'b01001101011: data <= 32'h3e513dd6;
    11'b01001101100: data <= 32'hb5053c7e;
    11'b01001101101: data <= 32'hbe73ad28;
    11'b01001101110: data <= 32'hb8b0bba6;
    11'b01001101111: data <= 32'h3db9b9af;
    11'b01001110000: data <= 32'h4023b586;
    11'b01001110001: data <= 32'h3ca4bb88;
    11'b01001110010: data <= 32'h35f8be69;
    11'b01001110011: data <= 32'h35c1b9fe;
    11'b01001110100: data <= 32'h2ea63c25;
    11'b01001110101: data <= 32'hbb243d81;
    11'b01001110110: data <= 32'hbe60b72b;
    11'b01001110111: data <= 32'hbcf3c06d;
    11'b01001111000: data <= 32'hb931bf24;
    11'b01001111001: data <= 32'hb9ba26a1;
    11'b01001111010: data <= 32'hb9f83ba5;
    11'b01001111011: data <= 32'h332d38d5;
    11'b01001111100: data <= 32'h3d383814;
    11'b01001111101: data <= 32'h39cd3d4d;
    11'b01001111110: data <= 32'hbcdd3f58;
    11'b01001111111: data <= 32'hc0183c85;
    11'b01010000000: data <= 32'hb82b2c84;
    11'b01010000001: data <= 32'h3e2fb451;
    11'b01010000010: data <= 32'h3f77b494;
    11'b01010000011: data <= 32'h3a91b9e2;
    11'b01010000100: data <= 32'h3796bbf1;
    11'b01010000101: data <= 32'h3cfba8fe;
    11'b01010000110: data <= 32'h3de93d45;
    11'b01010000111: data <= 32'h34483c46;
    11'b01010001000: data <= 32'hbc7ebbb1;
    11'b01010001001: data <= 32'hbd45c0ea;
    11'b01010001010: data <= 32'hb9f8bf0f;
    11'b01010001011: data <= 32'hb7a1b235;
    11'b01010001100: data <= 32'hb5a12c9e;
    11'b01010001101: data <= 32'h348bb9fe;
    11'b01010001110: data <= 32'h3a49b8ef;
    11'b01010001111: data <= 32'had513bd9;
    11'b01010010000: data <= 32'hbf314063;
    11'b01010010001: data <= 32'hc07e3e7f;
    11'b01010010010: data <= 32'hb9ca33e7;
    11'b01010010011: data <= 32'h3ae3b563;
    11'b01010010100: data <= 32'h39ebb0ad;
    11'b01010010101: data <= 32'hafabadfa;
    11'b01010010110: data <= 32'h357aaaee;
    11'b01010010111: data <= 32'h3fba398b;
    11'b01010011000: data <= 32'h40c93e52;
    11'b01010011001: data <= 32'h3aa93c82;
    11'b01010011010: data <= 32'hbb93b8f4;
    11'b01010011011: data <= 32'hbc65bee3;
    11'b01010011100: data <= 32'hb00bbc7f;
    11'b01010011101: data <= 32'h36a6b4a4;
    11'b01010011110: data <= 32'h3558bb0d;
    11'b01010011111: data <= 32'h3717c002;
    11'b01010100000: data <= 32'h38c5bdeb;
    11'b01010100001: data <= 32'hb0a83988;
    11'b01010100010: data <= 32'hbe0a4024;
    11'b01010100011: data <= 32'hbfc73cd9;
    11'b01010100100: data <= 32'hbc04b6f9;
    11'b01010100101: data <= 32'hb2febab0;
    11'b01010100110: data <= 32'hb967add6;
    11'b01010100111: data <= 32'hbc80365b;
    11'b01010101000: data <= 32'h2cc8365d;
    11'b01010101001: data <= 32'h401f3a60;
    11'b01010101010: data <= 32'h40b73e31;
    11'b01010101011: data <= 32'h37e73df7;
    11'b01010101100: data <= 32'hbcc936ab;
    11'b01010101101: data <= 32'hba98b5d5;
    11'b01010101110: data <= 32'h390db161;
    11'b01010101111: data <= 32'h3cb5b150;
    11'b01010110000: data <= 32'h399cbd5f;
    11'b01010110001: data <= 32'h383bc0de;
    11'b01010110010: data <= 32'h3b26be3a;
    11'b01010110011: data <= 32'h397d398c;
    11'b01010110100: data <= 32'hb64e3ead;
    11'b01010110101: data <= 32'hbcd23532;
    11'b01010110110: data <= 32'hbc74bd74;
    11'b01010110111: data <= 32'hbc11bd43;
    11'b01010111000: data <= 32'hbe27b004;
    11'b01010111001: data <= 32'hbe5a355a;
    11'b01010111010: data <= 32'haf0cadef;
    11'b01010111011: data <= 32'h3eb02730;
    11'b01010111100: data <= 32'h3e2e3c6a;
    11'b01010111101: data <= 32'hb6773f6f;
    11'b01010111110: data <= 32'hbe8f3df6;
    11'b01010111111: data <= 32'hb97f3a70;
    11'b01011000000: data <= 32'h3b593860;
    11'b01011000001: data <= 32'h3c772d74;
    11'b01011000010: data <= 32'h34edbc74;
    11'b01011000011: data <= 32'h358bbf8f;
    11'b01011000100: data <= 32'h3dc3bb16;
    11'b01011000101: data <= 32'h3fa73bcb;
    11'b01011000110: data <= 32'h3b4c3d44;
    11'b01011000111: data <= 32'hb6d2b521;
    11'b01011001000: data <= 32'hbba8bef1;
    11'b01011001001: data <= 32'hbc4abd0c;
    11'b01011001010: data <= 32'hbd8fae36;
    11'b01011001011: data <= 32'hbd1ab356;
    11'b01011001100: data <= 32'hac81bd2f;
    11'b01011001101: data <= 32'h3c83bcf8;
    11'b01011001110: data <= 32'h392136dd;
    11'b01011001111: data <= 32'hbc653fc4;
    11'b01011010000: data <= 32'hbf4e3fb3;
    11'b01011010001: data <= 32'hb9723c61;
    11'b01011010010: data <= 32'h383738e2;
    11'b01011010011: data <= 32'h307e346b;
    11'b01011010100: data <= 32'hba26b754;
    11'b01011010101: data <= 32'haff3bb20;
    11'b01011010110: data <= 32'h3f4dab94;
    11'b01011010111: data <= 32'h41813cf9;
    11'b01011011000: data <= 32'h3e733cd3;
    11'b01011011001: data <= 32'hac6db3c7;
    11'b01011011010: data <= 32'hb92dbc97;
    11'b01011011011: data <= 32'hb710b7fd;
    11'b01011011100: data <= 32'hb78a3090;
    11'b01011011101: data <= 32'hb82bbaef;
    11'b01011011110: data <= 32'h2ee6c0ed;
    11'b01011011111: data <= 32'h3a7ac084;
    11'b01011100000: data <= 32'h3584adb8;
    11'b01011100001: data <= 32'hbbb03ebc;
    11'b01011100010: data <= 32'hbdb13dfb;
    11'b01011100011: data <= 32'hb91d36b6;
    11'b01011100100: data <= 32'hb36a2ced;
    11'b01011100101: data <= 32'hbcb834fb;
    11'b01011100110: data <= 32'hbfc63013;
    11'b01011100111: data <= 32'hb94eb393;
    11'b01011101000: data <= 32'h3f1a3242;
    11'b01011101001: data <= 32'h41633c8e;
    11'b01011101010: data <= 32'h3d413d19;
    11'b01011101011: data <= 32'hb4f5379b;
    11'b01011101100: data <= 32'hb6152ed9;
    11'b01011101101: data <= 32'h362a3915;
    11'b01011101110: data <= 32'h37593894;
    11'b01011101111: data <= 32'h9de6bc74;
    11'b01011110000: data <= 32'h30dec1b9;
    11'b01011110001: data <= 32'h3ac1c0d1;
    11'b01011110010: data <= 32'h3af3b0a2;
    11'b01011110011: data <= 32'h29933d0f;
    11'b01011110100: data <= 32'hb80c3872;
    11'b01011110101: data <= 32'hb6b5b928;
    11'b01011110110: data <= 32'hba47b853;
    11'b01011110111: data <= 32'hc00334ab;
    11'b01011111000: data <= 32'hc10834a0;
    11'b01011111001: data <= 32'hbba9b6f4;
    11'b01011111010: data <= 32'h3d5db736;
    11'b01011111011: data <= 32'h3f593839;
    11'b01011111100: data <= 32'h34fb3d34;
    11'b01011111101: data <= 32'hbb003d1e;
    11'b01011111110: data <= 32'hb3e33cf2;
    11'b01011111111: data <= 32'h3ae23dfb;
    11'b01100000000: data <= 32'h39613be8;
    11'b01100000001: data <= 32'hb43bba6b;
    11'b01100000010: data <= 32'hb195c091;
    11'b01100000011: data <= 32'h3c38bead;
    11'b01100000100: data <= 32'h3f3d3373;
    11'b01100000101: data <= 32'h3d373b66;
    11'b01100000110: data <= 32'h3726b3e7;
    11'b01100000111: data <= 32'ha9bfbd14;
    11'b01100001000: data <= 32'hb9c7b90f;
    11'b01100001001: data <= 32'hbf5436f9;
    11'b01100001010: data <= 32'hc05929e1;
    11'b01100001011: data <= 32'hbad9bd61;
    11'b01100001100: data <= 32'h3a77beab;
    11'b01100001101: data <= 32'h3a6ab56e;
    11'b01100001110: data <= 32'hb8f03c7b;
    11'b01100001111: data <= 32'hbcdd3e3c;
    11'b01100010000: data <= 32'hb0f13e08;
    11'b01100010001: data <= 32'h3a223e4e;
    11'b01100010010: data <= 32'ha1683ca7;
    11'b01100010011: data <= 32'hbd1ab0bd;
    11'b01100010100: data <= 32'hbac2bcb3;
    11'b01100010101: data <= 32'h3c92b90e;
    11'b01100010110: data <= 32'h40ed394b;
    11'b01100010111: data <= 32'h3ff73a11;
    11'b01100011000: data <= 32'h3af5b712;
    11'b01100011001: data <= 32'h34dabbcb;
    11'b01100011010: data <= 32'haca22a79;
    11'b01100011011: data <= 32'hba9a3af8;
    11'b01100011100: data <= 32'hbcf4b469;
    11'b01100011101: data <= 32'hb82ac09a;
    11'b01100011110: data <= 32'h3759c159;
    11'b01100011111: data <= 32'h3423bbbf;
    11'b01100100000: data <= 32'hba273a21;
    11'b01100100001: data <= 32'hbb4a3c56;
    11'b01100100010: data <= 32'h2c6e3a1b;
    11'b01100100011: data <= 32'h354f3b2f;
    11'b01100100100: data <= 32'hbc683c39;
    11'b01100100101: data <= 32'hc0e33731;
    11'b01100100110: data <= 32'hbe22b4ce;
    11'b01100100111: data <= 32'h3b8cadb8;
    11'b01100101000: data <= 32'h40a8396c;
    11'b01100101001: data <= 32'h3e903954;
    11'b01100101010: data <= 32'h383aaa13;
    11'b01100101011: data <= 32'h374e28bb;
    11'b01100101100: data <= 32'h3a113cb6;
    11'b01100101101: data <= 32'h34cd3ded;
    11'b01100101110: data <= 32'hb712b532;
    11'b01100101111: data <= 32'hb554c132;
    11'b01100110000: data <= 32'h35ccc194;
    11'b01100110001: data <= 32'h3772bbc7;
    11'b01100110010: data <= 32'ha5cc36c0;
    11'b01100110011: data <= 32'ha03e3069;
    11'b01100110100: data <= 32'h37dcb78c;
    11'b01100110101: data <= 32'h245122f6;
    11'b01100110110: data <= 32'hbf373b02;
    11'b01100110111: data <= 32'hc20139b1;
    11'b01100111000: data <= 32'hbf50b237;
    11'b01100111001: data <= 32'h3847b76b;
    11'b01100111010: data <= 32'h3dd22e52;
    11'b01100111011: data <= 32'h37d237b5;
    11'b01100111100: data <= 32'hb48137cb;
    11'b01100111101: data <= 32'h36cb3c15;
    11'b01100111110: data <= 32'h3d3a4015;
    11'b01100111111: data <= 32'h3a693fce;
    11'b01101000000: data <= 32'hb6a92147;
    11'b01101000001: data <= 32'hb8d3bff4;
    11'b01101000010: data <= 32'h35e2bfb2;
    11'b01101000011: data <= 32'h3c76b611;
    11'b01101000100: data <= 32'h3c4933bf;
    11'b01101000101: data <= 32'h3bb6b9c1;
    11'b01101000110: data <= 32'h3bc3bd79;
    11'b01101000111: data <= 32'h30f5b5f3;
    11'b01101001000: data <= 32'hbe553b7d;
    11'b01101001001: data <= 32'hc11f3942;
    11'b01101001010: data <= 32'hbe32ba6a;
    11'b01101001011: data <= 32'h30aebdf8;
    11'b01101001100: data <= 32'h3607ba5a;
    11'b01101001101: data <= 32'hb99030e5;
    11'b01101001110: data <= 32'hbb613921;
    11'b01101001111: data <= 32'h367d3ced;
    11'b01101010000: data <= 32'h3d85401c;
    11'b01101010001: data <= 32'h36ce3ffd;
    11'b01101010010: data <= 32'hbce13861;
    11'b01101010011: data <= 32'hbd2ebabd;
    11'b01101010100: data <= 32'h346eb92e;
    11'b01101010101: data <= 32'h3e65359d;
    11'b01101010110: data <= 32'h3eba32b1;
    11'b01101010111: data <= 32'h3d68bc3c;
    11'b01101011000: data <= 32'h3cfdbd86;
    11'b01101011001: data <= 32'h39cb2d45;
    11'b01101011010: data <= 32'hb8543d85;
    11'b01101011011: data <= 32'hbda13841;
    11'b01101011100: data <= 32'hbb5cbe35;
    11'b01101011101: data <= 32'haab5c0d0;
    11'b01101011110: data <= 32'hb4a8bdac;
    11'b01101011111: data <= 32'hbca0b208;
    11'b01101100000: data <= 32'hbaf3327a;
    11'b01101100001: data <= 32'h38f13736;
    11'b01101100010: data <= 32'h3c973cc0;
    11'b01101100011: data <= 32'hb6ed3e77;
    11'b01101100100: data <= 32'hc08f3be5;
    11'b01101100101: data <= 32'hc001306e;
    11'b01101100110: data <= 32'h285c3287;
    11'b01101100111: data <= 32'h3dcf3924;
    11'b01101101000: data <= 32'h3d2a30f3;
    11'b01101101001: data <= 32'h3ad7baeb;
    11'b01101101010: data <= 32'h3ca4b8fe;
    11'b01101101011: data <= 32'h3d9b3c57;
    11'b01101101100: data <= 32'h3966400d;
    11'b01101101101: data <= 32'hb4e53896;
    11'b01101101110: data <= 32'hb6f4bf2c;
    11'b01101101111: data <= 32'had34c0f5;
    11'b01101110000: data <= 32'hb46dbd36;
    11'b01101110001: data <= 32'hb978b56a;
    11'b01101110010: data <= 32'haf25b8de;
    11'b01101110011: data <= 32'h3c55bae9;
    11'b01101110100: data <= 32'h3bb320a2;
    11'b01101110101: data <= 32'hbc2a3c7f;
    11'b01101110110: data <= 32'hc1943c9b;
    11'b01101110111: data <= 32'hc06f36c9;
    11'b01101111000: data <= 32'hb3692fd3;
    11'b01101111001: data <= 32'h39803397;
    11'b01101111010: data <= 32'h2c53ac77;
    11'b01101111011: data <= 32'hb372b7d6;
    11'b01101111100: data <= 32'h3a803365;
    11'b01101111101: data <= 32'h3f523f99;
    11'b01101111110: data <= 32'h3d5d40e9;
    11'b01101111111: data <= 32'h27243a91;
    11'b01110000000: data <= 32'hb7f7bd0a;
    11'b01110000001: data <= 32'hae75be30;
    11'b01110000010: data <= 32'h3239b74d;
    11'b01110000011: data <= 32'h33f8b2cf;
    11'b01110000100: data <= 32'h3a70bd55;
    11'b01110000101: data <= 32'h3e3dbfa6;
    11'b01110000110: data <= 32'h3c45b993;
    11'b01110000111: data <= 32'hbaea3b8b;
    11'b01110001000: data <= 32'hc0953c64;
    11'b01110001001: data <= 32'hbedd1de6;
    11'b01110001010: data <= 32'hb562b9b6;
    11'b01110001011: data <= 32'hb41bb8b3;
    11'b01110001100: data <= 32'hbd09b6cd;
    11'b01110001101: data <= 32'hbcceb5b1;
    11'b01110001110: data <= 32'h382e373c;
    11'b01110001111: data <= 32'h3f813f76;
    11'b01110010000: data <= 32'h3ca040a3;
    11'b01110010001: data <= 32'hb86e3c6d;
    11'b01110010010: data <= 32'hbc66b3c0;
    11'b01110010011: data <= 32'hb388b056;
    11'b01110010100: data <= 32'h38e338d8;
    11'b01110010101: data <= 32'h3ab12a59;
    11'b01110010110: data <= 32'h3ca1be7b;
    11'b01110010111: data <= 32'h3ecdc03b;
    11'b01110011000: data <= 32'h3db7b7e1;
    11'b01110011001: data <= 32'h2bf03d13;
    11'b01110011010: data <= 32'hbc0d3c14;
    11'b01110011011: data <= 32'hba12b923;
    11'b01110011100: data <= 32'hb32bbe4a;
    11'b01110011101: data <= 32'hbacdbcbb;
    11'b01110011110: data <= 32'hbfa5b96e;
    11'b01110011111: data <= 32'hbdb4b919;
    11'b01110100000: data <= 32'h38abb35e;
    11'b01110100001: data <= 32'h3ebd3b1b;
    11'b01110100010: data <= 32'h36d83e80;
    11'b01110100011: data <= 32'hbe1b3cec;
    11'b01110100100: data <= 32'hbf203930;
    11'b01110100101: data <= 32'hb6f13b43;
    11'b01110100110: data <= 32'h388d3cd1;
    11'b01110100111: data <= 32'h382e31db;
    11'b01110101000: data <= 32'h388dbdd0;
    11'b01110101001: data <= 32'h3d52be09;
    11'b01110101010: data <= 32'h3f333648;
    11'b01110101011: data <= 32'h3cb63f89;
    11'b01110101100: data <= 32'h34743c35;
    11'b01110101101: data <= 32'h2b8abb81;
    11'b01110101110: data <= 32'ha6e7becb;
    11'b01110101111: data <= 32'hbac4bbf9;
    11'b01110110000: data <= 32'hbe6db8ae;
    11'b01110110001: data <= 32'hba8fbca8;
    11'b01110110010: data <= 32'h3c06bdc4;
    11'b01110110011: data <= 32'h3e10b79b;
    11'b01110110100: data <= 32'hb2243a45;
    11'b01110110101: data <= 32'hc0233c89;
    11'b01110110110: data <= 32'hbfc73b64;
    11'b01110110111: data <= 32'hb8033c0a;
    11'b01110111000: data <= 32'h2af33be6;
    11'b01110111001: data <= 32'hb8d025cb;
    11'b01110111010: data <= 32'hb98cbc72;
    11'b01110111011: data <= 32'h3905b971;
    11'b01110111100: data <= 32'h3fc43cde;
    11'b01110111101: data <= 32'h3f414090;
    11'b01110111110: data <= 32'h3a7d3c98;
    11'b01110111111: data <= 32'h333fb8ec;
    11'b01111000000: data <= 32'h2a54badc;
    11'b01111000001: data <= 32'hb6a12160;
    11'b01111000010: data <= 32'hb9e1af2c;
    11'b01111000011: data <= 32'h2d57be5b;
    11'b01111000100: data <= 32'h3dddc0e3;
    11'b01111000101: data <= 32'h3e10bd90;
    11'b01111000110: data <= 32'hb1ee3549;
    11'b01111000111: data <= 32'hbe9d3b90;
    11'b01111001000: data <= 32'hbd353857;
    11'b01111001001: data <= 32'hb4723448;
    11'b01111001010: data <= 32'hb8b73295;
    11'b01111001011: data <= 32'hbf7fb531;
    11'b01111001100: data <= 32'hbf86bb52;
    11'b01111001101: data <= 32'h2780b545;
    11'b01111001110: data <= 32'h3f3f3d0b;
    11'b01111001111: data <= 32'h3ea1400f;
    11'b01111010000: data <= 32'h35a33c8b;
    11'b01111010001: data <= 32'hb4bd2f2c;
    11'b01111010010: data <= 32'haca937e9;
    11'b01111010011: data <= 32'h27713d2f;
    11'b01111010100: data <= 32'hab6837cb;
    11'b01111010101: data <= 32'h380dbea8;
    11'b01111010110: data <= 32'h3e17c154;
    11'b01111010111: data <= 32'h3e78bd59;
    11'b01111011000: data <= 32'h377e3847;
    11'b01111011001: data <= 32'hb6ff3ab4;
    11'b01111011010: data <= 32'hafd4aee7;
    11'b01111011011: data <= 32'h321ab922;
    11'b01111011100: data <= 32'hbb8bb733;
    11'b01111011101: data <= 32'hc111b832;
    11'b01111011110: data <= 32'hc090bbdb;
    11'b01111011111: data <= 32'hacedba1b;
    11'b01111100000: data <= 32'h3e42359d;
    11'b01111100001: data <= 32'h3b843c7e;
    11'b01111100010: data <= 32'hb9143b29;
    11'b01111100011: data <= 32'hbc1439ee;
    11'b01111100100: data <= 32'hb3c53e27;
    11'b01111100101: data <= 32'h30f74032;
    11'b01111100110: data <= 32'hb0df3aad;
    11'b01111100111: data <= 32'ha07cbda4;
    11'b01111101000: data <= 32'h3bb1c027;
    11'b01111101001: data <= 32'h3e85b78c;
    11'b01111101010: data <= 32'h3d3e3cae;
    11'b01111101011: data <= 32'h3acc3adb;
    11'b01111101100: data <= 32'h3b66b83b;
    11'b01111101101: data <= 32'h3930bba4;
    11'b01111101110: data <= 32'hba8ab579;
    11'b01111101111: data <= 32'hc081b450;
    11'b01111110000: data <= 32'hbeedbcb0;
    11'b01111110001: data <= 32'h355ebecb;
    11'b01111110010: data <= 32'h3d8cbc01;
    11'b01111110011: data <= 32'h335c286d;
    11'b01111110100: data <= 32'hbd5637ed;
    11'b01111110101: data <= 32'hbd103ae4;
    11'b01111110110: data <= 32'hb1d53ead;
    11'b01111110111: data <= 32'haafd3fe8;
    11'b01111111000: data <= 32'hbc0739c8;
    11'b01111111001: data <= 32'hbd02bc39;
    11'b01111111010: data <= 32'h1caabcbe;
    11'b01111111011: data <= 32'h3dbe37b1;
    11'b01111111100: data <= 32'h3f093e9a;
    11'b01111111101: data <= 32'h3da73ade;
    11'b01111111110: data <= 32'h3ceab798;
    11'b01111111111: data <= 32'h3a92b5f2;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    