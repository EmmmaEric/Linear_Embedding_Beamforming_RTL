
module memory_rom_30(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hb513be35;
    11'b00000000001: data <= 32'hb333bacf;
    11'b00000000010: data <= 32'h30b83b81;
    11'b00000000011: data <= 32'hb8203f35;
    11'b00000000100: data <= 32'hbea83775;
    11'b00000000101: data <= 32'hbf79bdc0;
    11'b00000000110: data <= 32'hbc6bbdd7;
    11'b00000000111: data <= 32'hb7ec33f4;
    11'b00000001000: data <= 32'hb35f3d57;
    11'b00000001001: data <= 32'h38103a4f;
    11'b00000001010: data <= 32'h3e283187;
    11'b00000001011: data <= 32'h3d973b00;
    11'b00000001100: data <= 32'hb4113fa0;
    11'b00000001101: data <= 32'hbde73e4a;
    11'b00000001110: data <= 32'hb8972dd2;
    11'b00000001111: data <= 32'h3d50bbac;
    11'b00000010000: data <= 32'h3f42bc56;
    11'b00000010001: data <= 32'h3951bc6f;
    11'b00000010010: data <= 32'ha626bce5;
    11'b00000010011: data <= 32'h3a51b8d5;
    11'b00000010100: data <= 32'h3e053965;
    11'b00000010101: data <= 32'h37753c18;
    11'b00000010110: data <= 32'hbdd5b576;
    11'b00000010111: data <= 32'hc06abf3b;
    11'b00000011000: data <= 32'hbdcebde0;
    11'b00000011001: data <= 32'hb89e298e;
    11'b00000011010: data <= 32'hb4743835;
    11'b00000011011: data <= 32'h2d28b606;
    11'b00000011100: data <= 32'h3933b915;
    11'b00000011101: data <= 32'h37333b54;
    11'b00000011110: data <= 32'hba19413d;
    11'b00000011111: data <= 32'hbdf440b3;
    11'b00000100000: data <= 32'hb8793845;
    11'b00000100001: data <= 32'h3b19b9b1;
    11'b00000100010: data <= 32'h3bfdb8ec;
    11'b00000100011: data <= 32'h2f08b433;
    11'b00000100100: data <= 32'h3400b545;
    11'b00000100101: data <= 32'h3f3fb0e0;
    11'b00000100110: data <= 32'h41473862;
    11'b00000100111: data <= 32'h3ca939aa;
    11'b00000101000: data <= 32'hbca6b552;
    11'b00000101001: data <= 32'hbf82bda0;
    11'b00000101010: data <= 32'hba97bcbe;
    11'b00000101011: data <= 32'h2ed6b61b;
    11'b00000101100: data <= 32'ha5e0b92b;
    11'b00000101101: data <= 32'hb482becc;
    11'b00000101110: data <= 32'h1f60bdcd;
    11'b00000101111: data <= 32'h2bbe39bc;
    11'b00000110000: data <= 32'hb9c84132;
    11'b00000110001: data <= 32'hbda44035;
    11'b00000110010: data <= 32'hbc0e3166;
    11'b00000110011: data <= 32'hb39db9cd;
    11'b00000110100: data <= 32'hb4bba461;
    11'b00000110101: data <= 32'hb940394a;
    11'b00000110110: data <= 32'h340535b6;
    11'b00000110111: data <= 32'h406127b3;
    11'b00000111000: data <= 32'h41bc383d;
    11'b00000111001: data <= 32'h3cae3c2d;
    11'b00000111010: data <= 32'hbbc63894;
    11'b00000111011: data <= 32'hbc9cb54d;
    11'b00000111100: data <= 32'h33e4b8ec;
    11'b00000111101: data <= 32'h3b90b91a;
    11'b00000111110: data <= 32'h32f7bda7;
    11'b00000111111: data <= 32'hb69cc0c3;
    11'b00001000000: data <= 32'h2c9ebf2f;
    11'b00001000001: data <= 32'h38f83693;
    11'b00001000010: data <= 32'h27313fac;
    11'b00001000011: data <= 32'hbc6e3c5e;
    11'b00001000100: data <= 32'hbe16b92e;
    11'b00001000101: data <= 32'hbd34bb18;
    11'b00001000110: data <= 32'hbd3335a4;
    11'b00001000111: data <= 32'hbce33bd7;
    11'b00001001000: data <= 32'haa3432a3;
    11'b00001001001: data <= 32'h3ee7b63b;
    11'b00001001010: data <= 32'h403f3746;
    11'b00001001011: data <= 32'h386e3ee1;
    11'b00001001100: data <= 32'hbbb13f2b;
    11'b00001001101: data <= 32'hb81b3a7b;
    11'b00001001110: data <= 32'h3bb5a0ef;
    11'b00001001111: data <= 32'h3ccfb7cb;
    11'b00001010000: data <= 32'h2c52bd26;
    11'b00001010001: data <= 32'hb63ec017;
    11'b00001010010: data <= 32'h3a03be05;
    11'b00001010011: data <= 32'h3f4d31f4;
    11'b00001010100: data <= 32'h3c853c45;
    11'b00001010101: data <= 32'hb90e2d26;
    11'b00001010110: data <= 32'hbe98bcdc;
    11'b00001010111: data <= 32'hbe5abb34;
    11'b00001011000: data <= 32'hbda23636;
    11'b00001011001: data <= 32'hbd1b37f3;
    11'b00001011010: data <= 32'hb763ba5c;
    11'b00001011011: data <= 32'h3a3abd44;
    11'b00001011100: data <= 32'h3c003275;
    11'b00001011101: data <= 32'hb0ac405e;
    11'b00001011110: data <= 32'hbc0240ff;
    11'b00001011111: data <= 32'hb4a03d40;
    11'b00001100000: data <= 32'h3aaf34d3;
    11'b00001100001: data <= 32'h387a1ab3;
    11'b00001100010: data <= 32'hb8c4b648;
    11'b00001100011: data <= 32'hb6bdbc05;
    11'b00001100100: data <= 32'h3dffbb02;
    11'b00001100101: data <= 32'h41c22ecc;
    11'b00001100110: data <= 32'h3fad3896;
    11'b00001100111: data <= 32'hb2e2b2bd;
    11'b00001101000: data <= 32'hbd04bbff;
    11'b00001101001: data <= 32'hbb4eb836;
    11'b00001101010: data <= 32'hb8eb344c;
    11'b00001101011: data <= 32'hbaf8b621;
    11'b00001101100: data <= 32'hba27c00e;
    11'b00001101101: data <= 32'ha2e6c07e;
    11'b00001101110: data <= 32'h3539b179;
    11'b00001101111: data <= 32'hb4e6401c;
    11'b00001110000: data <= 32'hbadf4069;
    11'b00001110001: data <= 32'hb7293b03;
    11'b00001110010: data <= 32'h230b31a4;
    11'b00001110011: data <= 32'hb9183869;
    11'b00001110100: data <= 32'hbdfd393f;
    11'b00001110101: data <= 32'hb91daae4;
    11'b00001110110: data <= 32'h3eedb7b9;
    11'b00001110111: data <= 32'h421e2adf;
    11'b00001111000: data <= 32'h3f93390f;
    11'b00001111001: data <= 32'hadae3622;
    11'b00001111010: data <= 32'hb880a88c;
    11'b00001111011: data <= 32'h3436320c;
    11'b00001111100: data <= 32'h3776344b;
    11'b00001111101: data <= 32'hb6a6bbc2;
    11'b00001111110: data <= 32'hbb3ec155;
    11'b00001111111: data <= 32'hb275c135;
    11'b00010000000: data <= 32'h3895b774;
    11'b00010000001: data <= 32'h35093d88;
    11'b00010000010: data <= 32'hb69d3c66;
    11'b00010000011: data <= 32'hb963b0ff;
    11'b00010000100: data <= 32'hbab8b23f;
    11'b00010000101: data <= 32'hbe653b3a;
    11'b00010000110: data <= 32'hc03d3ccf;
    11'b00010000111: data <= 32'hbbe02f18;
    11'b00010001000: data <= 32'h3cfaba00;
    11'b00010001001: data <= 32'h4077b0c5;
    11'b00010001010: data <= 32'h3c5e3c0d;
    11'b00010001011: data <= 32'hb45c3d79;
    11'b00010001100: data <= 32'h29dd3c40;
    11'b00010001101: data <= 32'h3cbd3b22;
    11'b00010001110: data <= 32'h3c23382d;
    11'b00010001111: data <= 32'hb641ba54;
    11'b00010010000: data <= 32'hbbe4c085;
    11'b00010010001: data <= 32'h31d3c055;
    11'b00010010010: data <= 32'h3e16b830;
    11'b00010010011: data <= 32'h3d78388a;
    11'b00010010100: data <= 32'h321bae47;
    11'b00010010101: data <= 32'hb927bc1f;
    11'b00010010110: data <= 32'hbc29b676;
    11'b00010010111: data <= 32'hbe9e3c10;
    11'b00010011000: data <= 32'hc0263c07;
    11'b00010011001: data <= 32'hbd13b8f5;
    11'b00010011010: data <= 32'h353fbe75;
    11'b00010011011: data <= 32'h3b88b863;
    11'b00010011100: data <= 32'h2e0a3d1b;
    11'b00010011101: data <= 32'hb8313fd5;
    11'b00010011110: data <= 32'h35203e1c;
    11'b00010011111: data <= 32'h3d583ca0;
    11'b00010100000: data <= 32'h396c3b74;
    11'b00010100001: data <= 32'hbbca2d74;
    11'b00010100010: data <= 32'hbcadbc4a;
    11'b00010100011: data <= 32'h3994bd06;
    11'b00010100100: data <= 32'h40dcb621;
    11'b00010100101: data <= 32'h404329f7;
    11'b00010100110: data <= 32'h38e8b941;
    11'b00010100111: data <= 32'hb469bc76;
    11'b00010101000: data <= 32'hb5dcb048;
    11'b00010101001: data <= 32'hb9dd3c2d;
    11'b00010101010: data <= 32'hbda9361b;
    11'b00010101011: data <= 32'hbd6fbebd;
    11'b00010101100: data <= 32'hb78cc10d;
    11'b00010101101: data <= 32'h2199bbcc;
    11'b00010101110: data <= 32'hb61d3c79;
    11'b00010101111: data <= 32'hb81c3e91;
    11'b00010110000: data <= 32'h34c23be3;
    11'b00010110001: data <= 32'h3a443a86;
    11'b00010110010: data <= 32'hb5403d1d;
    11'b00010110011: data <= 32'hbf713c84;
    11'b00010110100: data <= 32'hbdec2fd6;
    11'b00010110101: data <= 32'h3acab848;
    11'b00010110110: data <= 32'h4122b45b;
    11'b00010110111: data <= 32'h400ba177;
    11'b00010111000: data <= 32'h3891b579;
    11'b00010111001: data <= 32'h33ddb5db;
    11'b00010111010: data <= 32'h3a6c3882;
    11'b00010111011: data <= 32'h389a3cab;
    11'b00010111100: data <= 32'hb907ad16;
    11'b00010111101: data <= 32'hbd37c084;
    11'b00010111110: data <= 32'hba05c1a7;
    11'b00010111111: data <= 32'ha708bc9c;
    11'b00011000000: data <= 32'h991f389d;
    11'b00011000001: data <= 32'hae743851;
    11'b00011000010: data <= 32'h32e0b41a;
    11'b00011000011: data <= 32'h2df92fb5;
    11'b00011000100: data <= 32'hbcd63db1;
    11'b00011000101: data <= 32'hc0e73efc;
    11'b00011000110: data <= 32'hbf0d3897;
    11'b00011000111: data <= 32'h372bb842;
    11'b00011001000: data <= 32'h3ef1b6ad;
    11'b00011001001: data <= 32'h3c203307;
    11'b00011001010: data <= 32'h2d363723;
    11'b00011001011: data <= 32'h3921390e;
    11'b00011001100: data <= 32'h3f1c3d07;
    11'b00011001101: data <= 32'h3db83da6;
    11'b00011001110: data <= 32'hb4ea2b6e;
    11'b00011001111: data <= 32'hbd2fbf5e;
    11'b00011010000: data <= 32'hb820c074;
    11'b00011010001: data <= 32'h3996bb76;
    11'b00011010010: data <= 32'h3b67a820;
    11'b00011010011: data <= 32'h3811b99c;
    11'b00011010100: data <= 32'h348fbda9;
    11'b00011010101: data <= 32'hae8ab684;
    11'b00011010110: data <= 32'hbcfd3da8;
    11'b00011010111: data <= 32'hc08e3ebf;
    11'b00011011000: data <= 32'hbf3c2d92;
    11'b00011011001: data <= 32'hb471bcfa;
    11'b00011011010: data <= 32'h3685ba97;
    11'b00011011011: data <= 32'hb3e23670;
    11'b00011011100: data <= 32'hb80c3be4;
    11'b00011011101: data <= 32'h3a223c48;
    11'b00011011110: data <= 32'h401a3db8;
    11'b00011011111: data <= 32'h3d563e89;
    11'b00011100000: data <= 32'hb9a73a26;
    11'b00011100001: data <= 32'hbde8b8fa;
    11'b00011100010: data <= 32'haef0bc2f;
    11'b00011100011: data <= 32'h3e11b729;
    11'b00011100100: data <= 32'h3e9db618;
    11'b00011100101: data <= 32'h3b00bd7d;
    11'b00011100110: data <= 32'h382bbf1e;
    11'b00011100111: data <= 32'h3706b5ab;
    11'b00011101000: data <= 32'hb4cb3db1;
    11'b00011101001: data <= 32'hbd783cbd;
    11'b00011101010: data <= 32'hbe3bbad6;
    11'b00011101011: data <= 32'hbb1ec037;
    11'b00011101100: data <= 32'hb900bce6;
    11'b00011101101: data <= 32'hbc133523;
    11'b00011101110: data <= 32'hb9fe3a1f;
    11'b00011101111: data <= 32'h3998380f;
    11'b00011110000: data <= 32'h3e873af2;
    11'b00011110001: data <= 32'h37b63ea3;
    11'b00011110010: data <= 32'hbe1d3e7a;
    11'b00011110011: data <= 32'hbf233952;
    11'b00011110100: data <= 32'h2c83a3a1;
    11'b00011110101: data <= 32'h3ed8aa0d;
    11'b00011110110: data <= 32'h3e1cb5d8;
    11'b00011110111: data <= 32'h392fbcc7;
    11'b00011111000: data <= 32'h3a07bcdb;
    11'b00011111001: data <= 32'h3daf3416;
    11'b00011111010: data <= 32'h3c5e3e39;
    11'b00011111011: data <= 32'hb43839e8;
    11'b00011111100: data <= 32'hbcbbbdce;
    11'b00011111101: data <= 32'hbc45c0ca;
    11'b00011111110: data <= 32'hba6dbd07;
    11'b00011111111: data <= 32'hbadb26bc;
    11'b00100000000: data <= 32'hb746b146;
    11'b00100000001: data <= 32'h390aba7a;
    11'b00100000010: data <= 32'h3befb07f;
    11'b00100000011: data <= 32'hb63a3dda;
    11'b00100000100: data <= 32'hc0384036;
    11'b00100000101: data <= 32'hbfda3d04;
    11'b00100000110: data <= 32'hb02a33a3;
    11'b00100000111: data <= 32'h3c20a86a;
    11'b00100001000: data <= 32'h3785b07b;
    11'b00100001001: data <= 32'hb089b7c3;
    11'b00100001010: data <= 32'h3a6db425;
    11'b00100001011: data <= 32'h407e3b85;
    11'b00100001100: data <= 32'h402a3ef2;
    11'b00100001101: data <= 32'h356b39cb;
    11'b00100001110: data <= 32'hbbcabca8;
    11'b00100001111: data <= 32'hba89bef5;
    11'b00100010000: data <= 32'hb1afba13;
    11'b00100010001: data <= 32'h9f86b3d4;
    11'b00100010010: data <= 32'h306bbcfe;
    11'b00100010011: data <= 32'h395ac035;
    11'b00100010100: data <= 32'h398abbcd;
    11'b00100010101: data <= 32'hb8463cd8;
    11'b00100010110: data <= 32'hbf964005;
    11'b00100010111: data <= 32'hbf0d3b12;
    11'b00100011000: data <= 32'hb84ab5b5;
    11'b00100011001: data <= 32'hb06bb67f;
    11'b00100011010: data <= 32'hbb882a54;
    11'b00100011011: data <= 32'hbc392f4a;
    11'b00100011100: data <= 32'h3931343a;
    11'b00100011101: data <= 32'h40eb3c5e;
    11'b00100011110: data <= 32'h403b3f03;
    11'b00100011111: data <= 32'h2e193c93;
    11'b00100100000: data <= 32'hbc5dae6a;
    11'b00100100001: data <= 32'hb69fb6e5;
    11'b00100100010: data <= 32'h39482c0c;
    11'b00100100011: data <= 32'h3a3ab491;
    11'b00100100100: data <= 32'h3801bf5a;
    11'b00100100101: data <= 32'h39f8c137;
    11'b00100100110: data <= 32'h3bd4bc7a;
    11'b00100100111: data <= 32'h34333c7a;
    11'b00100101000: data <= 32'hbaf53e0c;
    11'b00100101001: data <= 32'hbcb2a9bc;
    11'b00100101010: data <= 32'hba92bd00;
    11'b00100101011: data <= 32'hbc4bba7e;
    11'b00100101100: data <= 32'hbf7a2d56;
    11'b00100101101: data <= 32'hbe262ed3;
    11'b00100101110: data <= 32'h370db104;
    11'b00100101111: data <= 32'h401336ee;
    11'b00100110000: data <= 32'h3d383dd2;
    11'b00100110001: data <= 32'hb9cc3ea4;
    11'b00100110010: data <= 32'hbd9e3c50;
    11'b00100110011: data <= 32'hb1043a23;
    11'b00100110100: data <= 32'h3c1b39f4;
    11'b00100110101: data <= 32'h3a46ad82;
    11'b00100110110: data <= 32'h3265be97;
    11'b00100110111: data <= 32'h3979c039;
    11'b00100111000: data <= 32'h3e88b860;
    11'b00100111001: data <= 32'h3e253d00;
    11'b00100111010: data <= 32'h36803c0f;
    11'b00100111011: data <= 32'hb7bfba34;
    11'b00100111100: data <= 32'hba30bea1;
    11'b00100111101: data <= 32'hbce7ba5d;
    11'b00100111110: data <= 32'hbf3729f4;
    11'b00100111111: data <= 32'hbd4cb81c;
    11'b00101000000: data <= 32'h359fbd67;
    11'b00101000001: data <= 32'h3d78b9f8;
    11'b00101000010: data <= 32'h35573b5e;
    11'b00101000011: data <= 32'hbda73f8a;
    11'b00101000100: data <= 32'hbe3a3e83;
    11'b00101000101: data <= 32'hb0773c96;
    11'b00101000110: data <= 32'h39103b19;
    11'b00101000111: data <= 32'hb0b83203;
    11'b00101001000: data <= 32'hba03bb5d;
    11'b00101001001: data <= 32'h362dbc5d;
    11'b00101001010: data <= 32'h40583359;
    11'b00101001011: data <= 32'h40f33db4;
    11'b00101001100: data <= 32'h3ca43a96;
    11'b00101001101: data <= 32'hadd5b9fb;
    11'b00101001110: data <= 32'hb6fbbc84;
    11'b00101001111: data <= 32'hb8b6b0e1;
    11'b00101010000: data <= 32'hbb642f9c;
    11'b00101010001: data <= 32'hb94ebd2e;
    11'b00101010010: data <= 32'h3667c12a;
    11'b00101010011: data <= 32'h3b6cbf05;
    11'b00101010100: data <= 32'ha99536f8;
    11'b00101010101: data <= 32'hbd543ea3;
    11'b00101010110: data <= 32'hbcf13cfb;
    11'b00101010111: data <= 32'hb2f73876;
    11'b00101011000: data <= 32'hb36737b4;
    11'b00101011001: data <= 32'hbdf735d6;
    11'b00101011010: data <= 32'hbf6db2e7;
    11'b00101011011: data <= 32'ha9afb5d0;
    11'b00101011100: data <= 32'h406e3827;
    11'b00101011101: data <= 32'h40fc3d67;
    11'b00101011110: data <= 32'h3bb13b83;
    11'b00101011111: data <= 32'hb25d22e7;
    11'b00101100000: data <= 32'ha8892ec0;
    11'b00101100001: data <= 32'h353e3af8;
    11'b00101100010: data <= 32'h28993634;
    11'b00101100011: data <= 32'hb12dbeba;
    11'b00101100100: data <= 32'h36afc225;
    11'b00101100101: data <= 32'h3b8bbfec;
    11'b00101100110: data <= 32'h3752348c;
    11'b00101100111: data <= 32'hb63c3c92;
    11'b00101101000: data <= 32'hb721341d;
    11'b00101101001: data <= 32'hb16fb7a3;
    11'b00101101010: data <= 32'hbb7eab3c;
    11'b00101101011: data <= 32'hc0ce36de;
    11'b00101101100: data <= 32'hc0eb222d;
    11'b00101101101: data <= 32'hb5d7b7fe;
    11'b00101101110: data <= 32'h3efaa95c;
    11'b00101101111: data <= 32'h3e8a3ae9;
    11'b00101110000: data <= 32'h28553c73;
    11'b00101110001: data <= 32'hb9083b85;
    11'b00101110010: data <= 32'h336d3d27;
    11'b00101110011: data <= 32'h3b273ed8;
    11'b00101110100: data <= 32'h34fb3a08;
    11'b00101110101: data <= 32'hb591bda6;
    11'b00101110110: data <= 32'h3215c114;
    11'b00101110111: data <= 32'h3d06bd5a;
    11'b00101111000: data <= 32'h3ddc380d;
    11'b00101111001: data <= 32'h3af23928;
    11'b00101111010: data <= 32'h36f7b924;
    11'b00101111011: data <= 32'h2e30bc8c;
    11'b00101111100: data <= 32'hbbd0b16d;
    11'b00101111101: data <= 32'hc0a13839;
    11'b00101111110: data <= 32'hc06fb484;
    11'b00101111111: data <= 32'hb65ebdac;
    11'b00110000000: data <= 32'h3c4abcc7;
    11'b00110000001: data <= 32'h38292f89;
    11'b00110000010: data <= 32'hbb1e3c4b;
    11'b00110000011: data <= 32'hbb613d63;
    11'b00110000100: data <= 32'h35a73ea2;
    11'b00110000101: data <= 32'h3a703f81;
    11'b00110000110: data <= 32'hb5763c10;
    11'b00110000111: data <= 32'hbd0ab967;
    11'b00110001000: data <= 32'hb53cbd97;
    11'b00110001001: data <= 32'h3dfeb592;
    11'b00110001010: data <= 32'h40763aa3;
    11'b00110001011: data <= 32'h3e80360a;
    11'b00110001100: data <= 32'h3b36bb2a;
    11'b00110001101: data <= 32'h3799bb1e;
    11'b00110001110: data <= 32'hb50a36b0;
    11'b00110001111: data <= 32'hbd593a84;
    11'b00110010000: data <= 32'hbd7cb9fd;
    11'b00110010001: data <= 32'hb27fc0e9;
    11'b00110010010: data <= 32'h38aac06d;
    11'b00110010011: data <= 32'haf5cb7d3;
    11'b00110010100: data <= 32'hbc5c3a00;
    11'b00110010101: data <= 32'hb9693b57;
    11'b00110010110: data <= 32'h379c3bf5;
    11'b00110010111: data <= 32'h34383d4a;
    11'b00110011000: data <= 32'hbde63c3d;
    11'b00110011001: data <= 32'hc0c32bd2;
    11'b00110011010: data <= 32'hbb5cb6f8;
    11'b00110011011: data <= 32'h3d90332a;
    11'b00110011100: data <= 32'h405b3ad5;
    11'b00110011101: data <= 32'h3d7f3507;
    11'b00110011110: data <= 32'h398bb757;
    11'b00110011111: data <= 32'h3a2a2fb5;
    11'b00110100000: data <= 32'h38fd3dd5;
    11'b00110100001: data <= 32'hb1533d1c;
    11'b00110100010: data <= 32'hb8bbbb81;
    11'b00110100011: data <= 32'habdec1b3;
    11'b00110100100: data <= 32'h3725c0d2;
    11'b00110100101: data <= 32'h2c3fb8bc;
    11'b00110100110: data <= 32'hb63434c8;
    11'b00110100111: data <= 32'h2fd3adf4;
    11'b00110101000: data <= 32'h39e8b341;
    11'b00110101001: data <= 32'hb2a13823;
    11'b00110101010: data <= 32'hc08b3bdb;
    11'b00110101011: data <= 32'hc1f53693;
    11'b00110101100: data <= 32'hbcfcb42d;
    11'b00110101101: data <= 32'h3b84ad20;
    11'b00110101110: data <= 32'h3d293600;
    11'b00110101111: data <= 32'h348f3438;
    11'b00110110000: data <= 32'h24713284;
    11'b00110110001: data <= 32'h3b1a3cb1;
    11'b00110110010: data <= 32'h3d2540a1;
    11'b00110110011: data <= 32'h36833ed0;
    11'b00110110100: data <= 32'hb809b91c;
    11'b00110110101: data <= 32'hb418c08e;
    11'b00110110110: data <= 32'h3851be89;
    11'b00110110111: data <= 32'h3a4cb0f6;
    11'b00110111000: data <= 32'h39c7aae5;
    11'b00110111001: data <= 32'h3c28bc47;
    11'b00110111010: data <= 32'h3c77bcae;
    11'b00110111011: data <= 32'hb1712f8a;
    11'b00110111100: data <= 32'hc0453c12;
    11'b00110111101: data <= 32'hc1443528;
    11'b00110111110: data <= 32'hbc6bbb09;
    11'b00110111111: data <= 32'h3659bc42;
    11'b00111000000: data <= 32'h2f0cb6a9;
    11'b00111000001: data <= 32'hbb432c68;
    11'b00111000010: data <= 32'hb89037ca;
    11'b00111000011: data <= 32'h3b593df0;
    11'b00111000100: data <= 32'h3d8740d3;
    11'b00111000101: data <= 32'h2bf23f5c;
    11'b00111000110: data <= 32'hbce89da2;
    11'b00111000111: data <= 32'hba85bc4f;
    11'b00111001000: data <= 32'h38c1b641;
    11'b00111001001: data <= 32'h3d8e376c;
    11'b00111001010: data <= 32'h3da5b2a5;
    11'b00111001011: data <= 32'h3de6bdf3;
    11'b00111001100: data <= 32'h3db5bcf0;
    11'b00111001101: data <= 32'h36c337de;
    11'b00111001110: data <= 32'hbc693d55;
    11'b00111001111: data <= 32'hbe392be5;
    11'b00111010000: data <= 32'hb8f7bedf;
    11'b00111010001: data <= 32'h28a5c002;
    11'b00111010010: data <= 32'hb960bc1b;
    11'b00111010011: data <= 32'hbdb2b3df;
    11'b00111010100: data <= 32'hb8812d83;
    11'b00111010101: data <= 32'h3c323a2b;
    11'b00111010110: data <= 32'h3c363ea1;
    11'b00111010111: data <= 32'hbac13e75;
    11'b00111011000: data <= 32'hc08238c2;
    11'b00111011001: data <= 32'hbdc123f0;
    11'b00111011010: data <= 32'h370437fe;
    11'b00111011011: data <= 32'h3d493a05;
    11'b00111011100: data <= 32'h3c73b40e;
    11'b00111011101: data <= 32'h3c69bd0c;
    11'b00111011110: data <= 32'h3df2b792;
    11'b00111011111: data <= 32'h3cea3db1;
    11'b00111100000: data <= 32'h31e53f61;
    11'b00111100001: data <= 32'hb756a822;
    11'b00111100010: data <= 32'hb21dc01d;
    11'b00111100011: data <= 32'haafac050;
    11'b00111100100: data <= 32'hb993bc08;
    11'b00111100101: data <= 32'hbbeeb80e;
    11'b00111100110: data <= 32'h2eceba75;
    11'b00111100111: data <= 32'h3d79b870;
    11'b00111101000: data <= 32'h39b9385a;
    11'b00111101001: data <= 32'hbe343cee;
    11'b00111101010: data <= 32'hc19d3af8;
    11'b00111101011: data <= 32'hbebf3634;
    11'b00111101100: data <= 32'h2ffd37cb;
    11'b00111101101: data <= 32'h383636e7;
    11'b00111101110: data <= 32'hac81b5bf;
    11'b00111101111: data <= 32'h3060ba19;
    11'b00111110000: data <= 32'h3d2e374e;
    11'b00111110001: data <= 32'h3f2e4079;
    11'b00111110010: data <= 32'h3b8f4078;
    11'b00111110011: data <= 32'haba531e1;
    11'b00111110100: data <= 32'hb232be32;
    11'b00111110101: data <= 32'h9ae3bd2d;
    11'b00111110110: data <= 32'hb11bb4e8;
    11'b00111110111: data <= 32'ha86fb87f;
    11'b00111111000: data <= 32'h3bd3beb4;
    11'b00111111001: data <= 32'h3effbeb3;
    11'b00111111010: data <= 32'h39c9b1db;
    11'b00111111011: data <= 32'hbdcc3c29;
    11'b00111111100: data <= 32'hc0c73a6a;
    11'b00111111101: data <= 32'hbd42a856;
    11'b00111111110: data <= 32'hb094b503;
    11'b00111111111: data <= 32'hb85bb4de;
    11'b01000000000: data <= 32'hbdb9b8b3;
    11'b01000000001: data <= 32'hba4fb7ff;
    11'b01000000010: data <= 32'h3c443a34;
    11'b01000000011: data <= 32'h3f89408e;
    11'b01000000100: data <= 32'h3a6c405d;
    11'b01000000101: data <= 32'hb886389a;
    11'b01000000110: data <= 32'hb96ab739;
    11'b01000000111: data <= 32'h93af2ef6;
    11'b01000001000: data <= 32'h3606393b;
    11'b01000001001: data <= 32'h3910b6ec;
    11'b01000001010: data <= 32'h3d7fc020;
    11'b01000001011: data <= 32'h3fadbfc8;
    11'b01000001100: data <= 32'h3c76ab43;
    11'b01000001101: data <= 32'hb8153d01;
    11'b01000001110: data <= 32'hbca738cb;
    11'b01000001111: data <= 32'hb7e4ba27;
    11'b01000010000: data <= 32'hb293bccf;
    11'b01000010001: data <= 32'hbd1cbb1c;
    11'b01000010010: data <= 32'hc050ba80;
    11'b01000010011: data <= 32'hbc3db9fd;
    11'b01000010100: data <= 32'h3c3c308e;
    11'b01000010101: data <= 32'h3e6f3d90;
    11'b01000010110: data <= 32'h27063e8b;
    11'b01000010111: data <= 32'hbe0c3afd;
    11'b01000011000: data <= 32'hbd1e38a2;
    11'b01000011001: data <= 32'haf3b3cd9;
    11'b01000011010: data <= 32'h36903d01;
    11'b01000011011: data <= 32'h3662b4da;
    11'b01000011100: data <= 32'h3b24bf84;
    11'b01000011101: data <= 32'h3ec0bd59;
    11'b01000011110: data <= 32'h3e833a19;
    11'b01000011111: data <= 32'h39a43ef5;
    11'b01000100000: data <= 32'h30c437f7;
    11'b01000100001: data <= 32'h345dbca6;
    11'b01000100010: data <= 32'had67bd9a;
    11'b01000100011: data <= 32'hbd51ba49;
    11'b01000100100: data <= 32'hbf97ba98;
    11'b01000100101: data <= 32'hb84abd7a;
    11'b01000100110: data <= 32'h3d5fbc6e;
    11'b01000100111: data <= 32'h3d282c42;
    11'b01000101000: data <= 32'hb9883b2f;
    11'b01000101001: data <= 32'hc0303b3c;
    11'b01000101010: data <= 32'hbddf3bb3;
    11'b01000101011: data <= 32'hb32f3d93;
    11'b01000101100: data <= 32'hb0a53c76;
    11'b01000101101: data <= 32'hb9adb5a8;
    11'b01000101110: data <= 32'hb45fbda9;
    11'b01000101111: data <= 32'h3c8ab6e8;
    11'b01000110000: data <= 32'h3fb23e59;
    11'b01000110001: data <= 32'h3dd8402f;
    11'b01000110010: data <= 32'h3a17387a;
    11'b01000110011: data <= 32'h37fabada;
    11'b01000110100: data <= 32'h2ab6b8df;
    11'b01000110101: data <= 32'hbab12e48;
    11'b01000110110: data <= 32'hbbffb834;
    11'b01000110111: data <= 32'h3532bfd2;
    11'b01000111000: data <= 32'h3ed1c06c;
    11'b01000111001: data <= 32'h3cc1bb1e;
    11'b01000111010: data <= 32'hba0936f2;
    11'b01000111011: data <= 32'hbef939b2;
    11'b01000111100: data <= 32'hbb7d38b2;
    11'b01000111101: data <= 32'hb119397e;
    11'b01000111110: data <= 32'hbb7636ae;
    11'b01000111111: data <= 32'hc017b895;
    11'b01001000000: data <= 32'hbdc1bc58;
    11'b01001000001: data <= 32'h38c523c5;
    11'b01001000010: data <= 32'h3f673ec4;
    11'b01001000011: data <= 32'h3d713fa2;
    11'b01001000100: data <= 32'h361a3931;
    11'b01001000101: data <= 32'h2dc2a829;
    11'b01001000110: data <= 32'h2c283a1d;
    11'b01001000111: data <= 32'hb4503d38;
    11'b01001001000: data <= 32'hb3b2ab44;
    11'b01001001001: data <= 32'h3a44c04a;
    11'b01001001010: data <= 32'h3f1bc108;
    11'b01001001011: data <= 32'h3d45bb5f;
    11'b01001001100: data <= 32'haca33836;
    11'b01001001101: data <= 32'hb86737c0;
    11'b01001001110: data <= 32'h3029b0e7;
    11'b01001001111: data <= 32'h3059b41d;
    11'b01001010000: data <= 32'hbdc5b322;
    11'b01001010001: data <= 32'hc199b9df;
    11'b01001010010: data <= 32'hbf98bc75;
    11'b01001010011: data <= 32'h36c2b61c;
    11'b01001010100: data <= 32'h3e193ac6;
    11'b01001010101: data <= 32'h38c73c83;
    11'b01001010110: data <= 32'hb8aa38a9;
    11'b01001010111: data <= 32'hb8703a0e;
    11'b01001011000: data <= 32'ha17e3f93;
    11'b01001011001: data <= 32'habf6403e;
    11'b01001011010: data <= 32'hb4363493;
    11'b01001011011: data <= 32'h35a8bf87;
    11'b01001011100: data <= 32'h3d56bfb8;
    11'b01001011101: data <= 32'h3de3afb4;
    11'b01001011110: data <= 32'h3b223c23;
    11'b01001011111: data <= 32'h3a4935d3;
    11'b01001100000: data <= 32'h3c91b96b;
    11'b01001100001: data <= 32'h3822b91c;
    11'b01001100010: data <= 32'hbd89b1d1;
    11'b01001100011: data <= 32'hc124b887;
    11'b01001100100: data <= 32'hbdb9bd97;
    11'b01001100101: data <= 32'h3992bd82;
    11'b01001100110: data <= 32'h3cc6b7f4;
    11'b01001100111: data <= 32'hb2fa2ff0;
    11'b01001101000: data <= 32'hbd4834ff;
    11'b01001101001: data <= 32'hba813bff;
    11'b01001101010: data <= 32'h2572403b;
    11'b01001101011: data <= 32'hb4f5402a;
    11'b01001101100: data <= 32'hbc7b348d;
    11'b01001101101: data <= 32'hba95bd9b;
    11'b01001101110: data <= 32'h380ebba7;
    11'b01001101111: data <= 32'h3dbc3aa9;
    11'b01001110000: data <= 32'h3deb3dd8;
    11'b01001110001: data <= 32'h3dca3516;
    11'b01001110010: data <= 32'h3e0bb926;
    11'b01001110011: data <= 32'h39fdadc0;
    11'b01001110100: data <= 32'hbae7399a;
    11'b01001110101: data <= 32'hbe85159a;
    11'b01001110110: data <= 32'hb789be87;
    11'b01001110111: data <= 32'h3c86c094;
    11'b01001111000: data <= 32'h3c0fbe09;
    11'b01001111001: data <= 32'hb822b839;
    11'b01001111010: data <= 32'hbccda713;
    11'b01001111011: data <= 32'hb4c4389d;
    11'b01001111100: data <= 32'h356a3d8e;
    11'b01001111101: data <= 32'hb9f23d49;
    11'b01001111110: data <= 32'hc07f1580;
    11'b01001111111: data <= 32'hc019bc14;
    11'b01010000000: data <= 32'hb425b4eb;
    11'b01010000001: data <= 32'h3ca53ca0;
    11'b01010000010: data <= 32'h3d3a3d40;
    11'b01010000011: data <= 32'h3c4831c1;
    11'b01010000100: data <= 32'h3c54b14d;
    11'b01010000101: data <= 32'h39c03c47;
    11'b01010000110: data <= 32'hb42d3fdf;
    11'b01010000111: data <= 32'hb99c39d1;
    11'b01010001000: data <= 32'h323fbe4e;
    11'b01010001001: data <= 32'h3d08c0fe;
    11'b01010001010: data <= 32'h3b94be42;
    11'b01010001011: data <= 32'hb14eb76f;
    11'b01010001100: data <= 32'hb345b3e6;
    11'b01010001101: data <= 32'h3a9bb21c;
    11'b01010001110: data <= 32'h3b4834eb;
    11'b01010001111: data <= 32'hbbc437d6;
    11'b01010010000: data <= 32'hc1c5b372;
    11'b01010010001: data <= 32'hc11abb1a;
    11'b01010010010: data <= 32'hb81cb64c;
    11'b01010010011: data <= 32'h3a663849;
    11'b01010010100: data <= 32'h381b37c2;
    11'b01010010101: data <= 32'h97ffb17c;
    11'b01010010110: data <= 32'h3451350b;
    11'b01010010111: data <= 32'h38794021;
    11'b01010011000: data <= 32'h2ca441b1;
    11'b01010011001: data <= 32'hb6fe3ccf;
    11'b01010011010: data <= 32'h9d54bcea;
    11'b01010011011: data <= 32'h3a4bbf7b;
    11'b01010011100: data <= 32'h3a91b979;
    11'b01010011101: data <= 32'h379231b2;
    11'b01010011110: data <= 32'h3bb1b48c;
    11'b01010011111: data <= 32'h3facba7f;
    11'b01010100000: data <= 32'h3de3b55c;
    11'b01010100001: data <= 32'hba3d34c2;
    11'b01010100010: data <= 32'hc136abfc;
    11'b01010100011: data <= 32'hc011bb42;
    11'b01010100100: data <= 32'hb09dbc39;
    11'b01010100101: data <= 32'h384db92d;
    11'b01010100110: data <= 32'hb60fb8e6;
    11'b01010100111: data <= 32'hbbcbb955;
    11'b01010101000: data <= 32'hb3193616;
    11'b01010101001: data <= 32'h38864072;
    11'b01010101010: data <= 32'h2bf84194;
    11'b01010101011: data <= 32'hbbb33c9b;
    11'b01010101100: data <= 32'hbc07ba5a;
    11'b01010101101: data <= 32'hb054baa9;
    11'b01010101110: data <= 32'h383337a7;
    11'b01010101111: data <= 32'h3abd3aa9;
    11'b01010110000: data <= 32'h3e32b47e;
    11'b01010110001: data <= 32'h409bbbe2;
    11'b01010110010: data <= 32'h3ed6af08;
    11'b01010110011: data <= 32'hb45d3beb;
    11'b01010110100: data <= 32'hbe6c38bb;
    11'b01010110101: data <= 32'hbb1ebae9;
    11'b01010110110: data <= 32'h380ebedc;
    11'b01010110111: data <= 32'h36d3be4d;
    11'b01010111000: data <= 32'hbad9bd43;
    11'b01010111001: data <= 32'hbcabbc48;
    11'b01010111010: data <= 32'h2db7ac5b;
    11'b01010111011: data <= 32'h3b9d3dc4;
    11'b01010111100: data <= 32'hada93f80;
    11'b01010111101: data <= 32'hbf413960;
    11'b01010111110: data <= 32'hc046b7d5;
    11'b01010111111: data <= 32'hbbdba797;
    11'b01011000000: data <= 32'h302d3c6a;
    11'b01011000001: data <= 32'h38ce3b39;
    11'b01011000010: data <= 32'h3c7bb76d;
    11'b01011000011: data <= 32'h3f08ba45;
    11'b01011000100: data <= 32'h3e0e3a0d;
    11'b01011000101: data <= 32'h340b404c;
    11'b01011000110: data <= 32'hb85b3dac;
    11'b01011000111: data <= 32'h2c44b915;
    11'b01011001000: data <= 32'h3af0bf3d;
    11'b01011001001: data <= 32'h3574be50;
    11'b01011001010: data <= 32'hba26bcb6;
    11'b01011001011: data <= 32'hb7f0bcad;
    11'b01011001100: data <= 32'h3c5eba2b;
    11'b01011001101: data <= 32'h3e8b33dd;
    11'b01011001110: data <= 32'hae953a26;
    11'b01011001111: data <= 32'hc0993233;
    11'b01011010000: data <= 32'hc12cb5e1;
    11'b01011010001: data <= 32'hbcd3302f;
    11'b01011010010: data <= 32'hb1423a5a;
    11'b01011010011: data <= 32'hb0db32d6;
    11'b01011010100: data <= 32'haa99bb6f;
    11'b01011010101: data <= 32'h398cb85b;
    11'b01011010110: data <= 32'h3c6e3e45;
    11'b01011010111: data <= 32'h386841f4;
    11'b01011011000: data <= 32'haaca3f9f;
    11'b01011011001: data <= 32'h31eab4bd;
    11'b01011011010: data <= 32'h3875bcc6;
    11'b01011011011: data <= 32'h2efcb8e2;
    11'b01011011100: data <= 32'hb63db4ff;
    11'b01011011101: data <= 32'h37b8bbc3;
    11'b01011011110: data <= 32'h4044bd5b;
    11'b01011011111: data <= 32'h4080b8d3;
    11'b01011100000: data <= 32'h3058340b;
    11'b01011100001: data <= 32'hbffa319f;
    11'b01011100010: data <= 32'hbff7b4d0;
    11'b01011100011: data <= 32'hb933b42f;
    11'b01011100100: data <= 32'hb2dfb0f1;
    11'b01011100101: data <= 32'hbbdfba9f;
    11'b01011100110: data <= 32'hbcd8be0b;
    11'b01011100111: data <= 32'hafc8b8a4;
    11'b01011101000: data <= 32'h3b323eaf;
    11'b01011101001: data <= 32'h38cc41b5;
    11'b01011101010: data <= 32'hb4ee3ed8;
    11'b01011101011: data <= 32'hb87aa8d4;
    11'b01011101100: data <= 32'hb4c3b2c2;
    11'b01011101101: data <= 32'hb4c439ca;
    11'b01011101110: data <= 32'hb16a3949;
    11'b01011101111: data <= 32'h3be2b9db;
    11'b01011110000: data <= 32'h40efbe2c;
    11'b01011110001: data <= 32'h40c8b922;
    11'b01011110010: data <= 32'h38153956;
    11'b01011110011: data <= 32'hbc2839f0;
    11'b01011110100: data <= 32'hb986b04c;
    11'b01011110101: data <= 32'h34efb9dc;
    11'b01011110110: data <= 32'had13bbc0;
    11'b01011110111: data <= 32'hbddfbdfb;
    11'b01011111000: data <= 32'hbea3bf7b;
    11'b01011111001: data <= 32'haee6bb93;
    11'b01011111010: data <= 32'h3caf3b57;
    11'b01011111011: data <= 32'h388f3f32;
    11'b01011111100: data <= 32'hbb8c3b8c;
    11'b01011111101: data <= 32'hbe3124cd;
    11'b01011111110: data <= 32'hbc7938a6;
    11'b01011111111: data <= 32'hb9993e63;
    11'b01100000000: data <= 32'hb6233c2f;
    11'b01100000001: data <= 32'h3885ba2b;
    11'b01100000010: data <= 32'h3f36bdcd;
    11'b01100000011: data <= 32'h3fc1a189;
    11'b01100000100: data <= 32'h3a613ea2;
    11'b01100000101: data <= 32'h12333e2f;
    11'b01100000110: data <= 32'h380c30a1;
    11'b01100000111: data <= 32'h3bfeba67;
    11'b01100001000: data <= 32'h20c4bbad;
    11'b01100001001: data <= 32'hbde3bd0c;
    11'b01100001010: data <= 32'hbcf1bf05;
    11'b01100001011: data <= 32'h399abdbc;
    11'b01100001100: data <= 32'h3f4fb404;
    11'b01100001101: data <= 32'h391a3762;
    11'b01100001110: data <= 32'hbd682fd9;
    11'b01100001111: data <= 32'hbfdbabf9;
    11'b01100010000: data <= 32'hbd183a82;
    11'b01100010001: data <= 32'hbaa63e2d;
    11'b01100010010: data <= 32'hbba438a1;
    11'b01100010011: data <= 32'hb8a3bcc6;
    11'b01100010100: data <= 32'h382bbd41;
    11'b01100010101: data <= 32'h3cc0397b;
    11'b01100010110: data <= 32'h3af340dc;
    11'b01100010111: data <= 32'h385c3ff3;
    11'b01100011000: data <= 32'h3b1e35fe;
    11'b01100011001: data <= 32'h3b8ab528;
    11'b01100011010: data <= 32'hb112a2a1;
    11'b01100011011: data <= 32'hbcd4b268;
    11'b01100011100: data <= 32'hb67dbce3;
    11'b01100011101: data <= 32'h3ea9bf0b;
    11'b01100011110: data <= 32'h40d5bc8a;
    11'b01100011111: data <= 32'h3a8fb53c;
    11'b01100100000: data <= 32'hbc8fb1d0;
    11'b01100100001: data <= 32'hbd86adb7;
    11'b01100100010: data <= 32'hb85b384d;
    11'b01100100011: data <= 32'hb8933a2e;
    11'b01100100100: data <= 32'hbe30b5d9;
    11'b01100100101: data <= 32'hbf0bbf10;
    11'b01100100110: data <= 32'hb88fbd5d;
    11'b01100100111: data <= 32'h394b3aae;
    11'b01100101000: data <= 32'h3a50409f;
    11'b01100101001: data <= 32'h36673e98;
    11'b01100101010: data <= 32'h359a35be;
    11'b01100101011: data <= 32'h32cc36f1;
    11'b01100101100: data <= 32'hb87f3d57;
    11'b01100101101: data <= 32'hbc133c30;
    11'b01100101110: data <= 32'h2e87b925;
    11'b01100101111: data <= 32'h3ffdbf36;
    11'b01100110000: data <= 32'h40e3bd17;
    11'b01100110001: data <= 32'h3bb6b08c;
    11'b01100110010: data <= 32'hb6333336;
    11'b01100110011: data <= 32'hac662c5c;
    11'b01100110100: data <= 32'h39733033;
    11'b01100110101: data <= 32'had579e84;
    11'b01100110110: data <= 32'hbf5ebc18;
    11'b01100110111: data <= 32'hc097c019;
    11'b01100111000: data <= 32'hba74be1b;
    11'b01100111001: data <= 32'h39e2341b;
    11'b01100111010: data <= 32'h39db3cfd;
    11'b01100111011: data <= 32'hb0bf3902;
    11'b01100111100: data <= 32'hb8852bc1;
    11'b01100111101: data <= 32'hb8b43c13;
    11'b01100111110: data <= 32'hbb5e4092;
    11'b01100111111: data <= 32'hbc6b3ecf;
    11'b01101000000: data <= 32'hb198b71c;
    11'b01101000001: data <= 32'h3d50bea0;
    11'b01101000010: data <= 32'h3f0ab9ea;
    11'b01101000011: data <= 32'h3b4039ed;
    11'b01101000100: data <= 32'h36ff3bed;
    11'b01101000101: data <= 32'h3ccb3547;
    11'b01101000110: data <= 32'h3ea4a2ab;
    11'b01101000111: data <= 32'h3481aec4;
    11'b01101001000: data <= 32'hbf0cba59;
    11'b01101001001: data <= 32'hbfe5beed;
    11'b01101001010: data <= 32'hb078bec4;
    11'b01101001011: data <= 32'h3d4fb994;
    11'b01101001100: data <= 32'h3a60b0fe;
    11'b01101001101: data <= 32'hb8b5b7f2;
    11'b01101001110: data <= 32'hbc36b54e;
    11'b01101001111: data <= 32'hba033c8e;
    11'b01101010000: data <= 32'hbb2140ad;
    11'b01101010001: data <= 32'hbd903da2;
    11'b01101010010: data <= 32'hbc74ba2e;
    11'b01101010011: data <= 32'ha1adbe13;
    11'b01101010100: data <= 32'h399baa1e;
    11'b01101010101: data <= 32'h391c3e33;
    11'b01101010110: data <= 32'h3abd3dc6;
    11'b01101010111: data <= 32'h3ec43705;
    11'b01101011000: data <= 32'h3f40332c;
    11'b01101011001: data <= 32'h33e13934;
    11'b01101011010: data <= 32'hbdf53512;
    11'b01101011011: data <= 32'hbcb4bb30;
    11'b01101011100: data <= 32'h3aa6bea8;
    11'b01101011101: data <= 32'h3fb5bdad;
    11'b01101011110: data <= 32'h3b2abc39;
    11'b01101011111: data <= 32'hb88fbc2f;
    11'b01101100000: data <= 32'hb91fb847;
    11'b01101100001: data <= 32'h22e33ab8;
    11'b01101100010: data <= 32'hb5983e7c;
    11'b01101100011: data <= 32'hbe8337de;
    11'b01101100100: data <= 32'hc03cbd65;
    11'b01101100101: data <= 32'hbcdabdfa;
    11'b01101100110: data <= 32'haea33404;
    11'b01101100111: data <= 32'h35603e51;
    11'b01101101000: data <= 32'h39383c54;
    11'b01101101001: data <= 32'h3ce7316e;
    11'b01101101010: data <= 32'h3c96391c;
    11'b01101101011: data <= 32'hb0b73f42;
    11'b01101101100: data <= 32'hbd183eb1;
    11'b01101101101: data <= 32'hb87ca35b;
    11'b01101101110: data <= 32'h3d29bdc1;
    11'b01101101111: data <= 32'h3fccbdf3;
    11'b01101110000: data <= 32'h3a92bbb3;
    11'b01101110001: data <= 32'hb054b9f8;
    11'b01101110010: data <= 32'h37d5b69d;
    11'b01101110011: data <= 32'h3d6136bd;
    11'b01101110100: data <= 32'h375b3a2d;
    11'b01101110101: data <= 32'hbe7bb458;
    11'b01101110110: data <= 32'hc11dbe91;
    11'b01101110111: data <= 32'hbe3abe01;
    11'b01101111000: data <= 32'hb1dba926;
    11'b01101111001: data <= 32'h3298398b;
    11'b01101111010: data <= 32'h2e1da8ca;
    11'b01101111011: data <= 32'h346ab744;
    11'b01101111100: data <= 32'h34403b31;
    11'b01101111101: data <= 32'hb83c414e;
    11'b01101111110: data <= 32'hbce340e5;
    11'b01101111111: data <= 32'hb8ad3621;
    11'b01110000000: data <= 32'h3a5abcb3;
    11'b01110000001: data <= 32'h3cb8bb83;
    11'b01110000010: data <= 32'h371dacd6;
    11'b01110000011: data <= 32'h35a52c57;
    11'b01110000100: data <= 32'h3e86afe7;
    11'b01110000101: data <= 32'h40e931b4;
    11'b01110000110: data <= 32'h3c44374d;
    11'b01110000111: data <= 32'hbd82b2b5;
    11'b01110001000: data <= 32'hc06abd0d;
    11'b01110001001: data <= 32'hbb4fbd77;
    11'b01110001010: data <= 32'h36b8b940;
    11'b01110001011: data <= 32'h34aab89b;
    11'b01110001100: data <= 32'hb69abd37;
    11'b01110001101: data <= 32'hb644bc81;
    11'b01110001110: data <= 32'hab7f3a80;
    11'b01110001111: data <= 32'hb76b4153;
    11'b01110010000: data <= 32'hbcf44069;
    11'b01110010001: data <= 32'hbcc52d8b;
    11'b01110010010: data <= 32'hb677bc28;
    11'b01110010011: data <= 32'ha6eab262;
    11'b01110010100: data <= 32'hb04b3b05;
    11'b01110010101: data <= 32'h3819395d;
    11'b01110010110: data <= 32'h4023a63d;
    11'b01110010111: data <= 32'h416031df;
    11'b01110011000: data <= 32'h3c713b33;
    11'b01110011001: data <= 32'hbc4f3a03;
    11'b01110011010: data <= 32'hbd7eb491;
    11'b01110011011: data <= 32'h3166bc08;
    11'b01110011100: data <= 32'h3c9cbc67;
    11'b01110011101: data <= 32'h3669bda4;
    11'b01110011110: data <= 32'hb8b0bfdb;
    11'b01110011111: data <= 32'hb448bdd9;
    11'b01110100000: data <= 32'h38683738;
    11'b01110100001: data <= 32'h32943fa8;
    11'b01110100010: data <= 32'hbc903cd6;
    11'b01110100011: data <= 32'hbf97b8d1;
    11'b01110100100: data <= 32'hbe20bc27;
    11'b01110100101: data <= 32'hbbc13419;
    11'b01110100110: data <= 32'hb8fd3cae;
    11'b01110100111: data <= 32'h330e3785;
    11'b01110101000: data <= 32'h3e4db661;
    11'b01110101001: data <= 32'h3fe83463;
    11'b01110101010: data <= 32'h39113f03;
    11'b01110101011: data <= 32'hbb1e400c;
    11'b01110101100: data <= 32'hb90c3a0f;
    11'b01110101101: data <= 32'h3af1b85e;
    11'b01110101110: data <= 32'h3d5dbc18;
    11'b01110101111: data <= 32'h33f1bd27;
    11'b01110110000: data <= 32'hb746bea0;
    11'b01110110001: data <= 32'h3865bd2f;
    11'b01110110010: data <= 32'h3f272aef;
    11'b01110110011: data <= 32'h3cbe3bb5;
    11'b01110110100: data <= 32'hbad83359;
    11'b01110110101: data <= 32'hc04dbc43;
    11'b01110110110: data <= 32'hbf5fbbf6;
    11'b01110110111: data <= 32'hbc5533bc;
    11'b01110111000: data <= 32'hba1338be;
    11'b01110111001: data <= 32'hb551b85e;
    11'b01110111010: data <= 32'h3859bcc9;
    11'b01110111011: data <= 32'h3b413355;
    11'b01110111100: data <= 32'h2d2f40be;
    11'b01110111101: data <= 32'hba894187;
    11'b01110111110: data <= 32'hb6843cec;
    11'b01110111111: data <= 32'h3964b30b;
    11'b01111000000: data <= 32'h3983b737;
    11'b01111000001: data <= 32'hb4b9b55e;
    11'b01111000010: data <= 32'hb498b97d;
    11'b01111000011: data <= 32'h3dcbbac4;
    11'b01111000100: data <= 32'h41bab1fc;
    11'b01111000101: data <= 32'h3fa036e3;
    11'b01111000110: data <= 32'hb7e59b10;
    11'b01111000111: data <= 32'hbefaba8f;
    11'b01111001000: data <= 32'hbc95b9ae;
    11'b01111001001: data <= 32'hb5c9aa48;
    11'b01111001010: data <= 32'hb849b6a6;
    11'b01111001011: data <= 32'hba99bf1b;
    11'b01111001100: data <= 32'hb4fbc008;
    11'b01111001101: data <= 32'h34c3a78d;
    11'b01111001110: data <= 32'h9e794093;
    11'b01111001111: data <= 32'hb9ab40f4;
    11'b01111010000: data <= 32'hb9923adb;
    11'b01111010001: data <= 32'hb400b205;
    11'b01111010010: data <= 32'hb7a03458;
    11'b01111010011: data <= 32'hbc313a3c;
    11'b01111010100: data <= 32'hb58c31fa;
    11'b01111010101: data <= 32'h3f0cb89c;
    11'b01111010110: data <= 32'h4220b463;
    11'b01111010111: data <= 32'h3fad388c;
    11'b01111011000: data <= 32'hb4123962;
    11'b01111011001: data <= 32'hbb552eaa;
    11'b01111011010: data <= 32'h2cedb13b;
    11'b01111011011: data <= 32'h38fbb38b;
    11'b01111011100: data <= 32'hb3e4bc64;
    11'b01111011101: data <= 32'hbc3ec0d4;
    11'b01111011110: data <= 32'hb790c0bd;
    11'b01111011111: data <= 32'h38e9b616;
    11'b01111100000: data <= 32'h38ba3e20;
    11'b01111100001: data <= 32'hb6bb3d6f;
    11'b01111100010: data <= 32'hbc74ab75;
    11'b01111100011: data <= 32'hbccbb5dc;
    11'b01111100100: data <= 32'hbda43a1e;
    11'b01111100101: data <= 32'hbe6d3d58;
    11'b01111100110: data <= 32'hb976348d;
    11'b01111100111: data <= 32'h3cf4bad7;
    11'b01111101000: data <= 32'h407fb5cc;
    11'b01111101001: data <= 32'h3cfc3c7a;
    11'b01111101010: data <= 32'hb38b3ef9;
    11'b01111101011: data <= 32'hb0e73c94;
    11'b01111101100: data <= 32'h3c1436a3;
    11'b01111101101: data <= 32'h3c73ab79;
    11'b01111101110: data <= 32'hb476bb63;
    11'b01111101111: data <= 32'hbc59c00f;
    11'b01111110000: data <= 32'h28a8c019;
    11'b01111110001: data <= 32'h3e85b908;
    11'b01111110010: data <= 32'h3e46388d;
    11'b01111110011: data <= 32'h246f30e0;
    11'b01111110100: data <= 32'hbcddba97;
    11'b01111110101: data <= 32'hbdbeb77b;
    11'b01111110110: data <= 32'hbde33b14;
    11'b01111110111: data <= 32'hbe8d3c42;
    11'b01111111000: data <= 32'hbc7bb7e3;
    11'b01111111001: data <= 32'h3256be91;
    11'b01111111010: data <= 32'h3bc6b8ac;
    11'b01111111011: data <= 32'h36533e2b;
    11'b01111111100: data <= 32'hb53f40c5;
    11'b01111111101: data <= 32'h31c73e5c;
    11'b01111111110: data <= 32'h3c84398c;
    11'b01111111111: data <= 32'h39bb3717;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    