
module memory_rom_27(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3990bdb2;
    11'b00000000001: data <= 32'h3570ba6f;
    11'b00000000010: data <= 32'hb7633ab6;
    11'b00000000011: data <= 32'hbe0d3c6d;
    11'b00000000100: data <= 32'hbe66b945;
    11'b00000000101: data <= 32'hb8c2c091;
    11'b00000000110: data <= 32'h246fbf4c;
    11'b00000000111: data <= 32'hb862ae46;
    11'b00000001000: data <= 32'hbbfa3b57;
    11'b00000001001: data <= 32'hacb13b79;
    11'b00000001010: data <= 32'h3c763c51;
    11'b00000001011: data <= 32'h38823e31;
    11'b00000001100: data <= 32'hbd7f3d66;
    11'b00000001101: data <= 32'hc0413565;
    11'b00000001110: data <= 32'hb7fab477;
    11'b00000001111: data <= 32'h3e942b0f;
    11'b00000010000: data <= 32'h403133fc;
    11'b00000010001: data <= 32'h3ccbb79c;
    11'b00000010010: data <= 32'h39d5bbdc;
    11'b00000010011: data <= 32'h3bf6222a;
    11'b00000010100: data <= 32'h3a353dd5;
    11'b00000010101: data <= 32'hb4303c59;
    11'b00000010110: data <= 32'hbb91bcb1;
    11'b00000010111: data <= 32'hb91ec190;
    11'b00000011000: data <= 32'hb403c015;
    11'b00000011001: data <= 32'hb7c3b4fd;
    11'b00000011010: data <= 32'hb85133da;
    11'b00000011011: data <= 32'h34c8b403;
    11'b00000011100: data <= 32'h3b38ae89;
    11'b00000011101: data <= 32'hb2d03c05;
    11'b00000011110: data <= 32'hc06c3e6d;
    11'b00000011111: data <= 32'hc1383b92;
    11'b00000100000: data <= 32'hba102d03;
    11'b00000100001: data <= 32'h3c91a521;
    11'b00000100010: data <= 32'h3ca62fdf;
    11'b00000100011: data <= 32'h33d3b08d;
    11'b00000100100: data <= 32'h3675aeba;
    11'b00000100101: data <= 32'h3e213bf3;
    11'b00000100110: data <= 32'h3f024019;
    11'b00000100111: data <= 32'h37b93d0e;
    11'b00000101000: data <= 32'hb9c2bbdf;
    11'b00000101001: data <= 32'hb8fdc085;
    11'b00000101010: data <= 32'h2ccfbdbd;
    11'b00000101011: data <= 32'h3516b37d;
    11'b00000101100: data <= 32'h360bb83e;
    11'b00000101101: data <= 32'h3a8bbe14;
    11'b00000101110: data <= 32'h3b1ebc8d;
    11'b00000101111: data <= 32'hb66338e7;
    11'b00000110000: data <= 32'hc0553e75;
    11'b00000110001: data <= 32'hc0cc3a60;
    11'b00000110010: data <= 32'hbb2db7d7;
    11'b00000110011: data <= 32'h3419b9be;
    11'b00000110100: data <= 32'hb34fb224;
    11'b00000110101: data <= 32'hbb642fe3;
    11'b00000110110: data <= 32'ha1bb3705;
    11'b00000110111: data <= 32'h3ee33d79;
    11'b00000111000: data <= 32'h3fc54059;
    11'b00000111001: data <= 32'h34763e23;
    11'b00000111010: data <= 32'hbc7cb0bd;
    11'b00000111011: data <= 32'hb9a2bbbb;
    11'b00000111100: data <= 32'h389cb550;
    11'b00000111101: data <= 32'h3c8e2c8e;
    11'b00000111110: data <= 32'h3c24bbf1;
    11'b00000111111: data <= 32'h3c84c047;
    11'b00001000000: data <= 32'h3c9cbd79;
    11'b00001000001: data <= 32'h337f39b6;
    11'b00001000010: data <= 32'hbc9e3e22;
    11'b00001000011: data <= 32'hbe2b31b4;
    11'b00001000100: data <= 32'hba70bdc9;
    11'b00001000101: data <= 32'hb7d5bdf9;
    11'b00001000110: data <= 32'hbcffb816;
    11'b00001000111: data <= 32'hbe41279b;
    11'b00001001000: data <= 32'hb0fa3058;
    11'b00001001001: data <= 32'h3e6f3a01;
    11'b00001001010: data <= 32'h3d963ea5;
    11'b00001001011: data <= 32'hb8fb3eca;
    11'b00001001100: data <= 32'hbf6d3a9d;
    11'b00001001101: data <= 32'hbb25353e;
    11'b00001001110: data <= 32'h3a3138a8;
    11'b00001001111: data <= 32'h3cfe3587;
    11'b00001010000: data <= 32'h3ab6bbe1;
    11'b00001010001: data <= 32'h3b8bbf6d;
    11'b00001010010: data <= 32'h3e10b9c7;
    11'b00001010011: data <= 32'h3d4f3d14;
    11'b00001010100: data <= 32'h33953e20;
    11'b00001010101: data <= 32'hb868b554;
    11'b00001010110: data <= 32'hb87ebfe4;
    11'b00001010111: data <= 32'hb9abbeb6;
    11'b00001011000: data <= 32'hbd6bb864;
    11'b00001011001: data <= 32'hbd3eb63a;
    11'b00001011010: data <= 32'h301fbb4d;
    11'b00001011011: data <= 32'h3db1b87d;
    11'b00001011100: data <= 32'h39473a38;
    11'b00001011101: data <= 32'hbdd63e90;
    11'b00001011110: data <= 32'hc0a33d74;
    11'b00001011111: data <= 32'hbc163ae3;
    11'b00001100000: data <= 32'h37b139fd;
    11'b00001100001: data <= 32'h37003573;
    11'b00001100010: data <= 32'hb376b970;
    11'b00001100011: data <= 32'h3497bc34;
    11'b00001100100: data <= 32'h3ee93368;
    11'b00001100101: data <= 32'h406c3f64;
    11'b00001100110: data <= 32'h3ca63e7b;
    11'b00001100111: data <= 32'ha9d1b4ec;
    11'b00001101000: data <= 32'hb61ebe3c;
    11'b00001101001: data <= 32'hb66ebbc1;
    11'b00001101010: data <= 32'hb937b131;
    11'b00001101011: data <= 32'hb73cbabc;
    11'b00001101100: data <= 32'h3917c028;
    11'b00001101101: data <= 32'h3d72bf1f;
    11'b00001101110: data <= 32'h35ac2cb6;
    11'b00001101111: data <= 32'hbe063dc5;
    11'b00001110000: data <= 32'hc00d3cde;
    11'b00001110001: data <= 32'hbb1136ad;
    11'b00001110010: data <= 32'hae3330ba;
    11'b00001110011: data <= 32'hbac629e0;
    11'b00001110100: data <= 32'hbe58b65e;
    11'b00001110101: data <= 32'hb76bb6e4;
    11'b00001110110: data <= 32'h3eb23977;
    11'b00001110111: data <= 32'h40c63fa9;
    11'b00001111000: data <= 32'h3c6a3e9c;
    11'b00001111001: data <= 32'hb4ef33c6;
    11'b00001111010: data <= 32'hb6beb5ef;
    11'b00001111011: data <= 32'h2e103508;
    11'b00001111100: data <= 32'h328d37e8;
    11'b00001111101: data <= 32'h343ebc20;
    11'b00001111110: data <= 32'h3b54c155;
    11'b00001111111: data <= 32'h3dbac05a;
    11'b00010000000: data <= 32'h39dba045;
    11'b00010000001: data <= 32'hb8cf3d27;
    11'b00010000010: data <= 32'hbbfc38e5;
    11'b00010000011: data <= 32'hb6f7b84f;
    11'b00010000100: data <= 32'hb865b954;
    11'b00010000101: data <= 32'hbf4cb42d;
    11'b00010000110: data <= 32'hc0d2b585;
    11'b00010000111: data <= 32'hbaafb81a;
    11'b00010001000: data <= 32'h3dce3181;
    11'b00010001001: data <= 32'h3f6b3d01;
    11'b00010001010: data <= 32'h338f3ddf;
    11'b00010001011: data <= 32'hbc373b50;
    11'b00010001100: data <= 32'hb8de3af9;
    11'b00010001101: data <= 32'h36573dba;
    11'b00010001110: data <= 32'h37fa3c28;
    11'b00010001111: data <= 32'h318fbb01;
    11'b00010010000: data <= 32'h38d7c0ca;
    11'b00010010001: data <= 32'h3de2be61;
    11'b00010010010: data <= 32'h3e163831;
    11'b00010010011: data <= 32'h39da3d21;
    11'b00010010100: data <= 32'h32b927ef;
    11'b00010010101: data <= 32'h2f97bcd9;
    11'b00010010110: data <= 32'hb8a9bb9d;
    11'b00010010111: data <= 32'hbfbfb294;
    11'b00010011000: data <= 32'hc082b798;
    11'b00010011001: data <= 32'hb8ebbd12;
    11'b00010011010: data <= 32'h3d01bc4b;
    11'b00010011011: data <= 32'h3c4c30b6;
    11'b00010011100: data <= 32'hb9b63c48;
    11'b00010011101: data <= 32'hbe713ceb;
    11'b00010011110: data <= 32'hb9633da0;
    11'b00010011111: data <= 32'h35a33eee;
    11'b00010100000: data <= 32'ha8c93c95;
    11'b00010100001: data <= 32'hba98b849;
    11'b00010100010: data <= 32'hb43abe41;
    11'b00010100011: data <= 32'h3d4eb87b;
    11'b00010100100: data <= 32'h40503cbf;
    11'b00010100101: data <= 32'h3e9e3d56;
    11'b00010100110: data <= 32'h3b13b0e3;
    11'b00010100111: data <= 32'h3762bc35;
    11'b00010101000: data <= 32'hb2cfb531;
    11'b00010101001: data <= 32'hbce3360d;
    11'b00010101010: data <= 32'hbd67b890;
    11'b00010101011: data <= 32'ha8d6c056;
    11'b00010101100: data <= 32'h3cb1c091;
    11'b00010101101: data <= 32'h38c7ba0d;
    11'b00010101110: data <= 32'hbbf0393f;
    11'b00010101111: data <= 32'hbda13be2;
    11'b00010110000: data <= 32'hb5c83bb3;
    11'b00010110001: data <= 32'h2fa53c7f;
    11'b00010110010: data <= 32'hbc323a77;
    11'b00010110011: data <= 32'hc054b3f2;
    11'b00010110100: data <= 32'hbcf3ba75;
    11'b00010110101: data <= 32'h3c092e80;
    11'b00010110110: data <= 32'h40653d6d;
    11'b00010110111: data <= 32'h3e693ce4;
    11'b00010111000: data <= 32'h39442cb5;
    11'b00010111001: data <= 32'h36b0b05e;
    11'b00010111010: data <= 32'h34a13b89;
    11'b00010111011: data <= 32'hb42c3d17;
    11'b00010111100: data <= 32'hb728b756;
    11'b00010111101: data <= 32'h35a5c12e;
    11'b00010111110: data <= 32'h3c88c162;
    11'b00010111111: data <= 32'h396cbb5c;
    11'b00011000000: data <= 32'hb5ba3754;
    11'b00011000001: data <= 32'hb68235ce;
    11'b00011000010: data <= 32'h3544aca1;
    11'b00011000011: data <= 32'h9ddd30f1;
    11'b00011000100: data <= 32'hbf583631;
    11'b00011000101: data <= 32'hc204afab;
    11'b00011000110: data <= 32'hbef1b8fd;
    11'b00011000111: data <= 32'h3985b096;
    11'b00011001000: data <= 32'h3e8339de;
    11'b00011001001: data <= 32'h39693a6c;
    11'b00011001010: data <= 32'hb2b3366f;
    11'b00011001011: data <= 32'h2ffd3b2d;
    11'b00011001100: data <= 32'h391d402c;
    11'b00011001101: data <= 32'h343f3ff2;
    11'b00011001110: data <= 32'hb478b0ef;
    11'b00011001111: data <= 32'h2ea9c083;
    11'b00011010000: data <= 32'h3ba6c024;
    11'b00011010001: data <= 32'h3c7cb4db;
    11'b00011010010: data <= 32'h3a023850;
    11'b00011010011: data <= 32'h3aa9b3fb;
    11'b00011010100: data <= 32'h3c5cbb92;
    11'b00011010101: data <= 32'h311eb616;
    11'b00011010110: data <= 32'hbf7135be;
    11'b00011010111: data <= 32'hc1aaabdd;
    11'b00011011000: data <= 32'hbde6bc28;
    11'b00011011001: data <= 32'h3860bc9c;
    11'b00011011010: data <= 32'h3a94b664;
    11'b00011011011: data <= 32'hb727316c;
    11'b00011011100: data <= 32'hbc013794;
    11'b00011011101: data <= 32'ha95b3d49;
    11'b00011011110: data <= 32'h3a0040c7;
    11'b00011011111: data <= 32'h2aa34034;
    11'b00011100000: data <= 32'hbc203152;
    11'b00011100001: data <= 32'hba45bd98;
    11'b00011100010: data <= 32'h387bbb1a;
    11'b00011100011: data <= 32'h3de7389f;
    11'b00011100100: data <= 32'h3e2a39a3;
    11'b00011100101: data <= 32'h3e20b875;
    11'b00011100110: data <= 32'h3dfebc5a;
    11'b00011100111: data <= 32'h38749d6c;
    11'b00011101000: data <= 32'hbc743b8d;
    11'b00011101001: data <= 32'hbf382e11;
    11'b00011101010: data <= 32'hb9a0be8a;
    11'b00011101011: data <= 32'h38b2c06c;
    11'b00011101100: data <= 32'h33f0bd62;
    11'b00011101101: data <= 32'hbc07b5d8;
    11'b00011101110: data <= 32'hbc3a30d0;
    11'b00011101111: data <= 32'h33fb3aab;
    11'b00011110000: data <= 32'h3a123ec0;
    11'b00011110001: data <= 32'hb9223e6a;
    11'b00011110010: data <= 32'hc0683575;
    11'b00011110011: data <= 32'hbf40b885;
    11'b00011110100: data <= 32'h2cbd28b3;
    11'b00011110101: data <= 32'h3d8b3c0a;
    11'b00011110110: data <= 32'h3db9391c;
    11'b00011110111: data <= 32'h3cf9b86e;
    11'b00011111000: data <= 32'h3d5bb7ef;
    11'b00011111001: data <= 32'h3bb73c50;
    11'b00011111010: data <= 32'hadd83f97;
    11'b00011111011: data <= 32'hb9473698;
    11'b00011111100: data <= 32'ha9d1bf85;
    11'b00011111101: data <= 32'h38f5c117;
    11'b00011111110: data <= 32'h3019bdeb;
    11'b00011111111: data <= 32'hb992b801;
    11'b00100000000: data <= 32'hb40fb68a;
    11'b00100000001: data <= 32'h3bfbb40f;
    11'b00100000010: data <= 32'h3aeb37fb;
    11'b00100000011: data <= 32'hbcdb3b5c;
    11'b00100000100: data <= 32'hc1eb35fc;
    11'b00100000101: data <= 32'hc09fb2a0;
    11'b00100000110: data <= 32'hb3ac2f33;
    11'b00100000111: data <= 32'h3ab638d4;
    11'b00100001000: data <= 32'h37463184;
    11'b00100001001: data <= 32'h31eeb78a;
    11'b00100001010: data <= 32'h3a6234b2;
    11'b00100001011: data <= 32'h3cd14040;
    11'b00100001100: data <= 32'h38ab4149;
    11'b00100001101: data <= 32'hb1a43a25;
    11'b00100001110: data <= 32'hab42be18;
    11'b00100001111: data <= 32'h36afbf7e;
    11'b00100010000: data <= 32'h3526b9a2;
    11'b00100010001: data <= 32'h30a0b260;
    11'b00100010010: data <= 32'h3b05bb43;
    11'b00100010011: data <= 32'h3f44bd04;
    11'b00100010100: data <= 32'h3c8bb57b;
    11'b00100010101: data <= 32'hbcb33913;
    11'b00100010110: data <= 32'hc17636da;
    11'b00100010111: data <= 32'hbfb5b617;
    11'b00100011000: data <= 32'hb269b8e0;
    11'b00100011001: data <= 32'h305ab67c;
    11'b00100011010: data <= 32'hba3cb84c;
    11'b00100011011: data <= 32'hbb37b86c;
    11'b00100011100: data <= 32'h35bf38e9;
    11'b00100011101: data <= 32'h3d1f40bf;
    11'b00100011110: data <= 32'h38c8415a;
    11'b00100011111: data <= 32'hb9053ba0;
    11'b00100100000: data <= 32'hba66ba00;
    11'b00100100001: data <= 32'habc0b8b7;
    11'b00100100010: data <= 32'h37c5374f;
    11'b00100100011: data <= 32'h3a5833d4;
    11'b00100100100: data <= 32'h3e18bc9f;
    11'b00100100101: data <= 32'h405fbe6d;
    11'b00100100110: data <= 32'h3dceb478;
    11'b00100100111: data <= 32'hb7c43c32;
    11'b00100101000: data <= 32'hbe743947;
    11'b00100101001: data <= 32'hbb2bba13;
    11'b00100101010: data <= 32'h2f67bdf8;
    11'b00100101011: data <= 32'hb5c1bd30;
    11'b00100101100: data <= 32'hbe23bc4d;
    11'b00100101101: data <= 32'hbd1bbad2;
    11'b00100101110: data <= 32'h373f30de;
    11'b00100101111: data <= 32'h3d633e5f;
    11'b00100110000: data <= 32'h304c3fca;
    11'b00100110001: data <= 32'hbe603aec;
    11'b00100110010: data <= 32'hbf119df0;
    11'b00100110011: data <= 32'hb8b23821;
    11'b00100110100: data <= 32'h35c53cde;
    11'b00100110101: data <= 32'h39663676;
    11'b00100110110: data <= 32'h3cacbcc0;
    11'b00100110111: data <= 32'h3f56bcfe;
    11'b00100111000: data <= 32'h3e7e3899;
    11'b00100111001: data <= 32'h37243fb8;
    11'b00100111010: data <= 32'hb4ca3c2c;
    11'b00100111011: data <= 32'h2dfdbb57;
    11'b00100111100: data <= 32'h3663bf23;
    11'b00100111101: data <= 32'hb7d7bd81;
    11'b00100111110: data <= 32'hbdd5bc43;
    11'b00100111111: data <= 32'hb9cfbcdd;
    11'b00101000000: data <= 32'h3c71bace;
    11'b00101000001: data <= 32'h3e233400;
    11'b00101000010: data <= 32'hb4f63b78;
    11'b00101000011: data <= 32'hc08d3901;
    11'b00101000100: data <= 32'hc0713566;
    11'b00101000101: data <= 32'hba703a9a;
    11'b00101000110: data <= 32'ha92d3c59;
    11'b00101000111: data <= 32'hb3722a94;
    11'b00101001000: data <= 32'ha766bcc3;
    11'b00101001001: data <= 32'h3bd1b8f4;
    11'b00101001010: data <= 32'h3e503e13;
    11'b00101001011: data <= 32'h3c554148;
    11'b00101001100: data <= 32'h369f3d67;
    11'b00101001101: data <= 32'h362ab93c;
    11'b00101001110: data <= 32'h357dbca2;
    11'b00101001111: data <= 32'hb608b7a5;
    11'b00101010000: data <= 32'hba6cb793;
    11'b00101010001: data <= 32'h3467bdbd;
    11'b00101010010: data <= 32'h3f9abf31;
    11'b00101010011: data <= 32'h3f34ba86;
    11'b00101010100: data <= 32'hb4ff3525;
    11'b00101010101: data <= 32'hc02537f8;
    11'b00101010110: data <= 32'hbeef335f;
    11'b00101010111: data <= 32'hb81234f3;
    11'b00101011000: data <= 32'hb7b2339a;
    11'b00101011001: data <= 32'hbda0b905;
    11'b00101011010: data <= 32'hbd55bd38;
    11'b00101011011: data <= 32'h323fb4e4;
    11'b00101011100: data <= 32'h3dc13f17;
    11'b00101011101: data <= 32'h3c93412e;
    11'b00101011110: data <= 32'h31e03d4a;
    11'b00101011111: data <= 32'hb14caf50;
    11'b00101100000: data <= 32'haded2c39;
    11'b00101100001: data <= 32'hb4623b22;
    11'b00101100010: data <= 32'hb2973527;
    11'b00101100011: data <= 32'h3b42bdc0;
    11'b00101100100: data <= 32'h406cc059;
    11'b00101100101: data <= 32'h3fcdbbde;
    11'b00101100110: data <= 32'h31be3812;
    11'b00101100111: data <= 32'hbc08394f;
    11'b00101101000: data <= 32'hb80aac9b;
    11'b00101101001: data <= 32'h3108b7b7;
    11'b00101101010: data <= 32'hb9b7b8f3;
    11'b00101101011: data <= 32'hc056bc87;
    11'b00101101100: data <= 32'hbfcabdf8;
    11'b00101101101: data <= 32'h26c1b8e4;
    11'b00101101110: data <= 32'h3da13c28;
    11'b00101101111: data <= 32'h3a143eba;
    11'b00101110000: data <= 32'hb9433b2b;
    11'b00101110001: data <= 32'hbc4935c4;
    11'b00101110010: data <= 32'hb8cf3cab;
    11'b00101110011: data <= 32'hb5663f9a;
    11'b00101110100: data <= 32'hb2cc3a38;
    11'b00101110101: data <= 32'h38bebd5a;
    11'b00101110110: data <= 32'h3ed3bf90;
    11'b00101110111: data <= 32'h3f3db483;
    11'b00101111000: data <= 32'h3ac23d33;
    11'b00101111001: data <= 32'h34b13c24;
    11'b00101111010: data <= 32'h39ebb3f1;
    11'b00101111011: data <= 32'h3a24babb;
    11'b00101111100: data <= 32'hb96db9d8;
    11'b00101111101: data <= 32'hc051bc00;
    11'b00101111110: data <= 32'hbe4dbe52;
    11'b00101111111: data <= 32'h387dbd73;
    11'b00110000000: data <= 32'h3e50b48f;
    11'b00110000001: data <= 32'h354a3698;
    11'b00110000010: data <= 32'hbd7634e2;
    11'b00110000011: data <= 32'hbe33380b;
    11'b00110000100: data <= 32'hb9d73e22;
    11'b00110000101: data <= 32'hb8153fe6;
    11'b00110000110: data <= 32'hbb2338af;
    11'b00110000111: data <= 32'hb8a5bd3e;
    11'b00110001000: data <= 32'h38cebd33;
    11'b00110001001: data <= 32'h3d9a3934;
    11'b00110001010: data <= 32'h3d08400b;
    11'b00110001011: data <= 32'h3c393d23;
    11'b00110001100: data <= 32'h3d0cb137;
    11'b00110001101: data <= 32'h3b52b697;
    11'b00110001110: data <= 32'hb819307c;
    11'b00110001111: data <= 32'hbe3ab1a7;
    11'b00110010000: data <= 32'hb8f5bdbf;
    11'b00110010001: data <= 32'h3d64c023;
    11'b00110010010: data <= 32'h3f3ebd90;
    11'b00110010011: data <= 32'h3257b744;
    11'b00110010100: data <= 32'hbd4dac93;
    11'b00110010101: data <= 32'hbc5e350d;
    11'b00110010110: data <= 32'hb3553c53;
    11'b00110010111: data <= 32'hb8d63cd2;
    11'b00110011000: data <= 32'hbf47ac78;
    11'b00110011001: data <= 32'hbfacbda3;
    11'b00110011010: data <= 32'hb742bb32;
    11'b00110011011: data <= 32'h3bbe3c24;
    11'b00110011100: data <= 32'h3cce4003;
    11'b00110011101: data <= 32'h3b283c53;
    11'b00110011110: data <= 32'h3aa22b88;
    11'b00110011111: data <= 32'h38443892;
    11'b00110100000: data <= 32'hb66e3e26;
    11'b00110100001: data <= 32'hbb4a3b36;
    11'b00110100010: data <= 32'h2f39bc74;
    11'b00110100011: data <= 32'h3ecbc097;
    11'b00110100100: data <= 32'h3f4bbe85;
    11'b00110100101: data <= 32'h3683b6c8;
    11'b00110100110: data <= 32'hb7d68835;
    11'b00110100111: data <= 32'h31121684;
    11'b00110101000: data <= 32'h39c6345f;
    11'b00110101001: data <= 32'hb7d5347d;
    11'b00110101010: data <= 32'hc0cfb8ef;
    11'b00110101011: data <= 32'hc135bdfc;
    11'b00110101100: data <= 32'hba89bbb3;
    11'b00110101101: data <= 32'h3a5f3822;
    11'b00110101110: data <= 32'h3a503c56;
    11'b00110101111: data <= 32'h2be73610;
    11'b00110110000: data <= 32'haf0c3197;
    11'b00110110001: data <= 32'ha3513dea;
    11'b00110110010: data <= 32'hb665413d;
    11'b00110110011: data <= 32'hb9bf3e59;
    11'b00110110100: data <= 32'h9a61ba98;
    11'b00110110101: data <= 32'h3cc7bfd7;
    11'b00110110110: data <= 32'h3db2bba7;
    11'b00110110111: data <= 32'h39b835cb;
    11'b00110111000: data <= 32'h38db3656;
    11'b00110111001: data <= 32'h3decb2d6;
    11'b00110111010: data <= 32'h3e61b3c2;
    11'b00110111011: data <= 32'hb2fba18d;
    11'b00110111100: data <= 32'hc0a3b807;
    11'b00110111101: data <= 32'hc08dbd6d;
    11'b00110111110: data <= 32'hb53cbd79;
    11'b00110111111: data <= 32'h3bbbb8c7;
    11'b00111000000: data <= 32'h355fb434;
    11'b00111000001: data <= 32'hba1cb801;
    11'b00111000010: data <= 32'hb9f8297f;
    11'b00111000011: data <= 32'hb1b93efb;
    11'b00111000100: data <= 32'hb6224182;
    11'b00111000101: data <= 32'hbc4f3df0;
    11'b00111000110: data <= 32'hbbb7ba19;
    11'b00111000111: data <= 32'h24a2bd64;
    11'b00111001000: data <= 32'h39af2bed;
    11'b00111001001: data <= 32'h3a893cdf;
    11'b00111001010: data <= 32'h3cfe398b;
    11'b00111001011: data <= 32'h4028b474;
    11'b00111001100: data <= 32'h3f83ae84;
    11'b00111001101: data <= 32'h26013932;
    11'b00111001110: data <= 32'hbec43607;
    11'b00111001111: data <= 32'hbd0cbb44;
    11'b00111010000: data <= 32'h3888bef6;
    11'b00111010001: data <= 32'h3d02be40;
    11'b00111010010: data <= 32'h2daabce4;
    11'b00111010011: data <= 32'hbbd4bc41;
    11'b00111010100: data <= 32'hb7e4b450;
    11'b00111010101: data <= 32'h35c53d08;
    11'b00111010110: data <= 32'hb1f03fd1;
    11'b00111010111: data <= 32'hbea53a07;
    11'b00111011000: data <= 32'hc04bbb4b;
    11'b00111011001: data <= 32'hbc91bae5;
    11'b00111011010: data <= 32'h29e2395d;
    11'b00111011011: data <= 32'h38b33d9c;
    11'b00111011100: data <= 32'h3c273792;
    11'b00111011101: data <= 32'h3e96b533;
    11'b00111011110: data <= 32'h3dd83853;
    11'b00111011111: data <= 32'h2e223f86;
    11'b00111100000: data <= 32'hbbdd3e44;
    11'b00111100001: data <= 32'hb562b50b;
    11'b00111100010: data <= 32'h3c71befe;
    11'b00111100011: data <= 32'h3d15bef3;
    11'b00111100100: data <= 32'h2b82bce3;
    11'b00111100101: data <= 32'hb792bc06;
    11'b00111100110: data <= 32'h38acb890;
    11'b00111100111: data <= 32'h3db0366e;
    11'b00111101000: data <= 32'h332a3aef;
    11'b00111101001: data <= 32'hbff62578;
    11'b00111101010: data <= 32'hc181bc1d;
    11'b00111101011: data <= 32'hbe42b9c0;
    11'b00111101100: data <= 32'hb23a3776;
    11'b00111101101: data <= 32'h30e43948;
    11'b00111101110: data <= 32'h3146b550;
    11'b00111101111: data <= 32'h389cb820;
    11'b00111110000: data <= 32'h39f63ca7;
    11'b00111110001: data <= 32'h2a5b41be;
    11'b00111110010: data <= 32'hb8f240ad;
    11'b00111110011: data <= 32'hb0f52e4a;
    11'b00111110100: data <= 32'h3a5fbd63;
    11'b00111110101: data <= 32'h3a49bc17;
    11'b00111110110: data <= 32'h2b88b56c;
    11'b00111110111: data <= 32'h3524b77e;
    11'b00111111000: data <= 32'h3f39b9d4;
    11'b00111111001: data <= 32'h40cfb40d;
    11'b00111111010: data <= 32'h396034c4;
    11'b00111111011: data <= 32'hbf2bac37;
    11'b00111111100: data <= 32'hc0c2baa0;
    11'b00111111101: data <= 32'hbc0cba9f;
    11'b00111111110: data <= 32'h2d1bb558;
    11'b00111111111: data <= 32'hb3f4b89e;
    11'b01000000000: data <= 32'hba32bd5e;
    11'b01000000001: data <= 32'hb50abaf7;
    11'b01000000010: data <= 32'h35f33d1c;
    11'b01000000011: data <= 32'h2e2b41ea;
    11'b01000000100: data <= 32'hb99b406b;
    11'b01000000101: data <= 32'hba612e79;
    11'b01000000110: data <= 32'hb41fba29;
    11'b01000000111: data <= 32'hac542dd2;
    11'b01000001000: data <= 32'hae6c39fb;
    11'b01000001001: data <= 32'h3a2e2904;
    11'b01000001010: data <= 32'h40b5ba5b;
    11'b01000001011: data <= 32'h4168b5cb;
    11'b01000001100: data <= 32'h3b40391f;
    11'b01000001101: data <= 32'hbcb33967;
    11'b01000001110: data <= 32'hbd21b3b9;
    11'b01000001111: data <= 32'h2d80bb4b;
    11'b01000010000: data <= 32'h388fbc50;
    11'b01000010001: data <= 32'hb796bdf2;
    11'b01000010010: data <= 32'hbcd7bfd9;
    11'b01000010011: data <= 32'hb600bcee;
    11'b01000010100: data <= 32'h3a073a27;
    11'b01000010101: data <= 32'h36ae402b;
    11'b01000010110: data <= 32'hbbe03d38;
    11'b01000010111: data <= 32'hbeedb39b;
    11'b01000011000: data <= 32'hbd75b51d;
    11'b01000011001: data <= 32'hbaa13b2b;
    11'b01000011010: data <= 32'hb7003cf4;
    11'b01000011011: data <= 32'h380f9afd;
    11'b01000011100: data <= 32'h3f71bb89;
    11'b01000011101: data <= 32'h404da4de;
    11'b01000011110: data <= 32'h3a843e6a;
    11'b01000011111: data <= 32'hb80f3f37;
    11'b01000100000: data <= 32'hb1cd37a4;
    11'b01000100001: data <= 32'h3b70ba0e;
    11'b01000100010: data <= 32'h3a45bca4;
    11'b01000100011: data <= 32'hb89fbdbe;
    11'b01000100100: data <= 32'hbbf7bf40;
    11'b01000100101: data <= 32'h36bdbda1;
    11'b01000100110: data <= 32'h3ef8aa55;
    11'b01000100111: data <= 32'h3bc63abb;
    11'b01000101000: data <= 32'hbc6c3488;
    11'b01000101001: data <= 32'hc06cb886;
    11'b01000101010: data <= 32'hbefcb02a;
    11'b01000101011: data <= 32'hbc1c3bc2;
    11'b01000101100: data <= 32'hba5d3a4f;
    11'b01000101101: data <= 32'hb578b9c3;
    11'b01000101110: data <= 32'h3939bd23;
    11'b01000101111: data <= 32'h3ca635cf;
    11'b01000110000: data <= 32'h386340e0;
    11'b01000110001: data <= 32'hafd14116;
    11'b01000110010: data <= 32'h343a3b32;
    11'b01000110011: data <= 32'h3b5ab605;
    11'b01000110100: data <= 32'h3689b730;
    11'b01000110101: data <= 32'hb9ceb6f6;
    11'b01000110110: data <= 32'hb76cbc1f;
    11'b01000110111: data <= 32'h3dd9bd64;
    11'b01000111000: data <= 32'h4166b9a1;
    11'b01000111001: data <= 32'h3de5261b;
    11'b01000111010: data <= 32'hbaf9afa8;
    11'b01000111011: data <= 32'hbf42b804;
    11'b01000111100: data <= 32'hbc61aeaa;
    11'b01000111101: data <= 32'hb85d3724;
    11'b01000111110: data <= 32'hbbf9b3df;
    11'b01000111111: data <= 32'hbd11bed5;
    11'b01001000000: data <= 32'hb785beef;
    11'b01001000001: data <= 32'h37713638;
    11'b01001000010: data <= 32'h36dc40f3;
    11'b01001000011: data <= 32'hadd240ac;
    11'b01001000100: data <= 32'hadf939eb;
    11'b01001000101: data <= 32'h2dcd27a6;
    11'b01001000110: data <= 32'hb6b6392f;
    11'b01001000111: data <= 32'hbc0b3aed;
    11'b01001001000: data <= 32'hb0b7b259;
    11'b01001001001: data <= 32'h3fc3bce3;
    11'b01001001010: data <= 32'h41e2bb35;
    11'b01001001011: data <= 32'h3e622d17;
    11'b01001001100: data <= 32'hb62c35f3;
    11'b01001001101: data <= 32'hb9d529d5;
    11'b01001001110: data <= 32'h326aa950;
    11'b01001001111: data <= 32'h342dafd7;
    11'b01001010000: data <= 32'hbc0cbc42;
    11'b01001010001: data <= 32'hbf11c097;
    11'b01001010010: data <= 32'hba83c012;
    11'b01001010011: data <= 32'h3893a844;
    11'b01001010100: data <= 32'h397e3e6c;
    11'b01001010101: data <= 32'hb3123d02;
    11'b01001010110: data <= 32'hba8d2e7b;
    11'b01001010111: data <= 32'hbb38343d;
    11'b01001011000: data <= 32'hbcac3dfd;
    11'b01001011001: data <= 32'hbd603e8c;
    11'b01001011010: data <= 32'hb6012b3c;
    11'b01001011011: data <= 32'h3dc0bd1a;
    11'b01001011100: data <= 32'h4078b9a5;
    11'b01001011101: data <= 32'h3ced3a7b;
    11'b01001011110: data <= 32'h2c913d73;
    11'b01001011111: data <= 32'h36783a1e;
    11'b01001100000: data <= 32'h3d47311c;
    11'b01001100001: data <= 32'h3a57b227;
    11'b01001100010: data <= 32'hbbefbbf5;
    11'b01001100011: data <= 32'hbec0c00b;
    11'b01001100100: data <= 32'hb44ebfe9;
    11'b01001100101: data <= 32'h3d97b942;
    11'b01001100110: data <= 32'h3cf83565;
    11'b01001100111: data <= 32'hb417a8fa;
    11'b01001101000: data <= 32'hbcf4b87a;
    11'b01001101001: data <= 32'hbd0434d2;
    11'b01001101010: data <= 32'hbd1c3ec5;
    11'b01001101011: data <= 32'hbe123dcf;
    11'b01001101100: data <= 32'hbc39b781;
    11'b01001101101: data <= 32'h32c0be72;
    11'b01001101110: data <= 32'h3be5b700;
    11'b01001101111: data <= 32'h38fc3e2c;
    11'b01001110000: data <= 32'h3477401e;
    11'b01001110001: data <= 32'h3ba63c86;
    11'b01001110010: data <= 32'h3e5b3699;
    11'b01001110011: data <= 32'h391d362e;
    11'b01001110100: data <= 32'hbc7825f8;
    11'b01001110101: data <= 32'hbd25bc00;
    11'b01001110110: data <= 32'h3916be52;
    11'b01001110111: data <= 32'h4098bc77;
    11'b01001111000: data <= 32'h3edfb896;
    11'b01001111001: data <= 32'hae02b9e2;
    11'b01001111010: data <= 32'hbb78ba07;
    11'b01001111011: data <= 32'hb8b0347e;
    11'b01001111100: data <= 32'hb8ab3d3b;
    11'b01001111101: data <= 32'hbd9a38ab;
    11'b01001111110: data <= 32'hbf1fbd87;
    11'b01001111111: data <= 32'hbbf1c01d;
    11'b01010000000: data <= 32'ha347b640;
    11'b01010000001: data <= 32'h32c83e87;
    11'b01010000010: data <= 32'h337c3f56;
    11'b01010000011: data <= 32'h39ec3a56;
    11'b01010000100: data <= 32'h3ba63842;
    11'b01010000101: data <= 32'hade23d28;
    11'b01010000110: data <= 32'hbda63d94;
    11'b01010000111: data <= 32'hbbf03077;
    11'b01010001000: data <= 32'h3c83bc87;
    11'b01010001001: data <= 32'h410bbcd2;
    11'b01010001010: data <= 32'h3ecbb942;
    11'b01010001011: data <= 32'h30b9b781;
    11'b01010001100: data <= 32'ha6aab551;
    11'b01010001101: data <= 32'h3a2f35b8;
    11'b01010001110: data <= 32'h38383a63;
    11'b01010001111: data <= 32'hbc4db2d5;
    11'b01010010000: data <= 32'hc049bfd1;
    11'b01010010001: data <= 32'hbde2c084;
    11'b01010010010: data <= 32'hb12ab8ed;
    11'b01010010011: data <= 32'h34e43b54;
    11'b01010010100: data <= 32'h2efc398b;
    11'b01010010101: data <= 32'h2ea2b06e;
    11'b01010010110: data <= 32'h24d036bd;
    11'b01010010111: data <= 32'hba983fee;
    11'b01010011000: data <= 32'hbebc4096;
    11'b01010011001: data <= 32'hbc4b3966;
    11'b01010011010: data <= 32'h3a0bbbd8;
    11'b01010011011: data <= 32'h3f10bbf8;
    11'b01010011100: data <= 32'h3c40a88c;
    11'b01010011101: data <= 32'h343d36e2;
    11'b01010011110: data <= 32'h3b8735cd;
    11'b01010011111: data <= 32'h4008383f;
    11'b01010100000: data <= 32'h3d723910;
    11'b01010100001: data <= 32'hba79b3ed;
    11'b01010100010: data <= 32'hc00cbe96;
    11'b01010100011: data <= 32'hbc30bfd5;
    11'b01010100100: data <= 32'h384abb58;
    11'b01010100101: data <= 32'h3a8db1de;
    11'b01010100110: data <= 32'h2c89b9c3;
    11'b01010100111: data <= 32'hb5d4bc7c;
    11'b01010101000: data <= 32'hb68b319b;
    11'b01010101001: data <= 32'hbb514039;
    11'b01010101010: data <= 32'hbea1407b;
    11'b01010101011: data <= 32'hbdd93503;
    11'b01010101100: data <= 32'hb4e5bcfc;
    11'b01010101101: data <= 32'h3670b9e2;
    11'b01010101110: data <= 32'h2fc739a4;
    11'b01010101111: data <= 32'h31273cb1;
    11'b01010110000: data <= 32'h3d9f39c7;
    11'b01010110001: data <= 32'h40da3908;
    11'b01010110010: data <= 32'h3da43bab;
    11'b01010110011: data <= 32'hbaa438e7;
    11'b01010110100: data <= 32'hbe85b826;
    11'b01010110101: data <= 32'hb157bcea;
    11'b01010110110: data <= 32'h3dd0bc2e;
    11'b01010110111: data <= 32'h3d2ebbe7;
    11'b01010111000: data <= 32'h2fc9be44;
    11'b01010111001: data <= 32'hb44cbe39;
    11'b01010111010: data <= 32'h2f462164;
    11'b01010111011: data <= 32'hb0373ee9;
    11'b01010111100: data <= 32'hbce23db1;
    11'b01010111101: data <= 32'hbf63b8b0;
    11'b01010111110: data <= 32'hbd8ebec6;
    11'b01010111111: data <= 32'hba0fb8eb;
    11'b01011000000: data <= 32'hb8913bab;
    11'b01011000001: data <= 32'hac9a3c51;
    11'b01011000010: data <= 32'h3cb53509;
    11'b01011000011: data <= 32'h3f7b3754;
    11'b01011000100: data <= 32'h39d13e1d;
    11'b01011000101: data <= 32'hbc7b3f6a;
    11'b01011000110: data <= 32'hbd2c3a44;
    11'b01011000111: data <= 32'h3735b776;
    11'b01011001000: data <= 32'h3f2dbb39;
    11'b01011001001: data <= 32'h3ceabc2b;
    11'b01011001010: data <= 32'h2ef1bd9d;
    11'b01011001011: data <= 32'h3537bce6;
    11'b01011001100: data <= 32'h3d5b2c20;
    11'b01011001101: data <= 32'h3c8e3cc8;
    11'b01011001110: data <= 32'hb87b384e;
    11'b01011001111: data <= 32'hbfc3bd09;
    11'b01011010000: data <= 32'hbf48bf7a;
    11'b01011010001: data <= 32'hbc20b901;
    11'b01011010010: data <= 32'hb8ea383d;
    11'b01011010011: data <= 32'hb3ef2c92;
    11'b01011010100: data <= 32'h383fba25;
    11'b01011010101: data <= 32'h3b0b13d9;
    11'b01011010110: data <= 32'hada43fb5;
    11'b01011010111: data <= 32'hbd8c4162;
    11'b01011011000: data <= 32'hbcce3ddf;
    11'b01011011001: data <= 32'h355bb010;
    11'b01011011010: data <= 32'h3caeb8d5;
    11'b01011011011: data <= 32'h3745b6a7;
    11'b01011011100: data <= 32'haf78b7c8;
    11'b01011011101: data <= 32'h3bddb78b;
    11'b01011011110: data <= 32'h410533ef;
    11'b01011011111: data <= 32'h40483b2f;
    11'b01011100000: data <= 32'hab73346f;
    11'b01011100001: data <= 32'hbec2bc57;
    11'b01011100010: data <= 32'hbd8dbdd0;
    11'b01011100011: data <= 32'hb59db8cc;
    11'b01011100100: data <= 32'hace2b416;
    11'b01011100101: data <= 32'hb45fbd0d;
    11'b01011100110: data <= 32'ha843bfbd;
    11'b01011100111: data <= 32'h3420b82e;
    11'b01011101000: data <= 32'hb5063f87;
    11'b01011101001: data <= 32'hbd17413f;
    11'b01011101010: data <= 32'hbd253ca0;
    11'b01011101011: data <= 32'hb6a7b603;
    11'b01011101100: data <= 32'haee7b588;
    11'b01011101101: data <= 32'hb972364a;
    11'b01011101110: data <= 32'hb84336af;
    11'b01011101111: data <= 32'h3cf325a9;
    11'b01011110000: data <= 32'h41cc34a2;
    11'b01011110001: data <= 32'h408d3ba3;
    11'b01011110010: data <= 32'ha3323ab2;
    11'b01011110011: data <= 32'hbd1baa9c;
    11'b01011110100: data <= 32'hb754b83a;
    11'b01011110101: data <= 32'h398eb642;
    11'b01011110110: data <= 32'h3834ba8f;
    11'b01011110111: data <= 32'hb402c02c;
    11'b01011111000: data <= 32'hb15ac0fb;
    11'b01011111001: data <= 32'h37edba6e;
    11'b01011111010: data <= 32'h35cf3dcc;
    11'b01011111011: data <= 32'hb93a3f12;
    11'b01011111100: data <= 32'hbd4c312e;
    11'b01011111101: data <= 32'hbcf1bb74;
    11'b01011111110: data <= 32'hbcf7b2f7;
    11'b01011111111: data <= 32'hbe1f3ab6;
    11'b01100000000: data <= 32'hbb7d38b7;
    11'b01100000001: data <= 32'h3b6db447;
    11'b01100000010: data <= 32'h40a1a95d;
    11'b01100000011: data <= 32'h3e213cba;
    11'b01100000100: data <= 32'hb63c3f33;
    11'b01100000101: data <= 32'hbb883ce1;
    11'b01100000110: data <= 32'h351b36bc;
    11'b01100000111: data <= 32'h3d1fa675;
    11'b01100001000: data <= 32'h38b4ba12;
    11'b01100001001: data <= 32'hb653bf9d;
    11'b01100001010: data <= 32'h2e69c048;
    11'b01100001011: data <= 32'h3dbeb995;
    11'b01100001100: data <= 32'h3e623b60;
    11'b01100001101: data <= 32'h32e239ff;
    11'b01100001110: data <= 32'hbc99b9e3;
    11'b01100001111: data <= 32'hbe10bcfd;
    11'b01100010000: data <= 32'hbe06b014;
    11'b01100010001: data <= 32'hbe6739b6;
    11'b01100010010: data <= 32'hbc6bb03c;
    11'b01100010011: data <= 32'h3472bd35;
    11'b01100010100: data <= 32'h3cddb9b6;
    11'b01100010101: data <= 32'h381d3d1c;
    11'b01100010110: data <= 32'hba6840e9;
    11'b01100010111: data <= 32'hba3b3f9b;
    11'b01100011000: data <= 32'h37b33ab1;
    11'b01100011001: data <= 32'h3b87351b;
    11'b01100011010: data <= 32'hafedaf0d;
    11'b01100011011: data <= 32'hbaa8bb33;
    11'b01100011100: data <= 32'h36f8bcdb;
    11'b01100011101: data <= 32'h40cdb5ef;
    11'b01100011110: data <= 32'h413338a3;
    11'b01100011111: data <= 32'h3ab63397;
    11'b01100100000: data <= 32'hba5dbac0;
    11'b01100100001: data <= 32'hbc26bb4a;
    11'b01100100010: data <= 32'hba132e39;
    11'b01100100011: data <= 32'hbb693422;
    11'b01100100100: data <= 32'hbc00bcf9;
    11'b01100100101: data <= 32'hb4f7c0f3;
    11'b01100100110: data <= 32'h35e8bd98;
    11'b01100100111: data <= 32'h20fa3c4e;
    11'b01100101000: data <= 32'hba52409f;
    11'b01100101001: data <= 32'hb9803e2c;
    11'b01100101010: data <= 32'h2bb937ed;
    11'b01100101011: data <= 32'hae783799;
    11'b01100101100: data <= 32'hbd1039b3;
    11'b01100101101: data <= 32'hbdc43278;
    11'b01100101110: data <= 32'h37c7b72b;
    11'b01100101111: data <= 32'h4161b281;
    11'b01100110000: data <= 32'h416a37d1;
    11'b01100110001: data <= 32'h3ab93797;
    11'b01100110010: data <= 32'hb724abb3;
    11'b01100110011: data <= 32'hade7234f;
    11'b01100110100: data <= 32'h3759382b;
    11'b01100110101: data <= 32'hac42ac05;
    11'b01100110110: data <= 32'hbaacbfc7;
    11'b01100110111: data <= 32'hb87dc20c;
    11'b01100111000: data <= 32'h34c1bec2;
    11'b01100111001: data <= 32'h36c6394b;
    11'b01100111010: data <= 32'hb1ef3dbb;
    11'b01100111011: data <= 32'hb8003662;
    11'b01100111100: data <= 32'hb7c2b4c0;
    11'b01100111101: data <= 32'hbc5f373e;
    11'b01100111110: data <= 32'hc0423cfd;
    11'b01100111111: data <= 32'hbfa23954;
    11'b01101000000: data <= 32'h30a2b765;
    11'b01101000001: data <= 32'h4023b7f0;
    11'b01101000010: data <= 32'h3f5b37eb;
    11'b01101000011: data <= 32'h34213c90;
    11'b01101000100: data <= 32'hb41d3c33;
    11'b01101000101: data <= 32'h3a063bf4;
    11'b01101000110: data <= 32'h3d483c02;
    11'b01101000111: data <= 32'h347c2d2f;
    11'b01101001000: data <= 32'hbb4cbeda;
    11'b01101001001: data <= 32'hb7f9c127;
    11'b01101001010: data <= 32'h3b6fbda9;
    11'b01101001011: data <= 32'h3de7343b;
    11'b01101001100: data <= 32'h39c535c0;
    11'b01101001101: data <= 32'hb14bba0f;
    11'b01101001110: data <= 32'hb911bb38;
    11'b01101001111: data <= 32'hbd2e3732;
    11'b01101010000: data <= 32'hc0463d38;
    11'b01101010001: data <= 32'hbfd4341c;
    11'b01101010010: data <= 32'hb668bd2f;
    11'b01101010011: data <= 32'h3b60bcd1;
    11'b01101010100: data <= 32'h38a23661;
    11'b01101010101: data <= 32'hb71d3e7b;
    11'b01101010110: data <= 32'hb2be3ea0;
    11'b01101010111: data <= 32'h3c4d3d85;
    11'b01101011000: data <= 32'h3d2c3d22;
    11'b01101011001: data <= 32'hb2c23948;
    11'b01101011010: data <= 32'hbd7eb953;
    11'b01101011011: data <= 32'hb5f7bdb8;
    11'b01101011100: data <= 32'h3ebbba6f;
    11'b01101011101: data <= 32'h40c82b1a;
    11'b01101011110: data <= 32'h3d63b4af;
    11'b01101011111: data <= 32'h31ecbcb7;
    11'b01101100000: data <= 32'hb1c8ba78;
    11'b01101100001: data <= 32'hb80b396f;
    11'b01101100010: data <= 32'hbd153c43;
    11'b01101100011: data <= 32'hbe5ab8ee;
    11'b01101100100: data <= 32'hbac7c0bb;
    11'b01101100101: data <= 32'ha9d7bfaa;
    11'b01101100110: data <= 32'hb3a030a4;
    11'b01101100111: data <= 32'hb9983dd4;
    11'b01101101000: data <= 32'hb0783d03;
    11'b01101101001: data <= 32'h3af53b12;
    11'b01101101010: data <= 32'h38163cd5;
    11'b01101101011: data <= 32'hbcef3d61;
    11'b01101101100: data <= 32'hc00e3854;
    11'b01101101101: data <= 32'hb6c6b5b3;
    11'b01101101110: data <= 32'h3fa2b595;
    11'b01101101111: data <= 32'h40e5234d;
    11'b01101110000: data <= 32'h3cedb434;
    11'b01101110001: data <= 32'h3591b963;
    11'b01101110010: data <= 32'h3924a5b4;
    11'b01101110011: data <= 32'h3a713ca2;
    11'b01101110100: data <= 32'haf473b15;
    11'b01101110101: data <= 32'hbc79bcdd;
    11'b01101110110: data <= 32'hbc12c1bb;
    11'b01101110111: data <= 32'hb4ffc043;
    11'b01101111000: data <= 32'hafbcb056;
    11'b01101111001: data <= 32'hb42a3964;
    11'b01101111010: data <= 32'h2e7c266a;
    11'b01101111011: data <= 32'h37eeb207;
    11'b01101111100: data <= 32'hb58b3b0b;
    11'b01101111101: data <= 32'hc0183f1b;
    11'b01101111110: data <= 32'hc0eb3cbe;
    11'b01101111111: data <= 32'hb97bab7d;
    11'b01110000000: data <= 32'h3d69b71b;
    11'b01110000001: data <= 32'h3e04a50c;
    11'b01110000010: data <= 32'h364c32c8;
    11'b01110000011: data <= 32'h33b83454;
    11'b01110000100: data <= 32'h3d7d3b3a;
    11'b01110000101: data <= 32'h3f553e93;
    11'b01110000110: data <= 32'h38743c05;
    11'b01110000111: data <= 32'hbbbbbc12;
    11'b01110001000: data <= 32'hbbc8c0b3;
    11'b01110001001: data <= 32'h2f76be88;
    11'b01110001010: data <= 32'h39dfb423;
    11'b01110001011: data <= 32'h38a6b481;
    11'b01110001100: data <= 32'h3787bd27;
    11'b01110001101: data <= 32'h3606bc80;
    11'b01110001110: data <= 32'hb86538ee;
    11'b01110001111: data <= 32'hbfff3f4d;
    11'b01110010000: data <= 32'hc0a63bdb;
    11'b01110010001: data <= 32'hbbeab955;
    11'b01110010010: data <= 32'h3518bc45;
    11'b01110010011: data <= 32'h2e2db16b;
    11'b01110010100: data <= 32'hb92638eb;
    11'b01110010101: data <= 32'h1a3b3ac2;
    11'b01110010110: data <= 32'h3ea33cfe;
    11'b01110010111: data <= 32'h40063f28;
    11'b01110011000: data <= 32'h351a3d8b;
    11'b01110011001: data <= 32'hbd43ac8a;
    11'b01110011010: data <= 32'hbb40bc44;
    11'b01110011011: data <= 32'h3a0eb988;
    11'b01110011100: data <= 32'h3e58b158;
    11'b01110011101: data <= 32'h3cb4bb05;
    11'b01110011110: data <= 32'h39e2bfa9;
    11'b01110011111: data <= 32'h3972bd40;
    11'b01110100000: data <= 32'h30fc399f;
    11'b01110100001: data <= 32'hbc0d3e8f;
    11'b01110100010: data <= 32'hbe9133fe;
    11'b01110100011: data <= 32'hbc85be91;
    11'b01110100100: data <= 32'hb89ebf03;
    11'b01110100101: data <= 32'hbb6ab61f;
    11'b01110100110: data <= 32'hbcd43860;
    11'b01110100111: data <= 32'haeb0380c;
    11'b01110101000: data <= 32'h3dfb3932;
    11'b01110101001: data <= 32'h3d903db7;
    11'b01110101010: data <= 32'hb8a43f18;
    11'b01110101011: data <= 32'hbfc43c36;
    11'b01110101100: data <= 32'hbba032c4;
    11'b01110101101: data <= 32'h3c1c2e4c;
    11'b01110101110: data <= 32'h3ebe1f93;
    11'b01110101111: data <= 32'h3bd6bafc;
    11'b01110110000: data <= 32'h393bbe5b;
    11'b01110110001: data <= 32'h3cebb975;
    11'b01110110010: data <= 32'h3d853c92;
    11'b01110110011: data <= 32'h357f3dee;
    11'b01110110100: data <= 32'hba91b5a2;
    11'b01110110101: data <= 32'hbc34c053;
    11'b01110110110: data <= 32'hbacebfa2;
    11'b01110110111: data <= 32'hbc06b770;
    11'b01110111000: data <= 32'hbbb01c22;
    11'b01110111001: data <= 32'h2cf0b91b;
    11'b01110111010: data <= 32'h3ca7b8e2;
    11'b01110111011: data <= 32'h389039f2;
    11'b01110111100: data <= 32'hbd933fb7;
    11'b01110111101: data <= 32'hc0ab3ebd;
    11'b01110111110: data <= 32'hbc4239c5;
    11'b01110111111: data <= 32'h39633393;
    11'b01111000000: data <= 32'h3a8b2c04;
    11'b01111000001: data <= 32'ha809b72e;
    11'b01111000010: data <= 32'h324eb9bd;
    11'b01111000011: data <= 32'h3eae331f;
    11'b01111000100: data <= 32'h40c23e6d;
    11'b01111000101: data <= 32'h3cf33e00;
    11'b01111000110: data <= 32'hb64fb506;
    11'b01111000111: data <= 32'hbb08bede;
    11'b01111001000: data <= 32'hb789bd07;
    11'b01111001001: data <= 32'hb419b41e;
    11'b01111001010: data <= 32'hb165b94b;
    11'b01111001011: data <= 32'h36fabfa8;
    11'b01111001100: data <= 32'h3be2bf1e;
    11'b01111001101: data <= 32'h33e5316a;
    11'b01111001110: data <= 32'hbda43f3e;
    11'b01111001111: data <= 32'hc0253e17;
    11'b01111010000: data <= 32'hbc4633ed;
    11'b01111010001: data <= 32'had38b4d4;
    11'b01111010010: data <= 32'hb862accd;
    11'b01111010011: data <= 32'hbd39a623;
    11'b01111010100: data <= 32'hb613ac06;
    11'b01111010101: data <= 32'h3f063901;
    11'b01111010110: data <= 32'h412e3ea1;
    11'b01111010111: data <= 32'h3ca53e7a;
    11'b01111011000: data <= 32'hb8f135ee;
    11'b01111011001: data <= 32'hba4ab7a8;
    11'b01111011010: data <= 32'h3149ad10;
    11'b01111011011: data <= 32'h39183222;
    11'b01111011100: data <= 32'h3799bc1c;
    11'b01111011101: data <= 32'h391cc121;
    11'b01111011110: data <= 32'h3c4cc050;
    11'b01111011111: data <= 32'h39b62d73;
    11'b01111100000: data <= 32'hb7953e4d;
    11'b01111100001: data <= 32'hbca73a7c;
    11'b01111100010: data <= 32'hbac0b9db;
    11'b01111100011: data <= 32'hb9d1bc15;
    11'b01111100100: data <= 32'hbe5bb40c;
    11'b01111100101: data <= 32'hc02c2cd6;
    11'b01111100110: data <= 32'hb9a1b22b;
    11'b01111100111: data <= 32'h3e0b2d5a;
    11'b01111101000: data <= 32'h3ffe3c5e;
    11'b01111101001: data <= 32'h34ae3e97;
    11'b01111101010: data <= 32'hbd053cee;
    11'b01111101011: data <= 32'hba853a80;
    11'b01111101100: data <= 32'h38793b9f;
    11'b01111101101: data <= 32'h3b513908;
    11'b01111101110: data <= 32'h3576bb48;
    11'b01111101111: data <= 32'h361fc08c;
    11'b01111110000: data <= 32'h3d24be5d;
    11'b01111110001: data <= 32'h3eb1380f;
    11'b01111110010: data <= 32'h3b1c3da1;
    11'b01111110011: data <= 32'had4a2fd5;
    11'b01111110100: data <= 32'hb75dbd99;
    11'b01111110101: data <= 32'hbad5bcf9;
    11'b01111110110: data <= 32'hbed6b240;
    11'b01111110111: data <= 32'hbfc7b128;
    11'b01111111000: data <= 32'hb89cbc50;
    11'b01111111001: data <= 32'h3ca9bcb3;
    11'b01111111010: data <= 32'h3c7b3075;
    11'b01111111011: data <= 32'hb91b3ddd;
    11'b01111111100: data <= 32'hbedf3ebf;
    11'b01111111101: data <= 32'hba923d78;
    11'b01111111110: data <= 32'h37933cf4;
    11'b01111111111: data <= 32'h34ac3a46;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    