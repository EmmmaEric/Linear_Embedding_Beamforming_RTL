
module memory_rom_18(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h3c2f3cc6;
    11'b00000000001: data <= 32'h38b938e6;
    11'b00000000010: data <= 32'hb8d2ba32;
    11'b00000000011: data <= 32'hb692bf51;
    11'b00000000100: data <= 32'h3d07bcc7;
    11'b00000000101: data <= 32'h40ac35cf;
    11'b00000000110: data <= 32'h3e9d39c3;
    11'b00000000111: data <= 32'h349ab7c6;
    11'b00000001000: data <= 32'hb760bd1a;
    11'b00000001001: data <= 32'hbab4b69c;
    11'b00000001010: data <= 32'hbdc038e0;
    11'b00000001011: data <= 32'hbe90aef4;
    11'b00000001100: data <= 32'hb97cbf40;
    11'b00000001101: data <= 32'h3840c027;
    11'b00000001110: data <= 32'h3707b518;
    11'b00000001111: data <= 32'hb9ab3e09;
    11'b00000010000: data <= 32'hbc2b3f4f;
    11'b00000010001: data <= 32'ha2dd3d21;
    11'b00000010010: data <= 32'h38ef3c38;
    11'b00000010011: data <= 32'hb6c23b3e;
    11'b00000010100: data <= 32'hbe9b302b;
    11'b00000010101: data <= 32'hbaf8b95f;
    11'b00000010110: data <= 32'h3dedb669;
    11'b00000010111: data <= 32'h41a03810;
    11'b00000011000: data <= 32'h3fd23877;
    11'b00000011001: data <= 32'h3760b565;
    11'b00000011010: data <= 32'ha347b8b0;
    11'b00000011011: data <= 32'h2f48363a;
    11'b00000011100: data <= 32'hb44a3ae9;
    11'b00000011101: data <= 32'hbac5b8f7;
    11'b00000011110: data <= 32'hb8d7c15e;
    11'b00000011111: data <= 32'h310ac182;
    11'b00000100000: data <= 32'h32f6b98d;
    11'b00000100001: data <= 32'hb6fc3c49;
    11'b00000100010: data <= 32'hb87f3c0b;
    11'b00000100011: data <= 32'h29803464;
    11'b00000100100: data <= 32'hacb736bd;
    11'b00000100101: data <= 32'hbe263c1b;
    11'b00000100110: data <= 32'hc1243a69;
    11'b00000100111: data <= 32'hbd46abb0;
    11'b00000101000: data <= 32'h3ce0b460;
    11'b00000101001: data <= 32'h40a53519;
    11'b00000101010: data <= 32'h3d133908;
    11'b00000101011: data <= 32'h2d5d3618;
    11'b00000101100: data <= 32'h35a33883;
    11'b00000101101: data <= 32'h3c563d6d;
    11'b00000101110: data <= 32'h397b3cfe;
    11'b00000101111: data <= 32'hb6bbb921;
    11'b00000110000: data <= 32'hb911c148;
    11'b00000110001: data <= 32'h32f6c100;
    11'b00000110010: data <= 32'h3a6db8da;
    11'b00000110011: data <= 32'h386f3825;
    11'b00000110100: data <= 32'h343cb0d7;
    11'b00000110101: data <= 32'h33dbbb33;
    11'b00000110110: data <= 32'hb6acb135;
    11'b00000110111: data <= 32'hbfd13c3e;
    11'b00000111000: data <= 32'hc1833b65;
    11'b00000111001: data <= 32'hbdf7b5c7;
    11'b00000111010: data <= 32'h38c8bbc8;
    11'b00000111011: data <= 32'h3ca1b416;
    11'b00000111100: data <= 32'h2c05395b;
    11'b00000111101: data <= 32'hb80d3c17;
    11'b00000111110: data <= 32'h383c3d64;
    11'b00000111111: data <= 32'h3e203f86;
    11'b00001000000: data <= 32'h3a4d3e53;
    11'b00001000001: data <= 32'hba1fade3;
    11'b00001000010: data <= 32'hbb97beb2;
    11'b00001000011: data <= 32'h3765bde5;
    11'b00001000100: data <= 32'h3e9eb11a;
    11'b00001000101: data <= 32'h3e3b2ffb;
    11'b00001000110: data <= 32'h3b9cbbbc;
    11'b00001000111: data <= 32'h38a1bdc7;
    11'b00001001000: data <= 32'had0bb178;
    11'b00001001001: data <= 32'hbd5a3cc8;
    11'b00001001010: data <= 32'hc02638e9;
    11'b00001001011: data <= 32'hbd32bd0b;
    11'b00001001100: data <= 32'ha5e0c00e;
    11'b00001001101: data <= 32'h28dbbb6b;
    11'b00001001110: data <= 32'hbaca37ff;
    11'b00001001111: data <= 32'hba583c11;
    11'b00001010000: data <= 32'h38cd3ca5;
    11'b00001010001: data <= 32'h3d583e66;
    11'b00001010010: data <= 32'h299b3eaf;
    11'b00001010011: data <= 32'hbed039a8;
    11'b00001010100: data <= 32'hbdedb63b;
    11'b00001010101: data <= 32'h386cb5e6;
    11'b00001010110: data <= 32'h40163427;
    11'b00001010111: data <= 32'h3f3da0a4;
    11'b00001011000: data <= 32'h3c1cbc2d;
    11'b00001011001: data <= 32'h3af9bc2a;
    11'b00001011010: data <= 32'h3a453800;
    11'b00001011011: data <= 32'hab0d3e1d;
    11'b00001011100: data <= 32'hbbd93459;
    11'b00001011101: data <= 32'hbb75c005;
    11'b00001011110: data <= 32'hb57bc151;
    11'b00001011111: data <= 32'hb664bd01;
    11'b00001100000: data <= 32'hbb0b3127;
    11'b00001100001: data <= 32'hb785343c;
    11'b00001100010: data <= 32'h39d92acc;
    11'b00001100011: data <= 32'h3abc3982;
    11'b00001100100: data <= 32'hbb5c3e06;
    11'b00001100101: data <= 32'hc1263d36;
    11'b00001100110: data <= 32'hbfad36cf;
    11'b00001100111: data <= 32'h354f2d12;
    11'b00001101000: data <= 32'h3e5a3423;
    11'b00001101001: data <= 32'h3c2410ee;
    11'b00001101010: data <= 32'h3674b852;
    11'b00001101011: data <= 32'h3bb9ac7e;
    11'b00001101100: data <= 32'h3eac3dac;
    11'b00001101101: data <= 32'h3c5b3fc3;
    11'b00001101110: data <= 32'hb31c3434;
    11'b00001101111: data <= 32'hb9e8bfe4;
    11'b00001110000: data <= 32'hb524c0a8;
    11'b00001110001: data <= 32'ha8f1bba4;
    11'b00001110010: data <= 32'hae3db0b6;
    11'b00001110011: data <= 32'h34c8ba7d;
    11'b00001110100: data <= 32'h3beebd34;
    11'b00001110101: data <= 32'h3879b384;
    11'b00001110110: data <= 32'hbd403d28;
    11'b00001110111: data <= 32'hc1673dc1;
    11'b00001111000: data <= 32'hbfb635aa;
    11'b00001111001: data <= 32'had35b61d;
    11'b00001111010: data <= 32'h3802b3a0;
    11'b00001111011: data <= 32'hb56da881;
    11'b00001111100: data <= 32'hb83396c4;
    11'b00001111101: data <= 32'h3af6394e;
    11'b00001111110: data <= 32'h40343f9a;
    11'b00001111111: data <= 32'h3db04051;
    11'b00010000000: data <= 32'hb4cb3930;
    11'b00010000001: data <= 32'hbb95bc4a;
    11'b00010000010: data <= 32'hb10dbc96;
    11'b00010000011: data <= 32'h3961b1bf;
    11'b00010000100: data <= 32'h3a9fb423;
    11'b00010000101: data <= 32'h3ba9be62;
    11'b00010000110: data <= 32'h3d0bc026;
    11'b00010000111: data <= 32'h3a43b84d;
    11'b00010001000: data <= 32'hb9fe3d23;
    11'b00010001001: data <= 32'hbf873ccf;
    11'b00010001010: data <= 32'hbdb6b610;
    11'b00010001011: data <= 32'hb6bcbd51;
    11'b00010001100: data <= 32'hb89cbb1c;
    11'b00010001101: data <= 32'hbdedb206;
    11'b00010001110: data <= 32'hbc882b16;
    11'b00010001111: data <= 32'h3a22381b;
    11'b00010010000: data <= 32'h3fe03e07;
    11'b00010010001: data <= 32'h3aeb3fe6;
    11'b00010010010: data <= 32'hbc643cb7;
    11'b00010010011: data <= 32'hbdd3313d;
    11'b00010010100: data <= 32'had9c3206;
    11'b00010010101: data <= 32'h3c4f38a9;
    11'b00010010110: data <= 32'h3c65b1ea;
    11'b00010010111: data <= 32'h3b95bee0;
    11'b00010011000: data <= 32'h3d4cbf81;
    11'b00010011001: data <= 32'h3d9ba8ed;
    11'b00010011010: data <= 32'h37b33e51;
    11'b00010011011: data <= 32'hb8843b40;
    11'b00010011100: data <= 32'hb99fbc67;
    11'b00010011101: data <= 32'hb807bfd8;
    11'b00010011110: data <= 32'hbc2dbc9d;
    11'b00010011111: data <= 32'hbef0b593;
    11'b00010100000: data <= 32'hbc12b7cc;
    11'b00010100001: data <= 32'h3ab7b858;
    11'b00010100010: data <= 32'h3e24362c;
    11'b00010100011: data <= 32'ha87e3dcc;
    11'b00010100100: data <= 32'hbfcf3e10;
    11'b00010100101: data <= 32'hbf6e3bf6;
    11'b00010100110: data <= 32'hb1cb3b00;
    11'b00010100111: data <= 32'h3a513aa4;
    11'b00010101000: data <= 32'h35f5ada3;
    11'b00010101001: data <= 32'h3050bd22;
    11'b00010101010: data <= 32'h3c48bc01;
    11'b00010101011: data <= 32'h40083ab9;
    11'b00010101100: data <= 32'h3e843fe4;
    11'b00010101101: data <= 32'h37283a88;
    11'b00010101110: data <= 32'hb308bcc3;
    11'b00010101111: data <= 32'hb5c1beb1;
    11'b00010110000: data <= 32'hba05b98e;
    11'b00010110001: data <= 32'hbc52b55e;
    11'b00010110010: data <= 32'hb508bd31;
    11'b00010110011: data <= 32'h3c5cbf91;
    11'b00010110100: data <= 32'h3cdaba64;
    11'b00010110101: data <= 32'hb8253b43;
    11'b00010110110: data <= 32'hc03c3df8;
    11'b00010110111: data <= 32'hbeef3be7;
    11'b00010111000: data <= 32'hb4f13898;
    11'b00010111001: data <= 32'ha9e836f4;
    11'b00010111010: data <= 32'hbbf1af38;
    11'b00010111011: data <= 32'hbc39b9ec;
    11'b00010111100: data <= 32'h3903b2de;
    11'b00010111101: data <= 32'h40843d6f;
    11'b00010111110: data <= 32'h400a402f;
    11'b00010111111: data <= 32'h387e3bac;
    11'b00011000000: data <= 32'hb490b82b;
    11'b00011000001: data <= 32'hb17ab80a;
    11'b00011000010: data <= 32'hac0c356a;
    11'b00011000011: data <= 32'hb06ead6f;
    11'b00011000100: data <= 32'h35fcbf77;
    11'b00011000101: data <= 32'h3d2ec16f;
    11'b00011000110: data <= 32'h3cf5bd4a;
    11'b00011000111: data <= 32'hb12639b3;
    11'b00011001000: data <= 32'hbd453cd2;
    11'b00011001001: data <= 32'hbbed34b5;
    11'b00011001010: data <= 32'hb491b5a4;
    11'b00011001011: data <= 32'hbb24b371;
    11'b00011001100: data <= 32'hc05db35f;
    11'b00011001101: data <= 32'hbfa5b845;
    11'b00011001110: data <= 32'h3495b1e5;
    11'b00011001111: data <= 32'h40173bf5;
    11'b00011010000: data <= 32'h3e0c3ec2;
    11'b00011010001: data <= 32'hb1bd3c8d;
    11'b00011010010: data <= 32'hba4b37a5;
    11'b00011010011: data <= 32'had583b00;
    11'b00011010100: data <= 32'h37263d7c;
    11'b00011010101: data <= 32'h348d3448;
    11'b00011010110: data <= 32'h3678bf84;
    11'b00011010111: data <= 32'h3cb3c126;
    11'b00011011000: data <= 32'h3e1fbb59;
    11'b00011011001: data <= 32'h3aa93bc2;
    11'b00011011010: data <= 32'h29273b2e;
    11'b00011011011: data <= 32'h2590b7f0;
    11'b00011011100: data <= 32'haabdbc6c;
    11'b00011011101: data <= 32'hbce4b85c;
    11'b00011011110: data <= 32'hc100b3dd;
    11'b00011011111: data <= 32'hbfbaba43;
    11'b00011100000: data <= 32'h3484bc0a;
    11'b00011100001: data <= 32'h3e61b111;
    11'b00011100010: data <= 32'h38943afb;
    11'b00011100011: data <= 32'hbc803c87;
    11'b00011100100: data <= 32'hbcf53c96;
    11'b00011100101: data <= 32'hac753e8b;
    11'b00011100110: data <= 32'h369c3f30;
    11'b00011100111: data <= 32'hb32437ca;
    11'b00011101000: data <= 32'hb6d4bda8;
    11'b00011101001: data <= 32'h391bbebe;
    11'b00011101010: data <= 32'h3f282554;
    11'b00011101011: data <= 32'h3f313da4;
    11'b00011101100: data <= 32'h3c8839dc;
    11'b00011101101: data <= 32'h39cfba67;
    11'b00011101110: data <= 32'h3436bc17;
    11'b00011101111: data <= 32'hbb12ad61;
    11'b00011110000: data <= 32'hbf6b2774;
    11'b00011110001: data <= 32'hbcd1bcf4;
    11'b00011110010: data <= 32'h388fc053;
    11'b00011110011: data <= 32'h3ce3bdb5;
    11'b00011110100: data <= 32'hada92ca3;
    11'b00011110101: data <= 32'hbdec3b17;
    11'b00011110110: data <= 32'hbc863c47;
    11'b00011110111: data <= 32'h28843d76;
    11'b00011111000: data <= 32'had2b3dae;
    11'b00011111001: data <= 32'hbd8c3724;
    11'b00011111010: data <= 32'hbecebab3;
    11'b00011111011: data <= 32'hadd1ba09;
    11'b00011111100: data <= 32'h3f1039b8;
    11'b00011111101: data <= 32'h40303e42;
    11'b00011111110: data <= 32'h3d333968;
    11'b00011111111: data <= 32'h39d4b73d;
    11'b00100000000: data <= 32'h3785ab6a;
    11'b00100000001: data <= 32'hb1613c1b;
    11'b00100000010: data <= 32'hba6738a3;
    11'b00100000011: data <= 32'hb5b8be08;
    11'b00100000100: data <= 32'h3a9dc1c0;
    11'b00100000101: data <= 32'h3c58c00b;
    11'b00100000110: data <= 32'ha76cb3ca;
    11'b00100000111: data <= 32'hbb16384d;
    11'b00100001000: data <= 32'hb5273590;
    11'b00100001001: data <= 32'h35c935bd;
    11'b00100001010: data <= 32'hb8dc38f7;
    11'b00100001011: data <= 32'hc0e53446;
    11'b00100001100: data <= 32'hc14ab808;
    11'b00100001101: data <= 32'hb8d1b73f;
    11'b00100001110: data <= 32'h3dc43877;
    11'b00100001111: data <= 32'h3e323c76;
    11'b00100010000: data <= 32'h3812387c;
    11'b00100010001: data <= 32'h302232e3;
    11'b00100010010: data <= 32'h37f53cba;
    11'b00100010011: data <= 32'h37024054;
    11'b00100010100: data <= 32'hb0523c98;
    11'b00100010101: data <= 32'haf81bd74;
    11'b00100010110: data <= 32'h397bc15d;
    11'b00100010111: data <= 32'h3c68be65;
    11'b00100011000: data <= 32'h390a2c76;
    11'b00100011001: data <= 32'h35263468;
    11'b00100011010: data <= 32'h3a76b822;
    11'b00100011011: data <= 32'h3aceb8db;
    11'b00100011100: data <= 32'hb9e52e66;
    11'b00100011101: data <= 32'hc16833d4;
    11'b00100011110: data <= 32'hc15bb810;
    11'b00100011111: data <= 32'hb8cabb97;
    11'b00100100000: data <= 32'h3c0bb6ea;
    11'b00100100001: data <= 32'h386331bd;
    11'b00100100010: data <= 32'hb8f7344d;
    11'b00100100011: data <= 32'hb82f392c;
    11'b00100100100: data <= 32'h37ac3f7e;
    11'b00100100101: data <= 32'h38ee4146;
    11'b00100100110: data <= 32'hb52f3da8;
    11'b00100100111: data <= 32'hba2fbb14;
    11'b00100101000: data <= 32'h2921bef3;
    11'b00100101001: data <= 32'h3c3cb808;
    11'b00100101010: data <= 32'h3d503990;
    11'b00100101011: data <= 32'h3d593111;
    11'b00100101100: data <= 32'h3e5ebc01;
    11'b00100101101: data <= 32'h3d14ba9f;
    11'b00100101110: data <= 32'hb58835f5;
    11'b00100101111: data <= 32'hc00338dd;
    11'b00100110000: data <= 32'hbf4fb946;
    11'b00100110001: data <= 32'hb0cabf40;
    11'b00100110010: data <= 32'h398dbe74;
    11'b00100110011: data <= 32'hb441b9d8;
    11'b00100110100: data <= 32'hbd0fb062;
    11'b00100110101: data <= 32'hb8ee379d;
    11'b00100110110: data <= 32'h392e3e39;
    11'b00100110111: data <= 32'h36a54059;
    11'b00100111000: data <= 32'hbcbe3cfc;
    11'b00100111001: data <= 32'hbfcab5c7;
    11'b00100111010: data <= 32'hba8cb965;
    11'b00100111011: data <= 32'h3a9c3767;
    11'b00100111100: data <= 32'h3df43c3f;
    11'b00100111101: data <= 32'h3dd42c42;
    11'b00100111110: data <= 32'h3e36bb6e;
    11'b00100111111: data <= 32'h3d94b17a;
    11'b00101000000: data <= 32'h35443d7b;
    11'b00101000001: data <= 32'hbab73d2f;
    11'b00101000010: data <= 32'hb9cfb976;
    11'b00101000011: data <= 32'h353ac0b3;
    11'b00101000100: data <= 32'h3866c053;
    11'b00101000101: data <= 32'hb762bc32;
    11'b00101000110: data <= 32'hbbd9b757;
    11'b00101000111: data <= 32'h2c24b351;
    11'b00101001000: data <= 32'h3c713738;
    11'b00101001001: data <= 32'h31213c95;
    11'b00101001010: data <= 32'hc0153ac8;
    11'b00101001011: data <= 32'hc1b2a9ae;
    11'b00101001100: data <= 32'hbd80b079;
    11'b00101001101: data <= 32'h378538f7;
    11'b00101001110: data <= 32'h3b703a17;
    11'b00101001111: data <= 32'h38acb198;
    11'b00101010000: data <= 32'h3a0db85f;
    11'b00101010001: data <= 32'h3cdd3abd;
    11'b00101010010: data <= 32'h3b3640ed;
    11'b00101010011: data <= 32'h28b63fcd;
    11'b00101010100: data <= 32'hb16eb72e;
    11'b00101010101: data <= 32'h35bdc039;
    11'b00101010110: data <= 32'h375dbead;
    11'b00101010111: data <= 32'hadf0b8a3;
    11'b00101011000: data <= 32'ha530b857;
    11'b00101011001: data <= 32'h3c95bc36;
    11'b00101011010: data <= 32'h3eddb9a2;
    11'b00101011011: data <= 32'h317734fc;
    11'b00101011100: data <= 32'hc0713905;
    11'b00101011101: data <= 32'hc1a527cc;
    11'b00101011110: data <= 32'hbd0bb590;
    11'b00101011111: data <= 32'h31bbaea2;
    11'b00101100000: data <= 32'ha8a0af70;
    11'b00101100001: data <= 32'hb9bcb8d8;
    11'b00101100010: data <= 32'hb264b4cc;
    11'b00101100011: data <= 32'h3bdb3db4;
    11'b00101100100: data <= 32'h3c8441c9;
    11'b00101100101: data <= 32'h3011404e;
    11'b00101100110: data <= 32'hb853ac0e;
    11'b00101100111: data <= 32'hb2abbcc0;
    11'b00101101000: data <= 32'h3447b6b8;
    11'b00101101001: data <= 32'h36263557;
    11'b00101101010: data <= 32'h3ae3b6f5;
    11'b00101101011: data <= 32'h3f9cbe3f;
    11'b00101101100: data <= 32'h4040bcc4;
    11'b00101101101: data <= 32'h38293485;
    11'b00101101110: data <= 32'hbe1c3b17;
    11'b00101101111: data <= 32'hbf562656;
    11'b00101110000: data <= 32'hb863bbb7;
    11'b00101110001: data <= 32'h2d56bc80;
    11'b00101110010: data <= 32'hbadcbc09;
    11'b00101110011: data <= 32'hbe77bc35;
    11'b00101110100: data <= 32'hb8ddb7ba;
    11'b00101110101: data <= 32'h3c103c60;
    11'b00101110110: data <= 32'h3c3d40a2;
    11'b00101110111: data <= 32'hb78a3f06;
    11'b00101111000: data <= 32'hbe1f3409;
    11'b00101111001: data <= 32'hbc37b017;
    11'b00101111010: data <= 32'haa4a3a55;
    11'b00101111011: data <= 32'h37ab3c1a;
    11'b00101111100: data <= 32'h3b95b5d3;
    11'b00101111101: data <= 32'h3f1abe67;
    11'b00101111110: data <= 32'h4021ba75;
    11'b00101111111: data <= 32'h3c0d3c48;
    11'b00110000000: data <= 32'hb5e23e38;
    11'b00110000001: data <= 32'hb8002f7b;
    11'b00110000010: data <= 32'h342dbd8e;
    11'b00110000011: data <= 32'h3016be7b;
    11'b00110000100: data <= 32'hbc93bd12;
    11'b00110000101: data <= 32'hbe71bcf8;
    11'b00110000110: data <= 32'hb12dbc2a;
    11'b00110000111: data <= 32'h3dc79b38;
    11'b00110001000: data <= 32'h3b813c47;
    11'b00110001001: data <= 32'hbcb33c1b;
    11'b00110001010: data <= 32'hc0b535c7;
    11'b00110001011: data <= 32'hbe4d37aa;
    11'b00110001100: data <= 32'hb54a3cee;
    11'b00110001101: data <= 32'h25763be7;
    11'b00110001110: data <= 32'h2cdbb865;
    11'b00110001111: data <= 32'h3a47bd71;
    11'b00110010000: data <= 32'h3e4825c1;
    11'b00110010001: data <= 32'h3d774023;
    11'b00110010010: data <= 32'h38824063;
    11'b00110010011: data <= 32'h357e3546;
    11'b00110010100: data <= 32'h38adbcce;
    11'b00110010101: data <= 32'h2fd6bc7a;
    11'b00110010110: data <= 32'hbb56b90e;
    11'b00110010111: data <= 32'hbadebc27;
    11'b00110011000: data <= 32'h3a6cbe9a;
    11'b00110011001: data <= 32'h4019bccd;
    11'b00110011010: data <= 32'h3bccaa93;
    11'b00110011011: data <= 32'hbd7137cb;
    11'b00110011100: data <= 32'hc0a03519;
    11'b00110011101: data <= 32'hbd4d367d;
    11'b00110011110: data <= 32'hb5fb39ee;
    11'b00110011111: data <= 32'hb9f73409;
    11'b00110100000: data <= 32'hbd07bbe3;
    11'b00110100001: data <= 32'hb742bcb7;
    11'b00110100010: data <= 32'h3bfa3893;
    11'b00110100011: data <= 32'h3dc740f3;
    11'b00110100100: data <= 32'h3a364097;
    11'b00110100101: data <= 32'h334b381f;
    11'b00110100110: data <= 32'h321eb739;
    11'b00110100111: data <= 32'hac85310e;
    11'b00110101000: data <= 32'hb84a386b;
    11'b00110101001: data <= 32'haa66b8ab;
    11'b00110101010: data <= 32'h3e1fbff0;
    11'b00110101011: data <= 32'h40c9bf30;
    11'b00110101100: data <= 32'h3cb4b5af;
    11'b00110101101: data <= 32'hba783847;
    11'b00110101110: data <= 32'hbd3334ba;
    11'b00110101111: data <= 32'hb5bfae02;
    11'b00110110000: data <= 32'hb00eb17c;
    11'b00110110001: data <= 32'hbd82b8d0;
    11'b00110110010: data <= 32'hc082bd99;
    11'b00110110011: data <= 32'hbc9cbd12;
    11'b00110110100: data <= 32'h3a41358e;
    11'b00110110101: data <= 32'h3d533f81;
    11'b00110110110: data <= 32'h34e43eae;
    11'b00110110111: data <= 32'hb8f33807;
    11'b00110111000: data <= 32'hb8c836a1;
    11'b00110111001: data <= 32'hb6193dd7;
    11'b00110111010: data <= 32'hb6623e32;
    11'b00110111011: data <= 32'h2f00b34e;
    11'b00110111100: data <= 32'h3d8dbfcc;
    11'b00110111101: data <= 32'h4047be2c;
    11'b00110111110: data <= 32'h3d7a3420;
    11'b00110111111: data <= 32'h31253c7d;
    11'b00111000000: data <= 32'h2f9e3655;
    11'b00111000001: data <= 32'h3a1db81f;
    11'b00111000010: data <= 32'h336eb9a1;
    11'b00111000011: data <= 32'hbe3ebad2;
    11'b00111000100: data <= 32'hc0c2bdbf;
    11'b00111000101: data <= 32'hbb4ebe43;
    11'b00111000110: data <= 32'h3c64b890;
    11'b00111000111: data <= 32'h3ce0386d;
    11'b00111001000: data <= 32'hb5be38fe;
    11'b00111001001: data <= 32'hbdc73469;
    11'b00111001010: data <= 32'hbc763b27;
    11'b00111001011: data <= 32'hb86c4011;
    11'b00111001100: data <= 32'hb9263eff;
    11'b00111001101: data <= 32'hb8cdb439;
    11'b00111001110: data <= 32'h354ebed6;
    11'b00111001111: data <= 32'h3d59ba3c;
    11'b00111010000: data <= 32'h3d803ce5;
    11'b00111010001: data <= 32'h3b913f05;
    11'b00111010010: data <= 32'h3c63384e;
    11'b00111010011: data <= 32'h3d6fb7da;
    11'b00111010100: data <= 32'h36afb57a;
    11'b00111010101: data <= 32'hbd47b13e;
    11'b00111010110: data <= 32'hbedcbb9a;
    11'b00111010111: data <= 32'ha28ebf51;
    11'b00111011000: data <= 32'h3ec2be6f;
    11'b00111011001: data <= 32'h3cdeb99f;
    11'b00111011010: data <= 32'hb947b2f1;
    11'b00111011011: data <= 32'hbe149488;
    11'b00111011100: data <= 32'hbaa03a4a;
    11'b00111011101: data <= 32'hb58b3e97;
    11'b00111011110: data <= 32'hbc563c74;
    11'b00111011111: data <= 32'hbf14b95f;
    11'b00111100000: data <= 32'hbc27be0d;
    11'b00111100001: data <= 32'h370ab104;
    11'b00111100010: data <= 32'h3cb63ee4;
    11'b00111100011: data <= 32'h3c673f58;
    11'b00111100100: data <= 32'h3c6a381b;
    11'b00111100101: data <= 32'h3c6da8e4;
    11'b00111100110: data <= 32'h34753a32;
    11'b00111100111: data <= 32'hbb803c94;
    11'b00111101000: data <= 32'hbaf7b11a;
    11'b00111101001: data <= 32'h3a47bf6d;
    11'b00111101010: data <= 32'h400dc03f;
    11'b00111101011: data <= 32'h3d00bc92;
    11'b00111101100: data <= 32'hb5edb5af;
    11'b00111101101: data <= 32'hb946af4f;
    11'b00111101110: data <= 32'h340b34a2;
    11'b00111101111: data <= 32'h338d39de;
    11'b00111110000: data <= 32'hbd8e32e3;
    11'b00111110001: data <= 32'hc155bc5f;
    11'b00111110010: data <= 32'hbf8bbde6;
    11'b00111110011: data <= 32'h9e26b0fc;
    11'b00111110100: data <= 32'h3b723d14;
    11'b00111110101: data <= 32'h39043c70;
    11'b00111110110: data <= 32'h349a31b6;
    11'b00111110111: data <= 32'h34e037ed;
    11'b00111111000: data <= 32'ha9a73fdc;
    11'b00111111001: data <= 32'hb9b5409a;
    11'b00111111010: data <= 32'hb8313779;
    11'b00111111011: data <= 32'h3a40be92;
    11'b00111111100: data <= 32'h3ec7bf6b;
    11'b00111111101: data <= 32'h3c92b8b6;
    11'b00111111110: data <= 32'h3455329e;
    11'b00111111111: data <= 32'h3923a088;
    11'b01000000000: data <= 32'h3e2cb1fb;
    11'b01000000001: data <= 32'h3b332ac9;
    11'b01000000010: data <= 32'hbd6ab153;
    11'b01000000011: data <= 32'hc186bc52;
    11'b01000000100: data <= 32'hbeedbe06;
    11'b01000000101: data <= 32'h33b2ba11;
    11'b01000000110: data <= 32'h3a6f2c6c;
    11'b01000000111: data <= 32'hac97aebe;
    11'b01000001000: data <= 32'hb932b617;
    11'b01000001001: data <= 32'hb54e39c5;
    11'b01000001010: data <= 32'hb22a40fe;
    11'b01000001011: data <= 32'hb9db413a;
    11'b01000001100: data <= 32'hbb833862;
    11'b01000001101: data <= 32'hb0b6bd6f;
    11'b01000001110: data <= 32'h39d8bc45;
    11'b01000001111: data <= 32'h3a6c3744;
    11'b01000010000: data <= 32'h3a323b87;
    11'b01000010001: data <= 32'h3e473034;
    11'b01000010010: data <= 32'h408fb58a;
    11'b01000010011: data <= 32'h3d0330a8;
    11'b01000010100: data <= 32'hbc213637;
    11'b01000010101: data <= 32'hc028b727;
    11'b01000010110: data <= 32'hba4dbdb2;
    11'b01000010111: data <= 32'h3b47bdfc;
    11'b01000011000: data <= 32'h3a7fbc82;
    11'b01000011001: data <= 32'hb825bc74;
    11'b01000011010: data <= 32'hbbb6bb02;
    11'b01000011011: data <= 32'hb1d937e9;
    11'b01000011100: data <= 32'h304e4030;
    11'b01000011101: data <= 32'hbabb3fe0;
    11'b01000011110: data <= 32'hbf332e02;
    11'b01000011111: data <= 32'hbdcbbcb3;
    11'b01000100000: data <= 32'hb5abb54a;
    11'b01000100001: data <= 32'h356e3ca9;
    11'b01000100010: data <= 32'h3a293ca6;
    11'b01000100011: data <= 32'h3e3d23b2;
    11'b01000100100: data <= 32'h401cb25c;
    11'b01000100101: data <= 32'h3c6d3ba6;
    11'b01000100110: data <= 32'hb9403e7b;
    11'b01000100111: data <= 32'hbc953853;
    11'b01000101000: data <= 32'h3243bc97;
    11'b01000101001: data <= 32'h3d8fbf42;
    11'b01000101010: data <= 32'h3a44be34;
    11'b01000101011: data <= 32'hb806bd4a;
    11'b01000101100: data <= 32'hb66dbc20;
    11'b01000101101: data <= 32'h3a7da352;
    11'b01000101110: data <= 32'h3b4e3c73;
    11'b01000101111: data <= 32'hba8d3b4e;
    11'b01000110000: data <= 32'hc0f1b77b;
    11'b01000110001: data <= 32'hc08ebc69;
    11'b01000110010: data <= 32'hbb4cad9d;
    11'b01000110011: data <= 32'h9e6f3bfe;
    11'b01000110100: data <= 32'h341e3848;
    11'b01000110101: data <= 32'h398ab80b;
    11'b01000110110: data <= 32'h3c869a38;
    11'b01000110111: data <= 32'h393e3f98;
    11'b01000111000: data <= 32'hb6b84183;
    11'b01000111001: data <= 32'hb8b83d43;
    11'b01000111010: data <= 32'h377dba3a;
    11'b01000111011: data <= 32'h3cafbde3;
    11'b01000111100: data <= 32'h3812bbac;
    11'b01000111101: data <= 32'hb259b96b;
    11'b01000111110: data <= 32'h391aba92;
    11'b01000111111: data <= 32'h4029b7d2;
    11'b01001000000: data <= 32'h3f07340b;
    11'b01001000001: data <= 32'hb89d344b;
    11'b01001000010: data <= 32'hc0eab8af;
    11'b01001000011: data <= 32'hc031bbf4;
    11'b01001000100: data <= 32'hb903b5d0;
    11'b01001000101: data <= 32'hac1d2c74;
    11'b01001000110: data <= 32'hb702b93c;
    11'b01001000111: data <= 32'hb652bd11;
    11'b01001001000: data <= 32'h33f3a6f7;
    11'b01001001001: data <= 32'h35c44095;
    11'b01001001010: data <= 32'hb54e421b;
    11'b01001001011: data <= 32'hb98f3d9f;
    11'b01001001100: data <= 32'hb1cfb823;
    11'b01001001101: data <= 32'h33c9b96e;
    11'b01001001110: data <= 32'ha9d932c0;
    11'b01001001111: data <= 32'h255d347b;
    11'b01001010000: data <= 32'h3d9ab836;
    11'b01001010001: data <= 32'h41a0b9c9;
    11'b01001010010: data <= 32'h40552b8f;
    11'b01001010011: data <= 32'hb349384f;
    11'b01001010100: data <= 32'hbf019f71;
    11'b01001010101: data <= 32'hbc2fb997;
    11'b01001010110: data <= 32'h3399ba56;
    11'b01001010111: data <= 32'h2e27bb87;
    11'b01001011000: data <= 32'hbb77beaf;
    11'b01001011001: data <= 32'hbbc5bf79;
    11'b01001011010: data <= 32'h2f10b55e;
    11'b01001011011: data <= 32'h38df3f62;
    11'b01001011100: data <= 32'hb3b340a4;
    11'b01001011101: data <= 32'hbcf03a52;
    11'b01001011110: data <= 32'hbd1bb78e;
    11'b01001011111: data <= 32'hbadc2dcd;
    11'b01001100000: data <= 32'hb9483ca4;
    11'b01001100001: data <= 32'haf903a4d;
    11'b01001100010: data <= 32'h3d4eb851;
    11'b01001100011: data <= 32'h410eba05;
    11'b01001100100: data <= 32'h3f9c3860;
    11'b01001100101: data <= 32'h28613e30;
    11'b01001100110: data <= 32'hba593bf7;
    11'b01001100111: data <= 32'h30f2b387;
    11'b01001101000: data <= 32'h3c00bb69;
    11'b01001101001: data <= 32'h3226bd1d;
    11'b01001101010: data <= 32'hbc46bf61;
    11'b01001101011: data <= 32'hb9cebfd5;
    11'b01001101100: data <= 32'h3aebba1d;
    11'b01001101101: data <= 32'h3d933ab9;
    11'b01001101110: data <= 32'ha1483c47;
    11'b01001101111: data <= 32'hbeb8a9db;
    11'b01001110000: data <= 32'hbfffb857;
    11'b01001110001: data <= 32'hbda03751;
    11'b01001110010: data <= 32'hbbfa3d36;
    11'b01001110011: data <= 32'hb8c436a3;
    11'b01001110100: data <= 32'h36edbc33;
    11'b01001110101: data <= 32'h3db9ba2f;
    11'b01001110110: data <= 32'h3cc63cee;
    11'b01001110111: data <= 32'h2f7e411c;
    11'b01001111000: data <= 32'hb0623f22;
    11'b01001111001: data <= 32'h39d031d2;
    11'b01001111010: data <= 32'h3c35b88c;
    11'b01001111011: data <= 32'haa63b936;
    11'b01001111100: data <= 32'hbbd1bc3a;
    11'b01001111101: data <= 32'h28bdbe13;
    11'b01001111110: data <= 32'h3ff5bc57;
    11'b01001111111: data <= 32'h4088ae50;
    11'b01010000000: data <= 32'h354b3050;
    11'b01010000001: data <= 32'hbe67b735;
    11'b01010000010: data <= 32'hbf15b7e6;
    11'b01010000011: data <= 32'hbc0a3629;
    11'b01010000100: data <= 32'hbaf03950;
    11'b01010000101: data <= 32'hbc9bb8e7;
    11'b01010000110: data <= 32'hb9c1bf67;
    11'b01010000111: data <= 32'h3457bb82;
    11'b01010001000: data <= 32'h38c93e0f;
    11'b01010001001: data <= 32'h2f6e4196;
    11'b01010001010: data <= 32'hab193f2f;
    11'b01010001011: data <= 32'h361334e3;
    11'b01010001100: data <= 32'h34e92f29;
    11'b01010001101: data <= 32'hb9293898;
    11'b01010001110: data <= 32'hbb75311a;
    11'b01010001111: data <= 32'h3931bb5b;
    11'b01010010000: data <= 32'h414fbcd0;
    11'b01010010001: data <= 32'h4145b757;
    11'b01010010010: data <= 32'h38c82e05;
    11'b01010010011: data <= 32'hbbc6ad30;
    11'b01010010100: data <= 32'hb957b15c;
    11'b01010010101: data <= 32'h2dcd30e3;
    11'b01010010110: data <= 32'hb692b125;
    11'b01010010111: data <= 32'hbe0dbe39;
    11'b01010011000: data <= 32'hbdc3c0e4;
    11'b01010011001: data <= 32'hb1dabce2;
    11'b01010011010: data <= 32'h38e03c6d;
    11'b01010011011: data <= 32'h32ee4006;
    11'b01010011100: data <= 32'hb6333bc6;
    11'b01010011101: data <= 32'hb7ff2cbb;
    11'b01010011110: data <= 32'hb9aa39ee;
    11'b01010011111: data <= 32'hbd223e9d;
    11'b01010100000: data <= 32'hbc673be1;
    11'b01010100001: data <= 32'h3898b958;
    11'b01010100010: data <= 32'h40a4bcdb;
    11'b01010100011: data <= 32'h4064b1bb;
    11'b01010100100: data <= 32'h38e83ae1;
    11'b01010100101: data <= 32'hb0c63a8d;
    11'b01010100110: data <= 32'h39343576;
    11'b01010100111: data <= 32'h3cae2e5d;
    11'b01010101000: data <= 32'ha6fbb756;
    11'b01010101001: data <= 32'hbe66bebe;
    11'b01010101010: data <= 32'hbd96c0cd;
    11'b01010101011: data <= 32'h34ebbdc7;
    11'b01010101100: data <= 32'h3d12332c;
    11'b01010101101: data <= 32'h38023936;
    11'b01010101110: data <= 32'hb9acb19d;
    11'b01010101111: data <= 32'hbc93b4cd;
    11'b01010110000: data <= 32'hbcde3c22;
    11'b01010110001: data <= 32'hbe203ff3;
    11'b01010110010: data <= 32'hbdb23b2b;
    11'b01010110011: data <= 32'hb2f4bc18;
    11'b01010110100: data <= 32'h3c81bd24;
    11'b01010110101: data <= 32'h3cbf35aa;
    11'b01010110110: data <= 32'h362b3f05;
    11'b01010110111: data <= 32'h369b3e45;
    11'b01010111000: data <= 32'h3da139b7;
    11'b01010111001: data <= 32'h3e1a35be;
    11'b01010111010: data <= 32'had4c2dec;
    11'b01010111011: data <= 32'hbe2fba7f;
    11'b01010111100: data <= 32'hba74bebf;
    11'b01010111101: data <= 32'h3d26bdd7;
    11'b01010111110: data <= 32'h4031b8db;
    11'b01010111111: data <= 32'h3ab1b762;
    11'b01011000000: data <= 32'hb962bb3a;
    11'b01011000001: data <= 32'hbbb2b78c;
    11'b01011000010: data <= 32'hba003bd7;
    11'b01011000011: data <= 32'hbca63e24;
    11'b01011000100: data <= 32'hbec6294f;
    11'b01011000101: data <= 32'hbd05bf15;
    11'b01011000110: data <= 32'hb27dbde6;
    11'b01011000111: data <= 32'h340d3906;
    11'b01011001000: data <= 32'h30244005;
    11'b01011001001: data <= 32'h37d83e18;
    11'b01011001010: data <= 32'h3d063922;
    11'b01011001011: data <= 32'h3bdf3a4b;
    11'b01011001100: data <= 32'hb8db3cd4;
    11'b01011001101: data <= 32'hbe2d3883;
    11'b01011001110: data <= 32'hb3d8b9ef;
    11'b01011001111: data <= 32'h3fc3bd2d;
    11'b01011010000: data <= 32'h40d8bb81;
    11'b01011010001: data <= 32'h3ba2b9a4;
    11'b01011010010: data <= 32'hb411ba2b;
    11'b01011010011: data <= 32'h2955b3c1;
    11'b01011010100: data <= 32'h37f83a67;
    11'b01011010101: data <= 32'hb5d93a5f;
    11'b01011010110: data <= 32'hbf03bae7;
    11'b01011010111: data <= 32'hbfb4c0ac;
    11'b01011011000: data <= 32'hbaeabe9e;
    11'b01011011001: data <= 32'ha00d3626;
    11'b01011011010: data <= 32'h2e493d40;
    11'b01011011011: data <= 32'h32b43888;
    11'b01011011100: data <= 32'h37e92d8d;
    11'b01011011101: data <= 32'h28803c70;
    11'b01011011110: data <= 32'hbce74070;
    11'b01011011111: data <= 32'hbea03e65;
    11'b01011100000: data <= 32'hb27bb1f1;
    11'b01011100001: data <= 32'h3eb5bc88;
    11'b01011100010: data <= 32'h3f79b997;
    11'b01011100011: data <= 32'h3961ad5b;
    11'b01011100100: data <= 32'h345827b0;
    11'b01011100101: data <= 32'h3d2433f1;
    11'b01011100110: data <= 32'h3f2639d6;
    11'b01011100111: data <= 32'h359736d7;
    11'b01011101000: data <= 32'hbe85bc31;
    11'b01011101001: data <= 32'hbf9fc067;
    11'b01011101010: data <= 32'hb851be78;
    11'b01011101011: data <= 32'h381db310;
    11'b01011101100: data <= 32'h35a62738;
    11'b01011101101: data <= 32'hae5dba52;
    11'b01011101110: data <= 32'hb1aab91a;
    11'b01011101111: data <= 32'hb81c3ca4;
    11'b01011110000: data <= 32'hbda6411f;
    11'b01011110001: data <= 32'hbf0e3ec7;
    11'b01011110010: data <= 32'hb9f3b5d8;
    11'b01011110011: data <= 32'h3877bc9b;
    11'b01011110100: data <= 32'h3944b248;
    11'b01011110101: data <= 32'h2d6b3a65;
    11'b01011110110: data <= 32'h38893a66;
    11'b01011110111: data <= 32'h401238ae;
    11'b01011111000: data <= 32'h40b13a97;
    11'b01011111001: data <= 32'h38173a19;
    11'b01011111010: data <= 32'hbdf8b403;
    11'b01011111011: data <= 32'hbd69bd33;
    11'b01011111100: data <= 32'h364abd19;
    11'b01011111101: data <= 32'h3d5dba28;
    11'b01011111110: data <= 32'h395dbc46;
    11'b01011111111: data <= 32'hb1c5bef5;
    11'b01100000000: data <= 32'hb188bc47;
    11'b01100000001: data <= 32'hafc73be8;
    11'b01100000010: data <= 32'hbb0b404b;
    11'b01100000011: data <= 32'hbec53b5a;
    11'b01100000100: data <= 32'hbdfabc54;
    11'b01100000101: data <= 32'hb9f8bd52;
    11'b01100000110: data <= 32'hb81a30e3;
    11'b01100000111: data <= 32'hb78d3cc5;
    11'b01100001000: data <= 32'h37d63a9f;
    11'b01100001001: data <= 32'h3faf3616;
    11'b01100001010: data <= 32'h3fa93b88;
    11'b01100001011: data <= 32'h2a663e63;
    11'b01100001100: data <= 32'hbdeb3c5f;
    11'b01100001101: data <= 32'hb9feaf11;
    11'b01100001110: data <= 32'h3c98ba32;
    11'b01100001111: data <= 32'h3ef0bb4a;
    11'b01100010000: data <= 32'h3981bd61;
    11'b01100010001: data <= 32'ha80bbf02;
    11'b01100010010: data <= 32'h3888bb8c;
    11'b01100010011: data <= 32'h3c5a3a4b;
    11'b01100010100: data <= 32'h311e3d91;
    11'b01100010101: data <= 32'hbd94aaf6;
    11'b01100010110: data <= 32'hbfc7bed6;
    11'b01100010111: data <= 32'hbdbebdc4;
    11'b01100011000: data <= 32'hbba1305e;
    11'b01100011001: data <= 32'hb93d39e6;
    11'b01100011010: data <= 32'h314dad6a;
    11'b01100011011: data <= 32'h3ca6b683;
    11'b01100011100: data <= 32'h3b743b34;
    11'b01100011101: data <= 32'hb8f640bb;
    11'b01100011110: data <= 32'hbe33404d;
    11'b01100011111: data <= 32'hb82c3943;
    11'b01100100000: data <= 32'h3c6ab690;
    11'b01100100001: data <= 32'h3cefb8ca;
    11'b01100100010: data <= 32'h3239b9ed;
    11'b01100100011: data <= 32'h305ebba0;
    11'b01100100100: data <= 32'h3e3bb6b9;
    11'b01100100101: data <= 32'h40cb398e;
    11'b01100100110: data <= 32'h3c743b04;
    11'b01100100111: data <= 32'hbc13b6f6;
    11'b01100101000: data <= 32'hbf45be8d;
    11'b01100101001: data <= 32'hbc8ebce1;
    11'b01100101010: data <= 32'hb79ab01a;
    11'b01100101011: data <= 32'hb65cb4ad;
    11'b01100101100: data <= 32'hb0efbdd4;
    11'b01100101101: data <= 32'h361fbd8e;
    11'b01100101110: data <= 32'h32c73943;
    11'b01100101111: data <= 32'hbb0b4123;
    11'b01100110000: data <= 32'hbe074090;
    11'b01100110001: data <= 32'hb9fc3884;
    11'b01100110010: data <= 32'h3394b63e;
    11'b01100110011: data <= 32'h2210ad4c;
    11'b01100110100: data <= 32'hb94c32fe;
    11'b01100110101: data <= 32'h2ee9a93b;
    11'b01100110110: data <= 32'h40499583;
    11'b01100110111: data <= 32'h41fe3967;
    11'b01100111000: data <= 32'h3d9f3b70;
    11'b01100111001: data <= 32'hba602f65;
    11'b01100111010: data <= 32'hbcf3b9e4;
    11'b01100111011: data <= 32'hb0f8b8e0;
    11'b01100111100: data <= 32'h3766b554;
    11'b01100111101: data <= 32'h160dbcd0;
    11'b01100111110: data <= 32'hb506c0ea;
    11'b01100111111: data <= 32'h3081bffa;
    11'b01101000000: data <= 32'h35d7359b;
    11'b01101000001: data <= 32'hb5dc4037;
    11'b01101000010: data <= 32'hbcb83de7;
    11'b01101000011: data <= 32'hbc95b349;
    11'b01101000100: data <= 32'hbaeeb91f;
    11'b01101000101: data <= 32'hbcde351c;
    11'b01101000110: data <= 32'hbdbc3a92;
    11'b01101000111: data <= 32'hb0f632e2;
    11'b01101001000: data <= 32'h3fd5b15e;
    11'b01101001001: data <= 32'h411d3882;
    11'b01101001010: data <= 32'h3b453da8;
    11'b01101001011: data <= 32'hbaaa3cfc;
    11'b01101001100: data <= 32'hb8c4381d;
    11'b01101001101: data <= 32'h3a393081;
    11'b01101001110: data <= 32'h3c48b3b4;
    11'b01101001111: data <= 32'h2cf2bd8d;
    11'b01101010000: data <= 32'hb5cbc0f7;
    11'b01101010001: data <= 32'h385dbf84;
    11'b01101010010: data <= 32'h3d683158;
    11'b01101010011: data <= 32'h39d73d48;
    11'b01101010100: data <= 32'hb8e135a9;
    11'b01101010101: data <= 32'hbd49bc37;
    11'b01101010110: data <= 32'hbdc6ba9b;
    11'b01101010111: data <= 32'hbec83775;
    11'b01101011000: data <= 32'hbeb8396f;
    11'b01101011001: data <= 32'hb801b785;
    11'b01101011010: data <= 32'h3cabbbfd;
    11'b01101011011: data <= 32'h3dce33bb;
    11'b01101011100: data <= 32'h2b953f85;
    11'b01101011101: data <= 32'hbbe74058;
    11'b01101011110: data <= 32'hb3953d5d;
    11'b01101011111: data <= 32'h3c1738fe;
    11'b01101100000: data <= 32'h3a663082;
    11'b01101100001: data <= 32'hb712b9f8;
    11'b01101100010: data <= 32'hb785be5e;
    11'b01101100011: data <= 32'h3cdcbcd2;
    11'b01101100100: data <= 32'h41073137;
    11'b01101100101: data <= 32'h3f09399e;
    11'b01101100110: data <= 32'hac16b4b9;
    11'b01101100111: data <= 32'hbc4bbcdd;
    11'b01101101000: data <= 32'hbc63b8ce;
    11'b01101101001: data <= 32'hbca03766;
    11'b01101101010: data <= 32'hbd3ea59a;
    11'b01101101011: data <= 32'hb9eebeba;
    11'b01101101100: data <= 32'h34e8c022;
    11'b01101101101: data <= 32'h37c7b2e3;
    11'b01101101110: data <= 32'hb7083fa7;
    11'b01101101111: data <= 32'hbbbf407a;
    11'b01101110000: data <= 32'hb32d3ce2;
    11'b01101110001: data <= 32'h37c138a5;
    11'b01101110010: data <= 32'hb3fb38cd;
    11'b01101110011: data <= 32'hbd8e3476;
    11'b01101110100: data <= 32'hb9f6b759;
    11'b01101110101: data <= 32'h3e5db862;
    11'b01101110110: data <= 32'h42143231;
    11'b01101110111: data <= 32'h401d3857;
    11'b01101111000: data <= 32'h30cfac74;
    11'b01101111001: data <= 32'hb822b803;
    11'b01101111010: data <= 32'hab282e1f;
    11'b01101111011: data <= 32'ha6d33835;
    11'b01101111100: data <= 32'hb978b987;
    11'b01101111101: data <= 32'hbaa4c132;
    11'b01101111110: data <= 32'haf91c16b;
    11'b01101111111: data <= 32'h3523b892;
    11'b01110000000: data <= 32'hb0223dbc;
    11'b01110000001: data <= 32'hb8913d83;
    11'b01110000010: data <= 32'hb5813446;
    11'b01110000011: data <= 32'hb59d2ff0;
    11'b01110000100: data <= 32'hbd8c3b5d;
    11'b01110000101: data <= 32'hc0753c26;
    11'b01110000110: data <= 32'hbc732eb2;
    11'b01110000111: data <= 32'h3d63b7e0;
    11'b01110001000: data <= 32'h41162888;
    11'b01110001001: data <= 32'h3dba3a02;
    11'b01110001010: data <= 32'habcd3a30;
    11'b01110001011: data <= 32'h29b0392c;
    11'b01110001100: data <= 32'h3c0b3b87;
    11'b01110001101: data <= 32'h3b023a32;
    11'b01110001110: data <= 32'hb5ebba35;
    11'b01110001111: data <= 32'hbb28c124;
    11'b01110010000: data <= 32'h25e8c103;
    11'b01110010001: data <= 32'h3c07b8f7;
    11'b01110010010: data <= 32'h3acb39b9;
    11'b01110010011: data <= 32'h2ef93069;
    11'b01110010100: data <= 32'hb518bab5;
    11'b01110010101: data <= 32'hba51b4f1;
    11'b01110010110: data <= 32'hbf413c37;
    11'b01110010111: data <= 32'hc0dd3c8f;
    11'b01110011000: data <= 32'hbd7fb452;
    11'b01110011001: data <= 32'h38d4bcbd;
    11'b01110011010: data <= 32'h3d53b65c;
    11'b01110011011: data <= 32'h35263bdc;
    11'b01110011100: data <= 32'hb7753e1a;
    11'b01110011101: data <= 32'h35e23db2;
    11'b01110011110: data <= 32'h3ded3db4;
    11'b01110011111: data <= 32'h3b5f3c84;
    11'b01110100000: data <= 32'hb9d2b0f4;
    11'b01110100001: data <= 32'hbc69be58;
    11'b01110100010: data <= 32'h3709be63;
    11'b01110100011: data <= 32'h3fdbb61a;
    11'b01110100100: data <= 32'h3f4e30cc;
    11'b01110100101: data <= 32'h3997b9c1;
    11'b01110100110: data <= 32'ha8dbbd4a;
    11'b01110100111: data <= 32'hb6ebb453;
    11'b01110101000: data <= 32'hbcc83c88;
    11'b01110101001: data <= 32'hbf72399a;
    11'b01110101010: data <= 32'hbd90bd04;
    11'b01110101011: data <= 32'hb244c064;
    11'b01110101100: data <= 32'h318dbb75;
    11'b01110101101: data <= 32'hb8053b6c;
    11'b01110101110: data <= 32'hb9433e31;
    11'b01110101111: data <= 32'h37093cf4;
    11'b01110110000: data <= 32'h3cd33ce8;
    11'b01110110001: data <= 32'h2fbe3d97;
    11'b01110110010: data <= 32'hbe6d3a79;
    11'b01110110011: data <= 32'hbdebb46b;
    11'b01110110100: data <= 32'h396fb8eb;
    11'b01110110101: data <= 32'h40d3af61;
    11'b01110110110: data <= 32'h4025a98e;
    11'b01110110111: data <= 32'h3a74ba0a;
    11'b01110111000: data <= 32'h35f8bb05;
    11'b01110111001: data <= 32'h38763579;
    11'b01110111010: data <= 32'h2e0a3d3e;
    11'b01110111011: data <= 32'hbb5a328b;
    11'b01110111100: data <= 32'hbce8c021;
    11'b01110111101: data <= 32'hb907c199;
    11'b01110111110: data <= 32'hb3edbced;
    11'b01110111111: data <= 32'hb7c13857;
    11'b01111000000: data <= 32'hb5e939c4;
    11'b01111000001: data <= 32'h36fc308c;
    11'b01111000010: data <= 32'h38963797;
    11'b01111000011: data <= 32'hbb153dd8;
    11'b01111000100: data <= 32'hc0d63e37;
    11'b01111000101: data <= 32'hbf5b384a;
    11'b01111000110: data <= 32'h379fb3d2;
    11'b01111000111: data <= 32'h3fb7b042;
    11'b01111001000: data <= 32'h3d4b2b4a;
    11'b01111001001: data <= 32'h354bb065;
    11'b01111001010: data <= 32'h39822f4c;
    11'b01111001011: data <= 32'h3e653ca9;
    11'b01111001100: data <= 32'h3cf23e62;
    11'b01111001101: data <= 32'hb45f3022;
    11'b01111001110: data <= 32'hbc78c00f;
    11'b01111001111: data <= 32'hb8a0c0fc;
    11'b01111010000: data <= 32'h3247bc39;
    11'b01111010001: data <= 32'h34ee29f9;
    11'b01111010010: data <= 32'h3491b7d6;
    11'b01111010011: data <= 32'h3847bcc6;
    11'b01111010100: data <= 32'h3229b4d2;
    11'b01111010101: data <= 32'hbd253d90;
    11'b01111010110: data <= 32'hc1173ee8;
    11'b01111010111: data <= 32'hbfb036a0;
    11'b01111011000: data <= 32'hacd8b9c4;
    11'b01111011001: data <= 32'h39f7b836;
    11'b01111011010: data <= 32'h9df1321d;
    11'b01111011011: data <= 32'hb6b7381c;
    11'b01111011100: data <= 32'h3a473ac7;
    11'b01111011101: data <= 32'h403d3e67;
    11'b01111011110: data <= 32'h3e2b3f4d;
    11'b01111011111: data <= 32'hb62038ca;
    11'b01111100000: data <= 32'hbd0cbc46;
    11'b01111100001: data <= 32'hb452bd85;
    11'b01111100010: data <= 32'h3c0fb7a6;
    11'b01111100011: data <= 32'h3ce0b476;
    11'b01111100100: data <= 32'h3accbd86;
    11'b01111100101: data <= 32'h39f6bfc7;
    11'b01111100110: data <= 32'h3714b856;
    11'b01111100111: data <= 32'hb97f3d81;
    11'b01111101000: data <= 32'hbf2e3d95;
    11'b01111101001: data <= 32'hbe7ab670;
    11'b01111101010: data <= 32'hb90fbe90;
    11'b01111101011: data <= 32'hb6f7bc33;
    11'b01111101100: data <= 32'hbc6a30fb;
    11'b01111101101: data <= 32'hbb5f38c6;
    11'b01111101110: data <= 32'h39da3964;
    11'b01111101111: data <= 32'h3fc93d02;
    11'b01111110000: data <= 32'h3b793f3a;
    11'b01111110001: data <= 32'hbc943d4f;
    11'b01111110010: data <= 32'hbe873416;
    11'b01111110011: data <= 32'haaa7afd4;
    11'b01111110100: data <= 32'h3deb2ffc;
    11'b01111110101: data <= 32'h3de0b509;
    11'b01111110110: data <= 32'h3abdbe0c;
    11'b01111110111: data <= 32'h3b50bedd;
    11'b01111111000: data <= 32'h3cdfad0d;
    11'b01111111001: data <= 32'h38e33e2b;
    11'b01111111010: data <= 32'hb8a53b9e;
    11'b01111111011: data <= 32'hbc67bcc2;
    11'b01111111100: data <= 32'hbb06c07a;
    11'b01111111101: data <= 32'hbb8bbd13;
    11'b01111111110: data <= 32'hbd4ea8e9;
    11'b01111111111: data <= 32'hba8da9bd;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    