
module memory_rom_61(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbc09bcd7;
    11'b00000000001: data <= 32'hb959b974;
    11'b00000000010: data <= 32'h385d395d;
    11'b00000000011: data <= 32'h37be3f38;
    11'b00000000100: data <= 32'hbc8c3d27;
    11'b00000000101: data <= 32'hc0a3b470;
    11'b00000000110: data <= 32'hbef7ba16;
    11'b00000000111: data <= 32'hb5e73639;
    11'b00000001000: data <= 32'h36e13d1b;
    11'b00000001001: data <= 32'h3a72380e;
    11'b00000001010: data <= 32'h3d97b8a8;
    11'b00000001011: data <= 32'h3ea51d95;
    11'b00000001100: data <= 32'h3a363edf;
    11'b00000001101: data <= 32'hb7b14044;
    11'b00000001110: data <= 32'hb7f3377d;
    11'b00000001111: data <= 32'h3919bdb4;
    11'b00000010000: data <= 32'h3c4cbf64;
    11'b00000010001: data <= 32'h2e56bd44;
    11'b00000010010: data <= 32'hb900bc3b;
    11'b00000010011: data <= 32'h3512bb75;
    11'b00000010100: data <= 32'h3e77b249;
    11'b00000010101: data <= 32'h3bfa3929;
    11'b00000010110: data <= 32'hbd4c3741;
    11'b00000010111: data <= 32'hc197b769;
    11'b00000011000: data <= 32'hc01eb8cd;
    11'b00000011001: data <= 32'hb850346a;
    11'b00000011010: data <= 32'h23b238ed;
    11'b00000011011: data <= 32'haf44b4fc;
    11'b00000011100: data <= 32'h3330bb20;
    11'b00000011101: data <= 32'h3a99378a;
    11'b00000011110: data <= 32'h392d412b;
    11'b00000011111: data <= 32'hafb741ac;
    11'b00000100000: data <= 32'hb3f13ada;
    11'b00000100001: data <= 32'h3657bc07;
    11'b00000100010: data <= 32'h38b4bc3d;
    11'b00000100011: data <= 32'h9d04b4e3;
    11'b00000100100: data <= 32'h2441b617;
    11'b00000100101: data <= 32'h3db1bc00;
    11'b00000100110: data <= 32'h4121bac5;
    11'b00000100111: data <= 32'h3de521d4;
    11'b00000101000: data <= 32'hbc4134aa;
    11'b00000101001: data <= 32'hc0a7b472;
    11'b00000101010: data <= 32'hbd7fb913;
    11'b00000101011: data <= 32'hafcdb659;
    11'b00000101100: data <= 32'hb4bcb82f;
    11'b00000101101: data <= 32'hbc3bbd3e;
    11'b00000101110: data <= 32'hba00bd44;
    11'b00000101111: data <= 32'h35ba37a7;
    11'b00000110000: data <= 32'h3946411d;
    11'b00000110001: data <= 32'hb0fb412d;
    11'b00000110010: data <= 32'hba5b39e9;
    11'b00000110011: data <= 32'hb8aab80b;
    11'b00000110100: data <= 32'hb4562cca;
    11'b00000110101: data <= 32'hb4193b20;
    11'b00000110110: data <= 32'h355c340c;
    11'b00000110111: data <= 32'h3f66bc04;
    11'b00000111000: data <= 32'h4188bbde;
    11'b00000111001: data <= 32'h3e87346e;
    11'b00000111010: data <= 32'hb7c23bd2;
    11'b00000111011: data <= 32'hbcc13536;
    11'b00000111100: data <= 32'hb0b6b8ff;
    11'b00000111101: data <= 32'h3831bc08;
    11'b00000111110: data <= 32'hb6e0bd42;
    11'b00000111111: data <= 32'hbe08bf6e;
    11'b00001000000: data <= 32'hbb19be9b;
    11'b00001000001: data <= 32'h3977a997;
    11'b00001000010: data <= 32'h3bfb3e76;
    11'b00001000011: data <= 32'hb5a13e2e;
    11'b00001000100: data <= 32'hbe743387;
    11'b00001000101: data <= 32'hbe61b144;
    11'b00001000110: data <= 32'hbbe63b11;
    11'b00001000111: data <= 32'hb8d73de1;
    11'b00001001000: data <= 32'h210d34a8;
    11'b00001001001: data <= 32'h3d02bc9a;
    11'b00001001010: data <= 32'h4024b9ba;
    11'b00001001011: data <= 32'h3d8e3c94;
    11'b00001001100: data <= 32'h2d364016;
    11'b00001001101: data <= 32'had523c24;
    11'b00001001110: data <= 32'h3a63b6d3;
    11'b00001001111: data <= 32'h3ad3bc04;
    11'b00001010000: data <= 32'hb7efbc92;
    11'b00001010001: data <= 32'hbd64be48;
    11'b00001010010: data <= 32'hb1a0becc;
    11'b00001010011: data <= 32'h3e84ba58;
    11'b00001010100: data <= 32'h3e4c3586;
    11'b00001010101: data <= 32'hb676367e;
    11'b00001010110: data <= 32'hbffeb385;
    11'b00001010111: data <= 32'hbf75aaa3;
    11'b00001011000: data <= 32'hbc443bdf;
    11'b00001011001: data <= 32'hbaf13c65;
    11'b00001011010: data <= 32'hba7cb61a;
    11'b00001011011: data <= 32'ha498be1a;
    11'b00001011100: data <= 32'h3b8cb6b7;
    11'b00001011101: data <= 32'h3bb63f88;
    11'b00001011110: data <= 32'h35e24163;
    11'b00001011111: data <= 32'h35de3d80;
    11'b00001100000: data <= 32'h3ae8aea7;
    11'b00001100001: data <= 32'h384eb495;
    11'b00001100010: data <= 32'hb948a9dd;
    11'b00001100011: data <= 32'hbb34b8fe;
    11'b00001100100: data <= 32'h3a2dbde5;
    11'b00001100101: data <= 32'h410cbd65;
    11'b00001100110: data <= 32'h4015b79e;
    11'b00001100111: data <= 32'hb1d7aceb;
    11'b00001101000: data <= 32'hbe45b40e;
    11'b00001101001: data <= 32'hbc68a93b;
    11'b00001101010: data <= 32'hb692382b;
    11'b00001101011: data <= 32'hbb3630b5;
    11'b00001101100: data <= 32'hbe9abd4b;
    11'b00001101101: data <= 32'hbcaabfea;
    11'b00001101110: data <= 32'h30a4b6d5;
    11'b00001101111: data <= 32'h39ea3f73;
    11'b00001110000: data <= 32'h35a840c2;
    11'b00001110001: data <= 32'h28fb3c3a;
    11'b00001110010: data <= 32'h2e5c30c6;
    11'b00001110011: data <= 32'hb40639f6;
    11'b00001110100: data <= 32'hbbb93d40;
    11'b00001110101: data <= 32'hb9293587;
    11'b00001110110: data <= 32'h3cb1bcda;
    11'b00001110111: data <= 32'h4158bdea;
    11'b00001111000: data <= 32'h4016b6e5;
    11'b00001111001: data <= 32'h31ff35d6;
    11'b00001111010: data <= 32'hb82f3428;
    11'b00001111011: data <= 32'h346e28e9;
    11'b00001111100: data <= 32'h388c23ed;
    11'b00001111101: data <= 32'hba01b8b7;
    11'b00001111110: data <= 32'hc023bf52;
    11'b00001111111: data <= 32'hbe17c068;
    11'b00010000000: data <= 32'h3255ba48;
    11'b00010000001: data <= 32'h3baa3bfb;
    11'b00010000010: data <= 32'h33543cca;
    11'b00010000011: data <= 32'hb91e3368;
    11'b00010000100: data <= 32'hbaa0324e;
    11'b00010000101: data <= 32'hbb843e03;
    11'b00010000110: data <= 32'hbd064037;
    11'b00010000111: data <= 32'hbadc3975;
    11'b00010001000: data <= 32'h3918bcd2;
    11'b00010001001: data <= 32'h3f6bbd18;
    11'b00010001010: data <= 32'h3dff3454;
    11'b00010001011: data <= 32'h37683d42;
    11'b00010001100: data <= 32'h382a3b8e;
    11'b00010001101: data <= 32'h3dc13320;
    11'b00010001110: data <= 32'h3ce1a944;
    11'b00010001111: data <= 32'hb904b761;
    11'b00010010000: data <= 32'hbfd3bdc5;
    11'b00010010001: data <= 32'hbbf7bff2;
    11'b00010010010: data <= 32'h3bf9bd08;
    11'b00010010011: data <= 32'h3e03b285;
    11'b00010010100: data <= 32'h3256b0fa;
    11'b00010010101: data <= 32'hbc24b8a9;
    11'b00010010110: data <= 32'hbc7a2d8c;
    11'b00010010111: data <= 32'hbb8a3e88;
    11'b00010011000: data <= 32'hbd2f3fc0;
    11'b00010011001: data <= 32'hbdb7320d;
    11'b00010011010: data <= 32'hb880be22;
    11'b00010011011: data <= 32'h3827bc16;
    11'b00010011100: data <= 32'h39be3bd2;
    11'b00010011101: data <= 32'h37f33fde;
    11'b00010011110: data <= 32'h3bdd3ced;
    11'b00010011111: data <= 32'h3ee035fc;
    11'b00010100000: data <= 32'h3c7c376e;
    11'b00010100001: data <= 32'hb9c7388d;
    11'b00010100010: data <= 32'hbe42b4d9;
    11'b00010100011: data <= 32'haf5cbd9c;
    11'b00010100100: data <= 32'h3f7dbe29;
    11'b00010100101: data <= 32'h3fc1bc16;
    11'b00010100110: data <= 32'h34c6baf2;
    11'b00010100111: data <= 32'hba33bad9;
    11'b00010101000: data <= 32'hb6ae98fc;
    11'b00010101001: data <= 32'haf4d3ced;
    11'b00010101010: data <= 32'hbbe53c56;
    11'b00010101011: data <= 32'hbff2b9ac;
    11'b00010101100: data <= 32'hbec7bfe0;
    11'b00010101101: data <= 32'hb82abba2;
    11'b00010101110: data <= 32'h32573c56;
    11'b00010101111: data <= 32'h35873ed2;
    11'b00010110000: data <= 32'h39b73a21;
    11'b00010110001: data <= 32'h3c5634fb;
    11'b00010110010: data <= 32'h36733ce0;
    11'b00010110011: data <= 32'hbc103f9b;
    11'b00010110100: data <= 32'hbd193b50;
    11'b00010110101: data <= 32'h35fdba82;
    11'b00010110110: data <= 32'h4022bdfb;
    11'b00010110111: data <= 32'h3f48bc1d;
    11'b00010111000: data <= 32'h363ab8b2;
    11'b00010111001: data <= 32'h20cdb738;
    11'b00010111010: data <= 32'h3b722be0;
    11'b00010111011: data <= 32'h3c7439cb;
    11'b00010111100: data <= 32'hb7c034c2;
    11'b00010111101: data <= 32'hc064bd07;
    11'b00010111110: data <= 32'hc02fc037;
    11'b00010111111: data <= 32'hb941bc4d;
    11'b00011000000: data <= 32'h343d3753;
    11'b00011000001: data <= 32'h320a3872;
    11'b00011000010: data <= 32'h2b83b4d3;
    11'b00011000011: data <= 32'h309d9c02;
    11'b00011000100: data <= 32'hb5113efa;
    11'b00011000101: data <= 32'hbd014176;
    11'b00011000110: data <= 32'hbd303dde;
    11'b00011000111: data <= 32'h2a6fb8db;
    11'b00011001000: data <= 32'h3d24bcec;
    11'b00011001001: data <= 32'h3c32b5d3;
    11'b00011001010: data <= 32'h34d5356c;
    11'b00011001011: data <= 32'h3a7333f9;
    11'b00011001100: data <= 32'h403e32f2;
    11'b00011001101: data <= 32'h40023833;
    11'b00011001110: data <= 32'haf7f33c3;
    11'b00011001111: data <= 32'hbff7bb50;
    11'b00011010000: data <= 32'hbe70bebf;
    11'b00011010001: data <= 32'h2d31bccb;
    11'b00011010010: data <= 32'h3a66b7dd;
    11'b00011010011: data <= 32'h309eba94;
    11'b00011010100: data <= 32'hb6fabd82;
    11'b00011010101: data <= 32'hb4c9b666;
    11'b00011010110: data <= 32'hb5f63f00;
    11'b00011010111: data <= 32'hbc7f4138;
    11'b00011011000: data <= 32'hbe2c3c48;
    11'b00011011001: data <= 32'hbb30bb24;
    11'b00011011010: data <= 32'hac72bbbe;
    11'b00011011011: data <= 32'ha02d367f;
    11'b00011011100: data <= 32'h235c3c72;
    11'b00011011101: data <= 32'h3c7638c1;
    11'b00011011110: data <= 32'h40e9339d;
    11'b00011011111: data <= 32'h401539f0;
    11'b00011100000: data <= 32'hb0223c1e;
    11'b00011100001: data <= 32'hbe53338e;
    11'b00011100010: data <= 32'hb98dba98;
    11'b00011100011: data <= 32'h3c2ebc88;
    11'b00011100100: data <= 32'h3d2dbc84;
    11'b00011100101: data <= 32'h30cfbe62;
    11'b00011100110: data <= 32'hb6c5bf50;
    11'b00011100111: data <= 32'h318fb8f2;
    11'b00011101000: data <= 32'h37453d42;
    11'b00011101001: data <= 32'hb85c3ef9;
    11'b00011101010: data <= 32'hbef82f66;
    11'b00011101011: data <= 32'hbf52bd85;
    11'b00011101100: data <= 32'hbcb2bab0;
    11'b00011101101: data <= 32'hb9f839c2;
    11'b00011101110: data <= 32'hb5123c3f;
    11'b00011101111: data <= 32'h3a5630a2;
    11'b00011110000: data <= 32'h3f51ac9c;
    11'b00011110001: data <= 32'h3d363c8f;
    11'b00011110010: data <= 32'hb765404c;
    11'b00011110011: data <= 32'hbd003e14;
    11'b00011110100: data <= 32'ha85b24aa;
    11'b00011110101: data <= 32'h3dbdbadd;
    11'b00011110110: data <= 32'h3cd5bc3a;
    11'b00011110111: data <= 32'h25e5bd5e;
    11'b00011111000: data <= 32'h24cebdc8;
    11'b00011111001: data <= 32'h3d37b851;
    11'b00011111010: data <= 32'h3efb3a3e;
    11'b00011111011: data <= 32'h33873a8e;
    11'b00011111100: data <= 32'hbeb5b8e3;
    11'b00011111101: data <= 32'hc03ebe45;
    11'b00011111110: data <= 32'hbd6dba30;
    11'b00011111111: data <= 32'hba01369f;
    11'b00100000000: data <= 32'hb7eb3031;
    11'b00100000001: data <= 32'h2f45bbd8;
    11'b00100000010: data <= 32'h3a45b96d;
    11'b00100000011: data <= 32'h36cc3d6f;
    11'b00100000100: data <= 32'hba1641b3;
    11'b00100000101: data <= 32'hbc7f4045;
    11'b00100000110: data <= 32'hac0e358d;
    11'b00100000111: data <= 32'h3afcb836;
    11'b00100001000: data <= 32'h3640b5d5;
    11'b00100001001: data <= 32'hb5b5b577;
    11'b00100001010: data <= 32'h37d2b8e9;
    11'b00100001011: data <= 32'h40b2b501;
    11'b00100001100: data <= 32'h416e3780;
    11'b00100001101: data <= 32'h3a3137f8;
    11'b00100001110: data <= 32'hbd6bb7cd;
    11'b00100001111: data <= 32'hbe65bc7b;
    11'b00100010000: data <= 32'hb895b8e9;
    11'b00100010001: data <= 32'hafabb256;
    11'b00100010010: data <= 32'hb78fbc5b;
    11'b00100010011: data <= 32'hb76fc04c;
    11'b00100010100: data <= 32'h2eacbd29;
    11'b00100010101: data <= 32'h30ca3ccb;
    11'b00100010110: data <= 32'hb90d4158;
    11'b00100010111: data <= 32'hbc6f3ee2;
    11'b00100011000: data <= 32'hb9632055;
    11'b00100011001: data <= 32'hb505b501;
    11'b00100011010: data <= 32'hba243780;
    11'b00100011011: data <= 32'hbb2f3918;
    11'b00100011100: data <= 32'h38b5aadb;
    11'b00100011101: data <= 32'h413ab446;
    11'b00100011110: data <= 32'h41873744;
    11'b00100011111: data <= 32'h3a0f3b9f;
    11'b00100100000: data <= 32'hbbbc37ba;
    11'b00100100001: data <= 32'hb90bb102;
    11'b00100100010: data <= 32'h388cb444;
    11'b00100100011: data <= 32'h38a0b8b7;
    11'b00100100100: data <= 32'hb6b4bf20;
    11'b00100100101: data <= 32'hb931c148;
    11'b00100100110: data <= 32'h3421be3b;
    11'b00100100111: data <= 32'h3a4639fe;
    11'b00100101000: data <= 32'h28b53f07;
    11'b00100101001: data <= 32'hbc0b38ef;
    11'b00100101010: data <= 32'hbd50b954;
    11'b00100101011: data <= 32'hbd4eb3c5;
    11'b00100101100: data <= 32'hbe523b96;
    11'b00100101101: data <= 32'hbd573b1d;
    11'b00100101110: data <= 32'h32b6b4cb;
    11'b00100101111: data <= 32'h3fc1b92b;
    11'b00100110000: data <= 32'h3fa03873;
    11'b00100110001: data <= 32'h34323f19;
    11'b00100110010: data <= 32'hb99e3ea6;
    11'b00100110011: data <= 32'h31693a4b;
    11'b00100110100: data <= 32'h3cf83174;
    11'b00100110101: data <= 32'h39a7b6aa;
    11'b00100110110: data <= 32'hb8b7bdeb;
    11'b00100110111: data <= 32'hb7d8c05b;
    11'b00100111000: data <= 32'h3c50bd68;
    11'b00100111001: data <= 32'h3fd6346f;
    11'b00100111010: data <= 32'h3b7a39b8;
    11'b00100111011: data <= 32'hb9e4b609;
    11'b00100111100: data <= 32'hbde7bc4f;
    11'b00100111101: data <= 32'hbdd6b146;
    11'b00100111110: data <= 32'hbe2d3b40;
    11'b00100111111: data <= 32'hbdbc345c;
    11'b00101000000: data <= 32'hb6bdbd2e;
    11'b00101000001: data <= 32'h3a57bd81;
    11'b00101000010: data <= 32'h3a3d383a;
    11'b00101000011: data <= 32'hb43f4095;
    11'b00101000100: data <= 32'hb8b34073;
    11'b00101000101: data <= 32'h361c3c79;
    11'b00101000110: data <= 32'h3bfa37a6;
    11'b00101000111: data <= 32'h288c3410;
    11'b00101001000: data <= 32'hbc5cb64a;
    11'b00101001001: data <= 32'hb4a2bc7e;
    11'b00101001010: data <= 32'h3fa3bb31;
    11'b00101001011: data <= 32'h41bf8c30;
    11'b00101001100: data <= 32'h3e113194;
    11'b00101001101: data <= 32'hb611b892;
    11'b00101001110: data <= 32'hbb86ba5d;
    11'b00101001111: data <= 32'hb8cd2e9f;
    11'b00101010000: data <= 32'hb9cb389c;
    11'b00101010001: data <= 32'hbccdb9b0;
    11'b00101010010: data <= 32'hbb98c0cf;
    11'b00101010011: data <= 32'had59c023;
    11'b00101010100: data <= 32'h3205346f;
    11'b00101010101: data <= 32'hb5374021;
    11'b00101010110: data <= 32'hb7c43efb;
    11'b00101010111: data <= 32'h2b523909;
    11'b00101011000: data <= 32'h2c483815;
    11'b00101011001: data <= 32'hbc3d3c22;
    11'b00101011010: data <= 32'hbef73a15;
    11'b00101011011: data <= 32'hb554b405;
    11'b00101011100: data <= 32'h402eb91f;
    11'b00101011101: data <= 32'h41bbacb9;
    11'b00101011110: data <= 32'h3d933594;
    11'b00101011111: data <= 32'hb0372fea;
    11'b00101100000: data <= 32'ha4a42ded;
    11'b00101100001: data <= 32'h399538a6;
    11'b00101100010: data <= 32'h346535f3;
    11'b00101100011: data <= 32'hbb56bd27;
    11'b00101100100: data <= 32'hbca7c1b5;
    11'b00101100101: data <= 32'hb261c08e;
    11'b00101100110: data <= 32'h383dad1a;
    11'b00101100111: data <= 32'h33e73cb9;
    11'b00101101000: data <= 32'hb3fc3800;
    11'b00101101001: data <= 32'hb601b541;
    11'b00101101010: data <= 32'hba6d3581;
    11'b00101101011: data <= 32'hbf5b3e12;
    11'b00101101100: data <= 32'hc0573d13;
    11'b00101101101: data <= 32'hb960b211;
    11'b00101101110: data <= 32'h3db5bb2d;
    11'b00101101111: data <= 32'h3f89aea9;
    11'b00101110000: data <= 32'h39203b62;
    11'b00101110001: data <= 32'hae4f3c89;
    11'b00101110010: data <= 32'h3a273c0b;
    11'b00101110011: data <= 32'h3e753c3c;
    11'b00101110100: data <= 32'h39c8387b;
    11'b00101110101: data <= 32'hbb7dbbce;
    11'b00101110110: data <= 32'hbc7bc091;
    11'b00101110111: data <= 32'h35c1bf63;
    11'b00101111000: data <= 32'h3e09b560;
    11'b00101111001: data <= 32'h3c7b311a;
    11'b00101111010: data <= 32'h2ed9b9cd;
    11'b00101111011: data <= 32'hb742bc45;
    11'b00101111100: data <= 32'hbb3833c3;
    11'b00101111101: data <= 32'hbee43e47;
    11'b00101111110: data <= 32'hc02d3b5c;
    11'b00101111111: data <= 32'hbc75bbb8;
    11'b00110000000: data <= 32'h34dfbe60;
    11'b00110000001: data <= 32'h384db3c0;
    11'b00110000010: data <= 32'hb3133d4b;
    11'b00110000011: data <= 32'hb2073e8e;
    11'b00110000100: data <= 32'h3c383d25;
    11'b00110000101: data <= 32'h3e903cf6;
    11'b00110000110: data <= 32'h34bd3c53;
    11'b00110000111: data <= 32'hbd8d2dc5;
    11'b00110001000: data <= 32'hbc2fbc1b;
    11'b00110001001: data <= 32'h3c23bc41;
    11'b00110001010: data <= 32'h40afb63e;
    11'b00110001011: data <= 32'h3eacb6f0;
    11'b00110001100: data <= 32'h364dbcc7;
    11'b00110001101: data <= 32'ha534bc3b;
    11'b00110001110: data <= 32'hab283704;
    11'b00110001111: data <= 32'hb9c53d7d;
    11'b00110010000: data <= 32'hbe2a2fe0;
    11'b00110010001: data <= 32'hbda4bfe2;
    11'b00110010010: data <= 32'hb8d9c089;
    11'b00110010011: data <= 32'hb54db79d;
    11'b00110010100: data <= 32'hb8a53c98;
    11'b00110010101: data <= 32'hb2033ca3;
    11'b00110010110: data <= 32'h3ae13924;
    11'b00110010111: data <= 32'h3b603be7;
    11'b00110011000: data <= 32'hb9633e88;
    11'b00110011001: data <= 32'hc0103d0f;
    11'b00110011010: data <= 32'hbc782fb8;
    11'b00110011011: data <= 32'h3ce1b7ad;
    11'b00110011100: data <= 32'h40a5b541;
    11'b00110011101: data <= 32'h3daeb614;
    11'b00110011110: data <= 32'h365eb9dd;
    11'b00110011111: data <= 32'h398cb526;
    11'b00110100000: data <= 32'h3d063b4e;
    11'b00110100001: data <= 32'h385f3cef;
    11'b00110100010: data <= 32'hbb52b6ab;
    11'b00110100011: data <= 32'hbdd3c0cc;
    11'b00110100100: data <= 32'hbaa1c0c4;
    11'b00110100101: data <= 32'hb3c9b919;
    11'b00110100110: data <= 32'hb22b371c;
    11'b00110100111: data <= 32'h28bdae2f;
    11'b00110101000: data <= 32'h382db894;
    11'b00110101001: data <= 32'h301b378e;
    11'b00110101010: data <= 32'hbdb03fb3;
    11'b00110101011: data <= 32'hc0cd3f75;
    11'b00110101100: data <= 32'hbd403740;
    11'b00110101101: data <= 32'h39a0b81d;
    11'b00110101110: data <= 32'h3d52b53f;
    11'b00110101111: data <= 32'h36d02d30;
    11'b00110110000: data <= 32'h2d91313e;
    11'b00110110001: data <= 32'h3d18386d;
    11'b00110110010: data <= 32'h40803d72;
    11'b00110110011: data <= 32'h3d1e3d54;
    11'b00110110100: data <= 32'hb965b2de;
    11'b00110110101: data <= 32'hbd6abf49;
    11'b00110110110: data <= 32'hb63fbef4;
    11'b00110110111: data <= 32'h38b4b888;
    11'b00110111000: data <= 32'h38f1b5df;
    11'b00110111001: data <= 32'h3633bd92;
    11'b00110111010: data <= 32'h367ebe6f;
    11'b00110111011: data <= 32'ha9932ce6;
    11'b00110111100: data <= 32'hbd343f8b;
    11'b00110111101: data <= 32'hc0463e8c;
    11'b00110111110: data <= 32'hbdd4b097;
    11'b00110111111: data <= 32'hb2e1bc7d;
    11'b00111000000: data <= 32'had1cb789;
    11'b00111000001: data <= 32'hb9ec3799;
    11'b00111000010: data <= 32'hb53639a1;
    11'b00111000011: data <= 32'h3dc13a9f;
    11'b00111000100: data <= 32'h40cb3d9a;
    11'b00111000101: data <= 32'h3c3e3e61;
    11'b00111000110: data <= 32'hbc033947;
    11'b00111000111: data <= 32'hbd23b80d;
    11'b00111001000: data <= 32'h33c7b933;
    11'b00111001001: data <= 32'h3daeb46d;
    11'b00111001010: data <= 32'h3ca9ba85;
    11'b00111001011: data <= 32'h3897bfeb;
    11'b00111001100: data <= 32'h390abf59;
    11'b00111001101: data <= 32'h390c2f33;
    11'b00111001110: data <= 32'hb4073eb9;
    11'b00111001111: data <= 32'hbd2f3b3f;
    11'b00111010000: data <= 32'hbd99bc75;
    11'b00111010001: data <= 32'hbbafbf2a;
    11'b00111010010: data <= 32'hbc44b921;
    11'b00111010011: data <= 32'hbd7a3757;
    11'b00111010100: data <= 32'hb83735f3;
    11'b00111010101: data <= 32'h3ce030bf;
    11'b00111010110: data <= 32'h3f0d3b06;
    11'b00111010111: data <= 32'h31213f31;
    11'b00111011000: data <= 32'hbe883ea0;
    11'b00111011001: data <= 32'hbd493a0f;
    11'b00111011010: data <= 32'h3851336c;
    11'b00111011011: data <= 32'h3e1527d3;
    11'b00111011100: data <= 32'h3b26b9b4;
    11'b00111011101: data <= 32'h3573be7a;
    11'b00111011110: data <= 32'h3c0ebcd2;
    11'b00111011111: data <= 32'h3f0b386e;
    11'b00111100000: data <= 32'h3c833e1d;
    11'b00111100001: data <= 32'hb59d34c1;
    11'b00111100010: data <= 32'hbca4be8c;
    11'b00111100011: data <= 32'hbc6fbf96;
    11'b00111100100: data <= 32'hbc60b8d5;
    11'b00111100101: data <= 32'hbc812ab7;
    11'b00111100110: data <= 32'hb5cdb9a9;
    11'b00111100111: data <= 32'h3b09bcb0;
    11'b00111101000: data <= 32'h3b802857;
    11'b00111101001: data <= 32'hb9443f17;
    11'b00111101010: data <= 32'hc0024050;
    11'b00111101011: data <= 32'hbd703cdd;
    11'b00111101100: data <= 32'h348c362e;
    11'b00111101101: data <= 32'h39923025;
    11'b00111101110: data <= 32'hb241b405;
    11'b00111101111: data <= 32'hb4bfb9cc;
    11'b00111110000: data <= 32'h3d0ab49a;
    11'b00111110001: data <= 32'h41463c10;
    11'b00111110010: data <= 32'h3ffd3e0b;
    11'b00111110011: data <= 32'h2fcb346c;
    11'b00111110100: data <= 32'hbb50bcdd;
    11'b00111110101: data <= 32'hb94abcae;
    11'b00111110110: data <= 32'hb4b5b30c;
    11'b00111110111: data <= 32'hb4e6b6b4;
    11'b00111111000: data <= 32'h1acabf7e;
    11'b00111111001: data <= 32'h397ac0b4;
    11'b00111111010: data <= 32'h38a8b90f;
    11'b00111111011: data <= 32'hb97b3e2e;
    11'b00111111100: data <= 32'hbeba3f9e;
    11'b00111111101: data <= 32'hbcdb396d;
    11'b00111111110: data <= 32'hb4cab222;
    11'b00111111111: data <= 32'hb89ea4db;
    11'b01000000000: data <= 32'hbe0c321c;
    11'b01000000001: data <= 32'hbc0da945;
    11'b01000000010: data <= 32'h3cc72ff2;
    11'b01000000011: data <= 32'h417b3c15;
    11'b01000000100: data <= 32'h3f713e14;
    11'b01000000101: data <= 32'hb0473aa5;
    11'b01000000110: data <= 32'hba9da97c;
    11'b01000000111: data <= 32'h17fd2c75;
    11'b01000001000: data <= 32'h3926365c;
    11'b01000001001: data <= 32'h35d0b8ce;
    11'b01000001010: data <= 32'h31c0c0ce;
    11'b01000001011: data <= 32'h398ec160;
    11'b01000001100: data <= 32'h3bacb9bd;
    11'b01000001101: data <= 32'h32fc3d2a;
    11'b01000001110: data <= 32'hb9913c9b;
    11'b01000001111: data <= 32'hba87b5d4;
    11'b01000010000: data <= 32'hba03bbb4;
    11'b01000010001: data <= 32'hbdfcb255;
    11'b01000010010: data <= 32'hc08c358c;
    11'b01000010011: data <= 32'hbd8aaea4;
    11'b01000010100: data <= 32'h3b19b67e;
    11'b01000010101: data <= 32'h402d35f1;
    11'b01000010110: data <= 32'h3b5c3d88;
    11'b01000010111: data <= 32'hbab83e10;
    11'b01000011000: data <= 32'hbb0f3c92;
    11'b01000011001: data <= 32'h36ee3c6f;
    11'b01000011010: data <= 32'h3bde3b69;
    11'b01000011011: data <= 32'h33ccb5ef;
    11'b01000011100: data <= 32'hb0f5c00b;
    11'b01000011101: data <= 32'h3a0dc019;
    11'b01000011110: data <= 32'h3f16b366;
    11'b01000011111: data <= 32'h3e0a3ca1;
    11'b01000100000: data <= 32'h36c73707;
    11'b01000100001: data <= 32'hb4edbc62;
    11'b01000100010: data <= 32'hb9d7bce2;
    11'b01000100011: data <= 32'hbe00ad98;
    11'b01000100100: data <= 32'hc01f338f;
    11'b01000100101: data <= 32'hbcdebaf3;
    11'b01000100110: data <= 32'h3873be84;
    11'b01000100111: data <= 32'h3cbab93d;
    11'b01000101000: data <= 32'had283c36;
    11'b01000101001: data <= 32'hbd743f3b;
    11'b01000101010: data <= 32'hbb003e4c;
    11'b01000101011: data <= 32'h37113d54;
    11'b01000101100: data <= 32'h37663c4a;
    11'b01000101101: data <= 32'hb9ea2e90;
    11'b01000101110: data <= 32'hbbc7bc44;
    11'b01000101111: data <= 32'h3966bbd5;
    11'b01000110000: data <= 32'h40d13607;
    11'b01000110001: data <= 32'h40b13c7b;
    11'b01000110010: data <= 32'h3c043201;
    11'b01000110011: data <= 32'h293fbbbd;
    11'b01000110100: data <= 32'hb3afb8e4;
    11'b01000110101: data <= 32'hb93a3770;
    11'b01000110110: data <= 32'hbc7d2e68;
    11'b01000110111: data <= 32'hb9c0bf17;
    11'b01000111000: data <= 32'h35cfc18c;
    11'b01000111001: data <= 32'h3908bddb;
    11'b01000111010: data <= 32'hb62c3953;
    11'b01000111011: data <= 32'hbcae3de8;
    11'b01000111100: data <= 32'hb8a73bfe;
    11'b01000111101: data <= 32'h321a3967;
    11'b01000111110: data <= 32'hb84a3a89;
    11'b01000111111: data <= 32'hc0083841;
    11'b01001000000: data <= 32'hbf70b2e7;
    11'b01001000001: data <= 32'h3661b4db;
    11'b01001000010: data <= 32'h40ca3839;
    11'b01001000011: data <= 32'h405c3c07;
    11'b01001000100: data <= 32'h39b436bc;
    11'b01001000101: data <= 32'h2badacf1;
    11'b01001000110: data <= 32'h369438ac;
    11'b01001000111: data <= 32'h36c93d19;
    11'b01001001000: data <= 32'hb2ac3180;
    11'b01001001001: data <= 32'hb61ec04f;
    11'b01001001010: data <= 32'h348cc22c;
    11'b01001001011: data <= 32'h39a1be3c;
    11'b01001001100: data <= 32'h334e36ed;
    11'b01001001101: data <= 32'hb3b339c9;
    11'b01001001110: data <= 32'h24dab122;
    11'b01001001111: data <= 32'h2683b510;
    11'b01001010000: data <= 32'hbd1e378f;
    11'b01001010001: data <= 32'hc18839f5;
    11'b01001010010: data <= 32'hc0939553;
    11'b01001010011: data <= 32'h2bc9b853;
    11'b01001010100: data <= 32'h3ee2aa03;
    11'b01001010101: data <= 32'h3c91395f;
    11'b01001010110: data <= 32'hb1e93a5f;
    11'b01001010111: data <= 32'hb1003b47;
    11'b01001011000: data <= 32'h3b003e7a;
    11'b01001011001: data <= 32'h3c0f3fa1;
    11'b01001011010: data <= 32'ha87a37cb;
    11'b01001011011: data <= 32'hb8f4beeb;
    11'b01001011100: data <= 32'h312fc0bc;
    11'b01001011101: data <= 32'h3cc7bb53;
    11'b01001011110: data <= 32'h3d33371c;
    11'b01001011111: data <= 32'h3b0b9f77;
    11'b01001100000: data <= 32'h3965bc7a;
    11'b01001100001: data <= 32'h31fabaeb;
    11'b01001100010: data <= 32'hbcdb3764;
    11'b01001100011: data <= 32'hc0fd3a5a;
    11'b01001100100: data <= 32'hc003b721;
    11'b01001100101: data <= 32'hb0d8be1a;
    11'b01001100110: data <= 32'h3a6ebc49;
    11'b01001100111: data <= 32'hac223128;
    11'b01001101000: data <= 32'hbbf13b2f;
    11'b01001101001: data <= 32'hb4a63cfe;
    11'b01001101010: data <= 32'h3c0f3f3c;
    11'b01001101011: data <= 32'h3a753ff6;
    11'b01001101100: data <= 32'hba203b07;
    11'b01001101101: data <= 32'hbdb3ba17;
    11'b01001101110: data <= 32'haf9bbc73;
    11'b01001101111: data <= 32'h3e67a82a;
    11'b01001110000: data <= 32'h400a3885;
    11'b01001110001: data <= 32'h3dcbb5d4;
    11'b01001110010: data <= 32'h3c11bd2c;
    11'b01001110011: data <= 32'h3922b82a;
    11'b01001110100: data <= 32'hb5983be2;
    11'b01001110101: data <= 32'hbd943ae8;
    11'b01001110110: data <= 32'hbd01bc5b;
    11'b01001110111: data <= 32'hb1b2c110;
    11'b01001111000: data <= 32'h3166bf8c;
    11'b01001111001: data <= 32'hb94cb46a;
    11'b01001111010: data <= 32'hbc523865;
    11'b01001111011: data <= 32'haa3e3924;
    11'b01001111100: data <= 32'h3bba3c11;
    11'b01001111101: data <= 32'h2da33e09;
    11'b01001111110: data <= 32'hbf8a3c93;
    11'b01001111111: data <= 32'hc0a930d7;
    11'b01010000000: data <= 32'hb7e9b102;
    11'b01010000001: data <= 32'h3e13369f;
    11'b01010000010: data <= 32'h3f3d3840;
    11'b01010000011: data <= 32'h3c36b520;
    11'b01010000100: data <= 32'h3acfb992;
    11'b01010000101: data <= 32'h3c9437fa;
    11'b01010000110: data <= 32'h3a353f4a;
    11'b01010000111: data <= 32'hb2d93c4d;
    11'b01010001000: data <= 32'hb8debd6b;
    11'b01010001001: data <= 32'hb0bfc192;
    11'b01010001010: data <= 32'h2ca9bfa3;
    11'b01010001011: data <= 32'hb59db5ff;
    11'b01010001100: data <= 32'hb58fad73;
    11'b01010001101: data <= 32'h38a0b878;
    11'b01010001110: data <= 32'h3bc6b31c;
    11'b01010001111: data <= 32'hb7fa3ad9;
    11'b01010010000: data <= 32'hc1203ce3;
    11'b01010010001: data <= 32'hc171381e;
    11'b01010010010: data <= 32'hba06ad63;
    11'b01010010011: data <= 32'h3b662be0;
    11'b01010010100: data <= 32'h39d531cc;
    11'b01010010101: data <= 32'hac7ab05c;
    11'b01010010110: data <= 32'h35622e57;
    11'b01010010111: data <= 32'h3dd43dcf;
    11'b01010011000: data <= 32'h3dfa40e5;
    11'b01010011001: data <= 32'h34583d78;
    11'b01010011010: data <= 32'hb8c3bbc1;
    11'b01010011011: data <= 32'hb432c00c;
    11'b01010011100: data <= 32'h35d2bc44;
    11'b01010011101: data <= 32'h37fead7a;
    11'b01010011110: data <= 32'h396cb948;
    11'b01010011111: data <= 32'h3d03be83;
    11'b01010100000: data <= 32'h3ca9bc54;
    11'b01010100001: data <= 32'hb6e9388d;
    11'b01010100010: data <= 32'hc0803cef;
    11'b01010100011: data <= 32'hc08b344b;
    11'b01010100100: data <= 32'hb9c1ba95;
    11'b01010100101: data <= 32'h3105baca;
    11'b01010100110: data <= 32'hb89cb5e3;
    11'b01010100111: data <= 32'hbcbfaf81;
    11'b01010101000: data <= 32'hae1d3651;
    11'b01010101001: data <= 32'h3e1f3e66;
    11'b01010101010: data <= 32'h3de640ce;
    11'b01010101011: data <= 32'hb21f3e38;
    11'b01010101100: data <= 32'hbd0bb04f;
    11'b01010101101: data <= 32'hb8b3b96e;
    11'b01010101110: data <= 32'h392b2f97;
    11'b01010101111: data <= 32'h3c8c358e;
    11'b01010110000: data <= 32'h3cd3bb64;
    11'b01010110001: data <= 32'h3e0dbfec;
    11'b01010110010: data <= 32'h3ddfbc18;
    11'b01010110011: data <= 32'h35283b64;
    11'b01010110100: data <= 32'hbc463d5e;
    11'b01010110101: data <= 32'hbce9b328;
    11'b01010110110: data <= 32'hb6d9bed6;
    11'b01010110111: data <= 32'hb5d5be7b;
    11'b01010111000: data <= 32'hbd5fba1d;
    11'b01010111001: data <= 32'hbe50b5ee;
    11'b01010111010: data <= 32'haaeab021;
    11'b01010111011: data <= 32'h3e0439e8;
    11'b01010111100: data <= 32'h3b673ea0;
    11'b01010111101: data <= 32'hbca43e09;
    11'b01010111110: data <= 32'hc03c3935;
    11'b01010111111: data <= 32'hbbaa3702;
    11'b01011000000: data <= 32'h38d33b17;
    11'b01011000001: data <= 32'h3bcc3862;
    11'b01011000010: data <= 32'h3a03bb0f;
    11'b01011000011: data <= 32'h3c79be41;
    11'b01011000100: data <= 32'h3ebab1e2;
    11'b01011000101: data <= 32'h3d433eca;
    11'b01011000110: data <= 32'h34393e4d;
    11'b01011000111: data <= 32'hb400b7a7;
    11'b01011001000: data <= 32'hb029bfeb;
    11'b01011001001: data <= 32'hb703be61;
    11'b01011001010: data <= 32'hbce0b969;
    11'b01011001011: data <= 32'hbc38ba01;
    11'b01011001100: data <= 32'h37debcd0;
    11'b01011001101: data <= 32'h3e32b923;
    11'b01011001110: data <= 32'h36453950;
    11'b01011001111: data <= 32'hbf4d3d2a;
    11'b01011010000: data <= 32'hc0f03bbb;
    11'b01011010001: data <= 32'hbc4d399f;
    11'b01011010010: data <= 32'h33093a36;
    11'b01011010011: data <= 32'h1fd234e8;
    11'b01011010100: data <= 32'hb803b9f3;
    11'b01011010101: data <= 32'h3451bada;
    11'b01011010110: data <= 32'h3eba39d2;
    11'b01011010111: data <= 32'h3fda4098;
    11'b01011011000: data <= 32'h3b8d3f16;
    11'b01011011001: data <= 32'h28fdb416;
    11'b01011011010: data <= 32'hae54bd41;
    11'b01011011011: data <= 32'hb20bb917;
    11'b01011011100: data <= 32'hb7cdac91;
    11'b01011011101: data <= 32'hae79bc0b;
    11'b01011011110: data <= 32'h3c96c05f;
    11'b01011011111: data <= 32'h3ec3bec9;
    11'b01011100000: data <= 32'h35802c89;
    11'b01011100001: data <= 32'hbe5b3c78;
    11'b01011100010: data <= 32'hbfaf39fb;
    11'b01011100011: data <= 32'hba062edd;
    11'b01011100100: data <= 32'hb3cba757;
    11'b01011100101: data <= 32'hbcd1b30b;
    11'b01011100110: data <= 32'hbf40b9af;
    11'b01011100111: data <= 32'hb7e5b7e3;
    11'b01011101000: data <= 32'h3e1e3b7d;
    11'b01011101001: data <= 32'h3fd0405a;
    11'b01011101010: data <= 32'h39263ed4;
    11'b01011101011: data <= 32'hb7be34ba;
    11'b01011101100: data <= 32'hb635ac07;
    11'b01011101101: data <= 32'h2d2139ee;
    11'b01011101110: data <= 32'h318939ae;
    11'b01011101111: data <= 32'h3783bc12;
    11'b01011110000: data <= 32'h3d6bc10e;
    11'b01011110001: data <= 32'h3f25bf45;
    11'b01011110010: data <= 32'h3abf33ca;
    11'b01011110011: data <= 32'hb8013ca7;
    11'b01011110100: data <= 32'hb98a348c;
    11'b01011110101: data <= 32'haeb6ba1b;
    11'b01011110110: data <= 32'hb7c0ba93;
    11'b01011110111: data <= 32'hbfc8b8b3;
    11'b01011111000: data <= 32'hc0ccba74;
    11'b01011111001: data <= 32'hb966ba63;
    11'b01011111010: data <= 32'h3da33149;
    11'b01011111011: data <= 32'h3dbe3d0a;
    11'b01011111100: data <= 32'hb4693d3b;
    11'b01011111101: data <= 32'hbd583a49;
    11'b01011111110: data <= 32'hb9f53c12;
    11'b01011111111: data <= 32'h30ae3ee1;
    11'b01100000000: data <= 32'h320b3cb3;
    11'b01100000001: data <= 32'h2e86bac4;
    11'b01100000010: data <= 32'h3a83c048;
    11'b01100000011: data <= 32'h3ea9bc3b;
    11'b01100000100: data <= 32'h3e273bdf;
    11'b01100000101: data <= 32'h3a4a3d8e;
    11'b01100000110: data <= 32'h3813a906;
    11'b01100000111: data <= 32'h37f5bcae;
    11'b01100001000: data <= 32'hb63dbb04;
    11'b01100001001: data <= 32'hbf64b621;
    11'b01100001010: data <= 32'hbff1bb13;
    11'b01100001011: data <= 32'hb250be54;
    11'b01100001100: data <= 32'h3dc4bca6;
    11'b01100001101: data <= 32'h3aeb28ae;
    11'b01100001110: data <= 32'hbc283a07;
    11'b01100001111: data <= 32'hbf0c3b2b;
    11'b01100010000: data <= 32'hba353d35;
    11'b01100010001: data <= 32'h26833f03;
    11'b01100010010: data <= 32'hb80c3c2d;
    11'b01100010011: data <= 32'hbc5eb972;
    11'b01100010100: data <= 32'hb42fbdaf;
    11'b01100010101: data <= 32'h3d3bad2c;
    11'b01100010110: data <= 32'h3fcc3e97;
    11'b01100010111: data <= 32'h3dea3e1c;
    11'b01100011000: data <= 32'h3bcba88f;
    11'b01100011001: data <= 32'h397eba06;
    11'b01100011010: data <= 32'hadca24a9;
    11'b01100011011: data <= 32'hbc7a36ff;
    11'b01100011100: data <= 32'hbc01ba3f;
    11'b01100011101: data <= 32'h3816c09d;
    11'b01100011110: data <= 32'h3e34c072;
    11'b01100011111: data <= 32'h391eba19;
    11'b01100100000: data <= 32'hbc1a35e9;
    11'b01100100001: data <= 32'hbd2138c3;
    11'b01100100010: data <= 32'hb42239c6;
    11'b01100100011: data <= 32'had4e3ba2;
    11'b01100100100: data <= 32'hbdcd37c3;
    11'b01100100101: data <= 32'hc0ceb911;
    11'b01100100110: data <= 32'hbd04bb5e;
    11'b01100100111: data <= 32'h3b2f3531;
    11'b01100101000: data <= 32'h3f483e6a;
    11'b01100101001: data <= 32'h3ccc3d2f;
    11'b01100101010: data <= 32'h37f631b9;
    11'b01100101011: data <= 32'h365d335c;
    11'b01100101100: data <= 32'h31ee3d91;
    11'b01100101101: data <= 32'hb5bb3ddd;
    11'b01100101110: data <= 32'hb42ab7d5;
    11'b01100101111: data <= 32'h3a70c0fe;
    11'b01100110000: data <= 32'h3e0cc0bc;
    11'b01100110001: data <= 32'h3aa4b96b;
    11'b01100110010: data <= 32'hb27235f9;
    11'b01100110011: data <= 32'hac132fa7;
    11'b01100110100: data <= 32'h392bb300;
    11'b01100110101: data <= 32'h1c8e253c;
    11'b01100110110: data <= 32'hc00526da;
    11'b01100110111: data <= 32'hc20ab90d;
    11'b01100111000: data <= 32'hbe43bb9b;
    11'b01100111001: data <= 32'h397eb20f;
    11'b01100111010: data <= 32'h3d1939ab;
    11'b01100111011: data <= 32'h33813923;
    11'b01100111100: data <= 32'hb7643526;
    11'b01100111101: data <= 32'ha9fc3c6f;
    11'b01100111110: data <= 32'h351240d0;
    11'b01100111111: data <= 32'haeaf4034;
    11'b01101000000: data <= 32'hb617b19e;
    11'b01101000001: data <= 32'h34d0c01e;
    11'b01101000010: data <= 32'h3c9abe53;
    11'b01101000011: data <= 32'h3cae3051;
    11'b01101000100: data <= 32'h3af03961;
    11'b01101000101: data <= 32'h3cb8b3dd;
    11'b01101000110: data <= 32'h3dd5ba9d;
    11'b01101000111: data <= 32'h34abb44c;
    11'b01101001000: data <= 32'hbf59319b;
    11'b01101001001: data <= 32'hc131b7ec;
    11'b01101001010: data <= 32'hbc39bd8a;
    11'b01101001011: data <= 32'h3a27bd26;
    11'b01101001100: data <= 32'h3965b875;
    11'b01101001101: data <= 32'hb996b0fd;
    11'b01101001110: data <= 32'hbc6c321f;
    11'b01101001111: data <= 32'hb0dc3d2b;
    11'b01101010000: data <= 32'h360740e6;
    11'b01101010001: data <= 32'hb7763ff0;
    11'b01101010010: data <= 32'hbd5aa758;
    11'b01101010011: data <= 32'hba7dbd40;
    11'b01101010100: data <= 32'h383cb76b;
    11'b01101010101: data <= 32'h3d323bfe;
    11'b01101010110: data <= 32'h3dbd3b33;
    11'b01101010111: data <= 32'h3eb3b639;
    11'b01101011000: data <= 32'h3edbb9c1;
    11'b01101011001: data <= 32'h38ec362d;
    11'b01101011010: data <= 32'hbc523c13;
    11'b01101011011: data <= 32'hbdfeafc0;
    11'b01101011100: data <= 32'hb16abf33;
    11'b01101011101: data <= 32'h3bcdc066;
    11'b01101011110: data <= 32'h3557bd9e;
    11'b01101011111: data <= 32'hbbc2b947;
    11'b01101100000: data <= 32'hbaf4b1df;
    11'b01101100001: data <= 32'h35f13964;
    11'b01101100010: data <= 32'h38423e42;
    11'b01101100011: data <= 32'hbc563d1b;
    11'b01101100100: data <= 32'hc0f8ad00;
    11'b01101100101: data <= 32'hbf77b9ca;
    11'b01101100110: data <= 32'haa723283;
    11'b01101100111: data <= 32'h3c2d3ccc;
    11'b01101101000: data <= 32'h3c6a397a;
    11'b01101101001: data <= 32'h3c91b6c2;
    11'b01101101010: data <= 32'h3d43ac64;
    11'b01101101011: data <= 32'h3a723e54;
    11'b01101101100: data <= 32'hb405403c;
    11'b01101101101: data <= 32'hb827361c;
    11'b01101101110: data <= 32'h35efbf40;
    11'b01101101111: data <= 32'h3bd4c08e;
    11'b01101110000: data <= 32'h34c9bd2d;
    11'b01101110001: data <= 32'hb79eb8c4;
    11'b01101110010: data <= 32'h3129b8ca;
    11'b01101110011: data <= 32'h3d65b522;
    11'b01101110100: data <= 32'h3ae636b3;
    11'b01101110101: data <= 32'hbdb63899;
    11'b01101110110: data <= 32'hc208b099;
    11'b01101110111: data <= 32'hc05db874;
    11'b01101111000: data <= 32'hb41a23ad;
    11'b01101111001: data <= 32'h382d380d;
    11'b01101111010: data <= 32'h2db6a8c3;
    11'b01101111011: data <= 32'h9631b855;
    11'b01101111100: data <= 32'h391e387b;
    11'b01101111101: data <= 32'h3acd4100;
    11'b01101111110: data <= 32'h316d4194;
    11'b01101111111: data <= 32'hb52b39f9;
    11'b01110000000: data <= 32'h2d82bd6c;
    11'b01110000001: data <= 32'h3886bdc3;
    11'b01110000010: data <= 32'h35e6b53e;
    11'b01110000011: data <= 32'h3513ada9;
    11'b01110000100: data <= 32'h3d32baf2;
    11'b01110000101: data <= 32'h4073bc46;
    11'b01110000110: data <= 32'h3d06b195;
    11'b01110000111: data <= 32'hbcc337cc;
    11'b01110001000: data <= 32'hc11524dd;
    11'b01110001001: data <= 32'hbe34b9cc;
    11'b01110001010: data <= 32'h153eba4f;
    11'b01110001011: data <= 32'h234eb920;
    11'b01110001100: data <= 32'hbbb2bb5d;
    11'b01110001101: data <= 32'hbb7abaa3;
    11'b01110001110: data <= 32'h3490391a;
    11'b01110001111: data <= 32'h3b4140fa;
    11'b01110010000: data <= 32'h2b99412c;
    11'b01110010001: data <= 32'hbbc93a16;
    11'b01110010010: data <= 32'hbb21b980;
    11'b01110010011: data <= 32'hb0e9b301;
    11'b01110010100: data <= 32'h34c03a79;
    11'b01110010101: data <= 32'h39e83656;
    11'b01110010110: data <= 32'h3ef5bbd6;
    11'b01110010111: data <= 32'h40e0bcc5;
    11'b01110011000: data <= 32'h3dfd314e;
    11'b01110011001: data <= 32'hb7ce3cb4;
    11'b01110011010: data <= 32'hbd6637d4;
    11'b01110011011: data <= 32'hb691bb42;
    11'b01110011100: data <= 32'h3770be14;
    11'b01110011101: data <= 32'hb45abdba;
    11'b01110011110: data <= 32'hbdc7bdb4;
    11'b01110011111: data <= 32'hbc10bcb8;
    11'b01110100000: data <= 32'h390b29a9;
    11'b01110100001: data <= 32'h3c963e17;
    11'b01110100010: data <= 32'hb4f03e9a;
    11'b01110100011: data <= 32'hbfa13765;
    11'b01110100100: data <= 32'hbf8ab161;
    11'b01110100101: data <= 32'hba323921;
    11'b01110100110: data <= 32'h1ded3d53;
    11'b01110100111: data <= 32'h365b361e;
    11'b01110101000: data <= 32'h3c8abc4f;
    11'b01110101001: data <= 32'h3f62ba61;
    11'b01110101010: data <= 32'h3dd73c80;
    11'b01110101011: data <= 32'h34384069;
    11'b01110101100: data <= 32'hb2343c42;
    11'b01110101101: data <= 32'h3742baa1;
    11'b01110101110: data <= 32'h398fbe32;
    11'b01110101111: data <= 32'hb58dbd0a;
    11'b01110110000: data <= 32'hbcd3bcd9;
    11'b01110110001: data <= 32'hb3c3bd9c;
    11'b01110110010: data <= 32'h3e1bbb00;
    11'b01110110011: data <= 32'h3e4832e8;
    11'b01110110100: data <= 32'hb81c3905;
    11'b01110110101: data <= 32'hc0b630b8;
    11'b01110110110: data <= 32'hc04c225e;
    11'b01110110111: data <= 32'hbb0939a2;
    11'b01110111000: data <= 32'hb5eb3b53;
    11'b01110111001: data <= 32'hb870b3ab;
    11'b01110111010: data <= 32'hb0e9bd34;
    11'b01110111011: data <= 32'h3ae1b57f;
    11'b01110111100: data <= 32'h3cf63fbb;
    11'b01110111101: data <= 32'h396041ab;
    11'b01110111110: data <= 32'h33e53d82;
    11'b01110111111: data <= 32'h3779b770;
    11'b01111000000: data <= 32'h3684ba08;
    11'b01111000001: data <= 32'hb61db149;
    11'b01111000010: data <= 32'hb8eeb6a8;
    11'b01111000011: data <= 32'h3a0cbda0;
    11'b01111000100: data <= 32'h40bcbe5c;
    11'b01111000101: data <= 32'h3fd5b8e6;
    11'b01111000110: data <= 32'hb50d3318;
    11'b01111000111: data <= 32'hbf9a30e4;
    11'b01111001000: data <= 32'hbd9fabde;
    11'b01111001001: data <= 32'hb5d13000;
    11'b01111001010: data <= 32'hb8feac3c;
    11'b01111001011: data <= 32'hbe3ebc5f;
    11'b01111001100: data <= 32'hbd3fbe80;
    11'b01111001101: data <= 32'h317ab476;
    11'b01111001110: data <= 32'h3c6c3faa;
    11'b01111001111: data <= 32'h39174114;
    11'b01111010000: data <= 32'hb1443cb0;
    11'b01111010001: data <= 32'hb50ba682;
    11'b01111010010: data <= 32'hb46b36b8;
    11'b01111010011: data <= 32'hb8323cbf;
    11'b01111010100: data <= 32'hb4193695;
    11'b01111010101: data <= 32'h3caebd2f;
    11'b01111010110: data <= 32'h4106bf0f;
    11'b01111010111: data <= 32'h400eb827;
    11'b01111011000: data <= 32'h3221397a;
    11'b01111011001: data <= 32'hba033892;
    11'b01111011010: data <= 32'habe9b0d9;
    11'b01111011011: data <= 32'h371bb801;
    11'b01111011100: data <= 32'hb958ba7a;
    11'b01111011101: data <= 32'hc025be36;
    11'b01111011110: data <= 32'hbe94bf6d;
    11'b01111011111: data <= 32'h3429b9bf;
    11'b01111100000: data <= 32'h3d123be3;
    11'b01111100001: data <= 32'h35e93da9;
    11'b01111100010: data <= 32'hbba9384d;
    11'b01111100011: data <= 32'hbcf333ae;
    11'b01111100100: data <= 32'hbaf93d2d;
    11'b01111100101: data <= 32'hba003fdd;
    11'b01111100110: data <= 32'hb7d7397a;
    11'b01111100111: data <= 32'h38c3bd24;
    11'b01111101000: data <= 32'h3f04bde0;
    11'b01111101001: data <= 32'h3eb13455;
    11'b01111101010: data <= 32'h39803e77;
    11'b01111101011: data <= 32'h36813c88;
    11'b01111101100: data <= 32'h3c41adb9;
    11'b01111101101: data <= 32'h3bebb8b8;
    11'b01111101110: data <= 32'hb8cfb942;
    11'b01111101111: data <= 32'hbfb4bccf;
    11'b01111110000: data <= 32'hbc42bf30;
    11'b01111110001: data <= 32'h3c1fbd92;
    11'b01111110010: data <= 32'h3eb7b50b;
    11'b01111110011: data <= 32'h31fe301e;
    11'b01111110100: data <= 32'hbdafaf8d;
    11'b01111110101: data <= 32'hbe0a33de;
    11'b01111110110: data <= 32'hbafa3dc0;
    11'b01111110111: data <= 32'hbb1e3f0f;
    11'b01111111000: data <= 32'hbcdf330f;
    11'b01111111001: data <= 32'hb975bdf5;
    11'b01111111010: data <= 32'h3816bc44;
    11'b01111111011: data <= 32'h3c623c34;
    11'b01111111100: data <= 32'h3b22407b;
    11'b01111111101: data <= 32'h3b553d7d;
    11'b01111111110: data <= 32'h3d422db8;
    11'b01111111111: data <= 32'h3b2f22dd;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    