
module memory_rom_1(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hb34bbe4b;
    11'b00000000001: data <= 32'hb097ba5c;
    11'b00000000010: data <= 32'h2c7d3c18;
    11'b00000000011: data <= 32'hb9933ef7;
    11'b00000000100: data <= 32'hbee633da;
    11'b00000000101: data <= 32'hbef0be7c;
    11'b00000000110: data <= 32'hbbb2bde9;
    11'b00000000111: data <= 32'hb80634b8;
    11'b00000001000: data <= 32'hb4ee3d4a;
    11'b00000001001: data <= 32'h38053a44;
    11'b00000001010: data <= 32'h3e363497;
    11'b00000001011: data <= 32'h3d1b3c1a;
    11'b00000001100: data <= 32'hb7a43f99;
    11'b00000001101: data <= 32'hbe5c3da1;
    11'b00000001110: data <= 32'hb7d3a2a9;
    11'b00000001111: data <= 32'h3ddabb07;
    11'b00000010000: data <= 32'h3f70bb97;
    11'b00000010001: data <= 32'h3978bc47;
    11'b00000010010: data <= 32'h2c99bcdd;
    11'b00000010011: data <= 32'h3b0bb7d3;
    11'b00000010100: data <= 32'h3dc73aa5;
    11'b00000010101: data <= 32'h34ed3c14;
    11'b00000010110: data <= 32'hbdfbb848;
    11'b00000010111: data <= 32'hc01ebff8;
    11'b00000011000: data <= 32'hbd30be06;
    11'b00000011001: data <= 32'hb8782bfe;
    11'b00000011010: data <= 32'hb4e137c0;
    11'b00000011011: data <= 32'h3062b697;
    11'b00000011100: data <= 32'h39a9b86a;
    11'b00000011101: data <= 32'h35623c27;
    11'b00000011110: data <= 32'hbc0a412f;
    11'b00000011111: data <= 32'hbe934059;
    11'b00000100000: data <= 32'hb825369b;
    11'b00000100001: data <= 32'h3bd8b94f;
    11'b00000100010: data <= 32'h3c06b82f;
    11'b00000100011: data <= 32'h2e44b405;
    11'b00000100100: data <= 32'h352db4fa;
    11'b00000100101: data <= 32'h3f912066;
    11'b00000100110: data <= 32'h41263a1f;
    11'b00000100111: data <= 32'h3c043a11;
    11'b00000101000: data <= 32'hbcd9b7be;
    11'b00000101001: data <= 32'hbeffbe3b;
    11'b00000101010: data <= 32'hb96dbccc;
    11'b00000101011: data <= 32'h30bcb5a2;
    11'b00000101100: data <= 32'h1fbbb988;
    11'b00000101101: data <= 32'hb0ecbefe;
    11'b00000101110: data <= 32'h2fe9bd84;
    11'b00000101111: data <= 32'ha4d23aac;
    11'b00000110000: data <= 32'hbba54124;
    11'b00000110001: data <= 32'hbe3d3fae;
    11'b00000110010: data <= 32'hbbd424cc;
    11'b00000110011: data <= 32'hb14ab9df;
    11'b00000110100: data <= 32'hb51c1e8c;
    11'b00000110101: data <= 32'hb99538f3;
    11'b00000110110: data <= 32'h34e735aa;
    11'b00000110111: data <= 32'h40853258;
    11'b00000111000: data <= 32'h41943a23;
    11'b00000111001: data <= 32'h3bd73c7b;
    11'b00000111010: data <= 32'hbc463746;
    11'b00000111011: data <= 32'hbc50b70d;
    11'b00000111100: data <= 32'h35a8b8b6;
    11'b00000111101: data <= 32'h3bdbb8ab;
    11'b00000111110: data <= 32'h346ebdcc;
    11'b00000111111: data <= 32'hb3b1c0d8;
    11'b00001000000: data <= 32'h3373bed3;
    11'b00001000001: data <= 32'h38aa387b;
    11'b00001000010: data <= 32'hb1333fb3;
    11'b00001000011: data <= 32'hbcdf3b67;
    11'b00001000100: data <= 32'hbddbba7d;
    11'b00001000101: data <= 32'hbce9bb86;
    11'b00001000110: data <= 32'hbd55350d;
    11'b00001000111: data <= 32'hbd0e3b0c;
    11'b00001001000: data <= 32'h2571312d;
    11'b00001001001: data <= 32'h3f3fb40d;
    11'b00001001010: data <= 32'h40173957;
    11'b00001001011: data <= 32'h35573f24;
    11'b00001001100: data <= 32'hbc743ebe;
    11'b00001001101: data <= 32'hb80739d1;
    11'b00001001110: data <= 32'h3c0e28f4;
    11'b00001001111: data <= 32'h3cd0b6d8;
    11'b00001010000: data <= 32'h2f16bd50;
    11'b00001010001: data <= 32'hb303c027;
    11'b00001010010: data <= 32'h3b62bd83;
    11'b00001010011: data <= 32'h3f413649;
    11'b00001010100: data <= 32'h3bd53c89;
    11'b00001010101: data <= 32'hb9a2a975;
    11'b00001010110: data <= 32'hbe47bd70;
    11'b00001010111: data <= 32'hbe0abbaa;
    11'b00001011000: data <= 32'hbdbb3549;
    11'b00001011001: data <= 32'hbd2735d7;
    11'b00001011010: data <= 32'hb579bb0e;
    11'b00001011011: data <= 32'h3b4dbce8;
    11'b00001011100: data <= 32'h3b9235f4;
    11'b00001011101: data <= 32'hb5e94072;
    11'b00001011110: data <= 32'hbcb740c6;
    11'b00001011111: data <= 32'hb51a3cec;
    11'b00001100000: data <= 32'h3ab63565;
    11'b00001100001: data <= 32'h381327ce;
    11'b00001100010: data <= 32'hb8cdb774;
    11'b00001100011: data <= 32'hb495bc2f;
    11'b00001100100: data <= 32'h3e9db9ce;
    11'b00001100101: data <= 32'h41bd35be;
    11'b00001100110: data <= 32'h3f21398a;
    11'b00001100111: data <= 32'hb47bb484;
    11'b00001101000: data <= 32'hbcbdbc62;
    11'b00001101001: data <= 32'hbaceb85a;
    11'b00001101010: data <= 32'hb9183378;
    11'b00001101011: data <= 32'hbac8b81e;
    11'b00001101100: data <= 32'hb8bcc045;
    11'b00001101101: data <= 32'h31bcc060;
    11'b00001101110: data <= 32'h3519a688;
    11'b00001101111: data <= 32'hb7f2402b;
    11'b00001110000: data <= 32'hbc0f402f;
    11'b00001110001: data <= 32'hb7903a48;
    11'b00001110010: data <= 32'h981231aa;
    11'b00001110011: data <= 32'hb9d1382e;
    11'b00001110100: data <= 32'hbe313837;
    11'b00001110101: data <= 32'hb854b027;
    11'b00001110110: data <= 32'h3f78b580;
    11'b00001110111: data <= 32'h421734f6;
    11'b00001111000: data <= 32'h3efd3a24;
    11'b00001111001: data <= 32'hb1be358a;
    11'b00001111010: data <= 32'hb849ad0c;
    11'b00001111011: data <= 32'h348a3352;
    11'b00001111100: data <= 32'h36c83466;
    11'b00001111101: data <= 32'hb620bc56;
    11'b00001111110: data <= 32'hb997c18c;
    11'b00001111111: data <= 32'h2751c117;
    11'b00010000000: data <= 32'h38e0b4f0;
    11'b00010000001: data <= 32'h31bb3dbf;
    11'b00010000010: data <= 32'hb81a3c0a;
    11'b00010000011: data <= 32'hb947b3ce;
    11'b00010000100: data <= 32'hbac7b301;
    11'b00010000101: data <= 32'hbed23aa0;
    11'b00010000110: data <= 32'hc0603c15;
    11'b00010000111: data <= 32'hbb23a339;
    11'b00010001000: data <= 32'h3d8bb942;
    11'b00010001001: data <= 32'h40722c32;
    11'b00010001010: data <= 32'h3b7a3c7e;
    11'b00010001011: data <= 32'hb65a3d58;
    11'b00010001100: data <= 32'h258d3c37;
    11'b00010001101: data <= 32'h3c9b3bc7;
    11'b00010001110: data <= 32'h3b95386d;
    11'b00010001111: data <= 32'hb63cbb31;
    11'b00010010000: data <= 32'hba63c0bb;
    11'b00010010001: data <= 32'h368dc02e;
    11'b00010010010: data <= 32'h3e52b547;
    11'b00010010011: data <= 32'h3d1e3957;
    11'b00010010100: data <= 32'h30bfb099;
    11'b00010010101: data <= 32'hb8b8bc59;
    11'b00010010110: data <= 32'hbc23b6a2;
    11'b00010010111: data <= 32'hbf093b7d;
    11'b00010011000: data <= 32'hc0443a71;
    11'b00010011001: data <= 32'hbc96ba45;
    11'b00010011010: data <= 32'h380bbe4f;
    11'b00010011011: data <= 32'h3babb654;
    11'b00010011100: data <= 32'haabb3d5d;
    11'b00010011101: data <= 32'hb9403fa5;
    11'b00010011110: data <= 32'h345b3e1a;
    11'b00010011111: data <= 32'h3d0d3cf9;
    11'b00010100000: data <= 32'h38503b9d;
    11'b00010100001: data <= 32'hbc1fa9b5;
    11'b00010100010: data <= 32'hbc26bcc1;
    11'b00010100011: data <= 32'h3b1bbcaf;
    11'b00010100100: data <= 32'h40f7b132;
    11'b00010100101: data <= 32'h402131e6;
    11'b00010100110: data <= 32'h38c8b942;
    11'b00010100111: data <= 32'hb2b9bc7b;
    11'b00010101000: data <= 32'hb5d5ade4;
    11'b00010101001: data <= 32'hbab63c06;
    11'b00010101010: data <= 32'hbdd1324c;
    11'b00010101011: data <= 32'hbccabf72;
    11'b00010101100: data <= 32'hb3f8c10e;
    11'b00010101101: data <= 32'h2c83baed;
    11'b00010101110: data <= 32'hb7d53c9c;
    11'b00010101111: data <= 32'hb8e13e57;
    11'b00010110000: data <= 32'h345a3bd6;
    11'b00010110001: data <= 32'h39a83b12;
    11'b00010110010: data <= 32'hb8013d0c;
    11'b00010110011: data <= 32'hbfe43ba6;
    11'b00010110100: data <= 32'hbd9ea6ef;
    11'b00010110101: data <= 32'h3c00b785;
    11'b00010110110: data <= 32'h4134ac0f;
    11'b00010110111: data <= 32'h3fcf3008;
    11'b00010111000: data <= 32'h3860b525;
    11'b00010111001: data <= 32'h349bb526;
    11'b00010111010: data <= 32'h3a31395f;
    11'b00010111011: data <= 32'h372d3cc3;
    11'b00010111100: data <= 32'hb95ab33e;
    11'b00010111101: data <= 32'hbc86c0d9;
    11'b00010111110: data <= 32'hb812c1ab;
    11'b00010111111: data <= 32'h2c30bc33;
    11'b00011000000: data <= 32'hab4238eb;
    11'b00011000001: data <= 32'hb02837e8;
    11'b00011000010: data <= 32'h33f2b41b;
    11'b00011000011: data <= 32'h29d431a6;
    11'b00011000100: data <= 32'hbd8c3d82;
    11'b00011000101: data <= 32'hc12d3e24;
    11'b00011000110: data <= 32'hbed83626;
    11'b00011000111: data <= 32'h38aeb81d;
    11'b00011001000: data <= 32'h3f11b434;
    11'b00011001001: data <= 32'h3ba134f9;
    11'b00011001010: data <= 32'h28cb373d;
    11'b00011001011: data <= 32'h3932399b;
    11'b00011001100: data <= 32'h3ed53da7;
    11'b00011001101: data <= 32'h3d0f3deb;
    11'b00011001110: data <= 32'hb61fabd9;
    11'b00011001111: data <= 32'hbc9fbffa;
    11'b00011010000: data <= 32'hb4b7c071;
    11'b00011010001: data <= 32'h3a5cba79;
    11'b00011010010: data <= 32'h3b4b2875;
    11'b00011010011: data <= 32'h385ab9b7;
    11'b00011010100: data <= 32'h360fbd8d;
    11'b00011010101: data <= 32'haf57b551;
    11'b00011010110: data <= 32'hbda63d83;
    11'b00011010111: data <= 32'hc0d03de5;
    11'b00011011000: data <= 32'hbefab003;
    11'b00011011001: data <= 32'hafd6bd1b;
    11'b00011011010: data <= 32'h3744b9ec;
    11'b00011011011: data <= 32'hb50b36d7;
    11'b00011011100: data <= 32'hb8663ba7;
    11'b00011011101: data <= 32'h3a1f3c8c;
    11'b00011011110: data <= 32'h3fd73e63;
    11'b00011011111: data <= 32'h3c873ed3;
    11'b00011100000: data <= 32'hbab2392b;
    11'b00011100001: data <= 32'hbd9cba33;
    11'b00011100010: data <= 32'h2b07bc20;
    11'b00011100011: data <= 32'h3e58b4e9;
    11'b00011100100: data <= 32'h3e9ab4a9;
    11'b00011100101: data <= 32'h3b8cbd6c;
    11'b00011100110: data <= 32'h3926bed9;
    11'b00011100111: data <= 32'h370fb34d;
    11'b00011101000: data <= 32'hb7493dc1;
    11'b00011101001: data <= 32'hbdea3c0c;
    11'b00011101010: data <= 32'hbdddbc3c;
    11'b00011101011: data <= 32'hb9a4c056;
    11'b00011101100: data <= 32'hb867bcc5;
    11'b00011101101: data <= 32'hbc3a34be;
    11'b00011101110: data <= 32'hba0b39a4;
    11'b00011101111: data <= 32'h39de3878;
    11'b00011110000: data <= 32'h3e3c3c13;
    11'b00011110001: data <= 32'h343f3ed4;
    11'b00011110010: data <= 32'hbed23de1;
    11'b00011110011: data <= 32'hbf1937df;
    11'b00011110100: data <= 32'h318da326;
    11'b00011110101: data <= 32'h3ef82cff;
    11'b00011110110: data <= 32'h3e0ab4a4;
    11'b00011110111: data <= 32'h39b1bcb6;
    11'b00011111000: data <= 32'h3aefbc76;
    11'b00011111001: data <= 32'h3da2370f;
    11'b00011111010: data <= 32'h3b6c3e92;
    11'b00011111011: data <= 32'hb5f838ff;
    11'b00011111100: data <= 32'hbc55be7d;
    11'b00011111101: data <= 32'hbb01c0e7;
    11'b00011111110: data <= 32'hb9b6bcf2;
    11'b00011111111: data <= 32'hbadca0df;
    11'b00100000000: data <= 32'hb660b35e;
    11'b00100000001: data <= 32'h39deba1e;
    11'b00100000010: data <= 32'h3bbf9c66;
    11'b00100000011: data <= 32'hb8b63df4;
    11'b00100000100: data <= 32'hc0993fbc;
    11'b00100000101: data <= 32'hbfee3c3c;
    11'b00100000110: data <= 32'hab763298;
    11'b00100000111: data <= 32'h3c282904;
    11'b00100001000: data <= 32'h36f2afd1;
    11'b00100001001: data <= 32'hae5ab808;
    11'b00100001010: data <= 32'h3b1fb10a;
    11'b00100001011: data <= 32'h406a3ca7;
    11'b00100001100: data <= 32'h3f953f7f;
    11'b00100001101: data <= 32'h32973940;
    11'b00100001110: data <= 32'hbb3fbd34;
    11'b00100001111: data <= 32'hb949bf15;
    11'b00100010000: data <= 32'haed4b9bd;
    11'b00100010001: data <= 32'h2212b42c;
    11'b00100010010: data <= 32'h3400bd2f;
    11'b00100010011: data <= 32'h3abac017;
    11'b00100010100: data <= 32'h39cbbaa2;
    11'b00100010101: data <= 32'hb99c3cfd;
    11'b00100010110: data <= 32'hc0233f64;
    11'b00100010111: data <= 32'hbf15397e;
    11'b00100011000: data <= 32'hb751b6bb;
    11'b00100011001: data <= 32'hb022b656;
    11'b00100011010: data <= 32'hbbd9a018;
    11'b00100011011: data <= 32'hbc1428d7;
    11'b00100011100: data <= 32'h39d53576;
    11'b00100011101: data <= 32'h40d33d42;
    11'b00100011110: data <= 32'h3fa53f98;
    11'b00100011111: data <= 32'hacc33c57;
    11'b00100100000: data <= 32'hbc55b320;
    11'b00100100001: data <= 32'hb538b70d;
    11'b00100100010: data <= 32'h39753015;
    11'b00100100011: data <= 32'h3a4bb487;
    11'b00100100100: data <= 32'h3913bf7a;
    11'b00100100101: data <= 32'h3b9bc10e;
    11'b00100100110: data <= 32'h3c28bb81;
    11'b00100100111: data <= 32'h2fd93cd1;
    11'b00100101000: data <= 32'hbc0c3d9b;
    11'b00100101001: data <= 32'hbc9bb2be;
    11'b00100101010: data <= 32'hb9c0bd48;
    11'b00100101011: data <= 32'hbc33babf;
    11'b00100101100: data <= 32'hbf94a797;
    11'b00100101101: data <= 32'hbde9a446;
    11'b00100101110: data <= 32'h386eaf3a;
    11'b00100101111: data <= 32'h400a3906;
    11'b00100110000: data <= 32'h3c703e4b;
    11'b00100110001: data <= 32'hbb593e53;
    11'b00100110010: data <= 32'hbdcf3b97;
    11'b00100110011: data <= 32'hb0653a12;
    11'b00100110100: data <= 32'h3bef3a6f;
    11'b00100110101: data <= 32'h3a12ae38;
    11'b00100110110: data <= 32'h3512bec3;
    11'b00100110111: data <= 32'h3b06c00b;
    11'b00100111000: data <= 32'h3ec0b53b;
    11'b00100111001: data <= 32'h3d9b3d98;
    11'b00100111010: data <= 32'h34813bc9;
    11'b00100111011: data <= 32'hb71abb1a;
    11'b00100111100: data <= 32'hb950bece;
    11'b00100111101: data <= 32'hbcccba9d;
    11'b00100111110: data <= 32'hbf40ad05;
    11'b00100111111: data <= 32'hbce2b938;
    11'b00101000000: data <= 32'h3838bd4f;
    11'b00101000001: data <= 32'h3da4b8a4;
    11'b00101000010: data <= 32'h31aa3c08;
    11'b00101000011: data <= 32'hbe663f24;
    11'b00101000100: data <= 32'hbe7f3df4;
    11'b00101000101: data <= 32'hb0ec3c7f;
    11'b00101000110: data <= 32'h387e3b4e;
    11'b00101000111: data <= 32'hb2a32ff2;
    11'b00101001000: data <= 32'hb959bc0b;
    11'b00101001001: data <= 32'h3860bc15;
    11'b00101001010: data <= 32'h40673772;
    11'b00101001011: data <= 32'h40a93e75;
    11'b00101001100: data <= 32'h3c203aa8;
    11'b00101001101: data <= 32'hac4fba7d;
    11'b00101001110: data <= 32'hb5c0bc87;
    11'b00101001111: data <= 32'hb8c0b0cf;
    11'b00101010000: data <= 32'hbb7c24d7;
    11'b00101010001: data <= 32'hb834bdae;
    11'b00101010010: data <= 32'h3915c11e;
    11'b00101010011: data <= 32'h3c22be62;
    11'b00101010100: data <= 32'hb0cc3827;
    11'b00101010101: data <= 32'hbdee3e46;
    11'b00101010110: data <= 32'hbd1d3c78;
    11'b00101010111: data <= 32'hb3163836;
    11'b00101011000: data <= 32'hb4e8376c;
    11'b00101011001: data <= 32'hbe453378;
    11'b00101011010: data <= 32'hbf2fb5f3;
    11'b00101011011: data <= 32'h2e31b565;
    11'b00101011100: data <= 32'h407839e0;
    11'b00101011101: data <= 32'h40b03e23;
    11'b00101011110: data <= 32'h3a893ba5;
    11'b00101011111: data <= 32'hb2e9a712;
    11'b00101100000: data <= 32'ha5673067;
    11'b00101100001: data <= 32'h34373b4a;
    11'b00101100010: data <= 32'h9fc63515;
    11'b00101100011: data <= 32'ha5d2bf28;
    11'b00101100100: data <= 32'h3965c213;
    11'b00101100101: data <= 32'h3c4fbf3b;
    11'b00101100110: data <= 32'h36343660;
    11'b00101100111: data <= 32'hb7e93c63;
    11'b00101101000: data <= 32'hb7153187;
    11'b00101101001: data <= 32'hb07ab7e2;
    11'b00101101010: data <= 32'hbbfbae16;
    11'b00101101011: data <= 32'hc0f4340a;
    11'b00101101100: data <= 32'hc0cab233;
    11'b00101101101: data <= 32'hb2a9b827;
    11'b00101101110: data <= 32'h3f293023;
    11'b00101101111: data <= 32'h3e083c06;
    11'b00101110000: data <= 32'haf363c66;
    11'b00101110001: data <= 32'hb9733b27;
    11'b00101110010: data <= 32'h31fd3d56;
    11'b00101110011: data <= 32'h3a243f10;
    11'b00101110100: data <= 32'h3306397d;
    11'b00101110101: data <= 32'hb3c8be1c;
    11'b00101110110: data <= 32'h36bec105;
    11'b00101110111: data <= 32'h3d82bc99;
    11'b00101111000: data <= 32'h3d9d394f;
    11'b00101111001: data <= 32'h3a593949;
    11'b00101111010: data <= 32'h3792b954;
    11'b00101111011: data <= 32'h30b9bc70;
    11'b00101111100: data <= 32'hbc22b210;
    11'b00101111101: data <= 32'hc0c535a4;
    11'b00101111110: data <= 32'hc044b7fa;
    11'b00101111111: data <= 32'hb251bdda;
    11'b00110000000: data <= 32'h3cb2bc43;
    11'b00110000001: data <= 32'h370e32c1;
    11'b00110000010: data <= 32'hbc093c1b;
    11'b00110000011: data <= 32'hbbcc3d27;
    11'b00110000100: data <= 32'h34963ecf;
    11'b00110000101: data <= 32'h39273fab;
    11'b00110000110: data <= 32'hb7993b4f;
    11'b00110000111: data <= 32'hbcd1baab;
    11'b00110001000: data <= 32'hb0abbd97;
    11'b00110001001: data <= 32'h3e55b142;
    11'b00110001010: data <= 32'h40513c07;
    11'b00110001011: data <= 32'h3e3b36f0;
    11'b00110001100: data <= 32'h3b8dbaf5;
    11'b00110001101: data <= 32'h3816ba7d;
    11'b00110001110: data <= 32'hb65c3728;
    11'b00110001111: data <= 32'hbdb03972;
    11'b00110010000: data <= 32'hbd17bb84;
    11'b00110010001: data <= 32'h28b6c100;
    11'b00110010010: data <= 32'h39e4c036;
    11'b00110010011: data <= 32'hb07fb6b6;
    11'b00110010100: data <= 32'hbca53990;
    11'b00110010101: data <= 32'hb9823af0;
    11'b00110010110: data <= 32'h36f63c2b;
    11'b00110010111: data <= 32'h2efa3d5e;
    11'b00110011000: data <= 32'hbe803b47;
    11'b00110011001: data <= 32'hc0b8b0f0;
    11'b00110011010: data <= 32'hba39b7c2;
    11'b00110011011: data <= 32'h3dcc35f6;
    11'b00110011100: data <= 32'h40323c0a;
    11'b00110011101: data <= 32'h3d3735d3;
    11'b00110011110: data <= 32'h39bab6b0;
    11'b00110011111: data <= 32'h3a1a3391;
    11'b00110100000: data <= 32'h37d03e27;
    11'b00110100001: data <= 32'hb4a63cc5;
    11'b00110100010: data <= 32'hb810bc62;
    11'b00110100011: data <= 32'h31cec1c3;
    11'b00110100100: data <= 32'h38eec09a;
    11'b00110100101: data <= 32'h2ca7b81b;
    11'b00110100110: data <= 32'hb687345a;
    11'b00110100111: data <= 32'h3177aebd;
    11'b00110101000: data <= 32'h3a00b0ee;
    11'b00110101001: data <= 32'hb5513845;
    11'b00110101010: data <= 32'hc0d63a70;
    11'b00110101011: data <= 32'hc1ef310d;
    11'b00110101100: data <= 32'hbc71b5aa;
    11'b00110101101: data <= 32'h3c06243f;
    11'b00110101110: data <= 32'h3ce93794;
    11'b00110101111: data <= 32'h332d3443;
    11'b00110110000: data <= 32'h26363339;
    11'b00110110001: data <= 32'h3ab63d33;
    11'b00110110010: data <= 32'h3c6540d8;
    11'b00110110011: data <= 32'h337f3e91;
    11'b00110110100: data <= 32'hb772ba4b;
    11'b00110110101: data <= 32'haafbc09e;
    11'b00110110110: data <= 32'h396dbe13;
    11'b00110110111: data <= 32'h3a52aad5;
    11'b00110111000: data <= 32'h39daa8c7;
    11'b00110111001: data <= 32'h3c8bbc1e;
    11'b00110111010: data <= 32'h3caebc35;
    11'b00110111011: data <= 32'hb45e3149;
    11'b00110111100: data <= 32'hc08c3adf;
    11'b00110111101: data <= 32'hc1392cd2;
    11'b00110111110: data <= 32'hbb90bbe6;
    11'b00110111111: data <= 32'h3800bc0c;
    11'b00111000000: data <= 32'h2dafb614;
    11'b00111000001: data <= 32'hbb7d2421;
    11'b00111000010: data <= 32'hb86537ae;
    11'b00111000011: data <= 32'h3aec3e6d;
    11'b00111000100: data <= 32'h3cb44109;
    11'b00111000101: data <= 32'hb09f3f10;
    11'b00111000110: data <= 32'hbcf5b1b4;
    11'b00111000111: data <= 32'hb96ebc88;
    11'b00111001000: data <= 32'h3967b49e;
    11'b00111001001: data <= 32'h3d743890;
    11'b00111001010: data <= 32'h3db3b164;
    11'b00111001011: data <= 32'h3e5abda4;
    11'b00111001100: data <= 32'h3df2bc47;
    11'b00111001101: data <= 32'h34fa38bf;
    11'b00111001110: data <= 32'hbd003ced;
    11'b00111001111: data <= 32'hbe1eb075;
    11'b00111010000: data <= 32'hb708bf3c;
    11'b00111010001: data <= 32'h3196bfe1;
    11'b00111010010: data <= 32'hb934bc1c;
    11'b00111010011: data <= 32'hbd9fb53f;
    11'b00111010100: data <= 32'hb7e62c74;
    11'b00111010101: data <= 32'h3c263b23;
    11'b00111010110: data <= 32'h3afa3f01;
    11'b00111010111: data <= 32'hbc373e0a;
    11'b00111011000: data <= 32'hc09a361c;
    11'b00111011001: data <= 32'hbd6cad16;
    11'b00111011010: data <= 32'h378d3886;
    11'b00111011011: data <= 32'h3d153a9e;
    11'b00111011100: data <= 32'h3c7ab397;
    11'b00111011101: data <= 32'h3cd3bcc1;
    11'b00111011110: data <= 32'h3e15b48b;
    11'b00111011111: data <= 32'h3c533e4d;
    11'b00111100000: data <= 32'h1dd43f39;
    11'b00111100001: data <= 32'hb737b1b1;
    11'b00111100010: data <= 32'ha4dcc03b;
    11'b00111100011: data <= 32'h2d51c03a;
    11'b00111100100: data <= 32'hb948bc0a;
    11'b00111100101: data <= 32'hbb75b8a4;
    11'b00111100110: data <= 32'h3398ba6b;
    11'b00111100111: data <= 32'h3db3b6a4;
    11'b00111101000: data <= 32'h38b1391e;
    11'b00111101001: data <= 32'hbef33c75;
    11'b00111101010: data <= 32'hc1b73919;
    11'b00111101011: data <= 32'hbe7b343a;
    11'b00111101100: data <= 32'h30ad3812;
    11'b00111101101: data <= 32'h379f371d;
    11'b00111101110: data <= 32'habb9b67d;
    11'b00111101111: data <= 32'h3367b9d6;
    11'b00111110000: data <= 32'h3d36391e;
    11'b00111110001: data <= 32'h3e7340d3;
    11'b00111110010: data <= 32'h39d84076;
    11'b00111110011: data <= 32'haddd2c67;
    11'b00111110100: data <= 32'hac6ebe5d;
    11'b00111110101: data <= 32'h2d92bcf9;
    11'b00111110110: data <= 32'hb0bab4b5;
    11'b00111110111: data <= 32'h28d3b8dc;
    11'b00111111000: data <= 32'h3c9ebe8a;
    11'b00111111001: data <= 32'h3f71be00;
    11'b00111111010: data <= 32'h391aab88;
    11'b00111111011: data <= 32'hbe703b97;
    11'b00111111100: data <= 32'hc0da38ba;
    11'b00111111101: data <= 32'hbcf0b0dd;
    11'b00111111110: data <= 32'hae80b521;
    11'b00111111111: data <= 32'hb88db5a4;
    11'b01000000000: data <= 32'hbd97b9a0;
    11'b01000000001: data <= 32'hb970b825;
    11'b01000000010: data <= 32'h3c513b7b;
    11'b01000000011: data <= 32'h3ecc40e4;
    11'b01000000100: data <= 32'h3897405a;
    11'b01000000101: data <= 32'hb9183741;
    11'b01000000110: data <= 32'hb8f2b805;
    11'b01000000111: data <= 32'h243230f0;
    11'b01000001000: data <= 32'h3565395a;
    11'b01000001001: data <= 32'h3987b775;
    11'b01000001010: data <= 32'h3e40c000;
    11'b01000001011: data <= 32'h4018bef7;
    11'b01000001100: data <= 32'h3c292f20;
    11'b01000001101: data <= 32'hb94f3ce0;
    11'b01000001110: data <= 32'hbcc13737;
    11'b01000001111: data <= 32'hb655bac7;
    11'b01000010000: data <= 32'hb084bcd6;
    11'b01000010001: data <= 32'hbd19bbc2;
    11'b01000010010: data <= 32'hc02ebbc2;
    11'b01000010011: data <= 32'hbb49ba5f;
    11'b01000010100: data <= 32'h3c783489;
    11'b01000010101: data <= 32'h3ddd3e2b;
    11'b01000010110: data <= 32'hb1ce3e6c;
    11'b01000010111: data <= 32'hbe6639cc;
    11'b01000011000: data <= 32'hbd163807;
    11'b01000011001: data <= 32'hb1053cf0;
    11'b01000011010: data <= 32'h35323cf5;
    11'b01000011011: data <= 32'h36edb5d9;
    11'b01000011100: data <= 32'h3c44bf59;
    11'b01000011101: data <= 32'h3f30bc86;
    11'b01000011110: data <= 32'h3e203bb8;
    11'b01000011111: data <= 32'h384a3f13;
    11'b01000100000: data <= 32'h2f5d36b8;
    11'b01000100001: data <= 32'h35d1bcbf;
    11'b01000100010: data <= 32'ha744bd88;
    11'b01000100011: data <= 32'hbd4fbae9;
    11'b01000100100: data <= 32'hbf3fbbd8;
    11'b01000100101: data <= 32'hb56fbda6;
    11'b01000100110: data <= 32'h3de0bbb5;
    11'b01000100111: data <= 32'h3cdc32bb;
    11'b01000101000: data <= 32'hbad43ad5;
    11'b01000101001: data <= 32'hc05639f3;
    11'b01000101010: data <= 32'hbde43aff;
    11'b01000101011: data <= 32'hb4a33d8f;
    11'b01000101100: data <= 32'hb3e53c37;
    11'b01000101101: data <= 32'hb980b7ae;
    11'b01000101110: data <= 32'haf81bdb9;
    11'b01000101111: data <= 32'h3ce0b416;
    11'b01000110000: data <= 32'h3f353f2d;
    11'b01000110001: data <= 32'h3d17404e;
    11'b01000110010: data <= 32'h39a33830;
    11'b01000110011: data <= 32'h3869bac3;
    11'b01000110100: data <= 32'h2b66b888;
    11'b01000110101: data <= 32'hbb042970;
    11'b01000110110: data <= 32'hbb65b940;
    11'b01000110111: data <= 32'h3864bfe2;
    11'b01000111000: data <= 32'h3f88c018;
    11'b01000111001: data <= 32'h3cafb9db;
    11'b01000111010: data <= 32'hbaf6368a;
    11'b01000111011: data <= 32'hbf2438a2;
    11'b01000111100: data <= 32'hbb5e382d;
    11'b01000111101: data <= 32'hb2ad3969;
    11'b01000111110: data <= 32'hbc1434fc;
    11'b01000111111: data <= 32'hc007ba24;
    11'b01001000000: data <= 32'hbd20bcab;
    11'b01001000001: data <= 32'h396f30a9;
    11'b01001000010: data <= 32'h3eee3f80;
    11'b01001000011: data <= 32'h3cb23fd8;
    11'b01001000100: data <= 32'h34ea38e5;
    11'b01001000101: data <= 32'h2de3a450;
    11'b01001000110: data <= 32'h99a63a87;
    11'b01001000111: data <= 32'hb6083d0d;
    11'b01001001000: data <= 32'hb279b17f;
    11'b01001001001: data <= 32'h3c01c04c;
    11'b01001001010: data <= 32'h3fdec0ad;
    11'b01001001011: data <= 32'h3d45b9eb;
    11'b01001001100: data <= 32'hb1523861;
    11'b01001001101: data <= 32'hb88936a8;
    11'b01001001110: data <= 32'h318bb124;
    11'b01001001111: data <= 32'h2f22b3c9;
    11'b01001010000: data <= 32'hbe0ab57e;
    11'b01001010001: data <= 32'hc181bbb9;
    11'b01001010010: data <= 32'hbee1bcf1;
    11'b01001010011: data <= 32'h3852b494;
    11'b01001010100: data <= 32'h3dcf3bf6;
    11'b01001010101: data <= 32'h37313c96;
    11'b01001010110: data <= 32'hb9333825;
    11'b01001010111: data <= 32'hb8af3a0e;
    11'b01001011000: data <= 32'hb05e3fbf;
    11'b01001011001: data <= 32'hb3434023;
    11'b01001011010: data <= 32'hb44830dd;
    11'b01001011011: data <= 32'h3850bfa2;
    11'b01001011100: data <= 32'h3dfcbf13;
    11'b01001011101: data <= 32'h3dce2c90;
    11'b01001011110: data <= 32'h3a553c66;
    11'b01001011111: data <= 32'h3a3635d5;
    11'b01001100000: data <= 32'h3cc6b8f2;
    11'b01001100001: data <= 32'h37dfb8a6;
    11'b01001100010: data <= 32'hbdd4b482;
    11'b01001100011: data <= 32'hc10bba4e;
    11'b01001100100: data <= 32'hbce9be10;
    11'b01001100101: data <= 32'h3aecbd28;
    11'b01001100110: data <= 32'h3cc1b5ed;
    11'b01001100111: data <= 32'hb4dd2f5f;
    11'b01001101000: data <= 32'hbd683359;
    11'b01001101001: data <= 32'hbab73bf0;
    11'b01001101010: data <= 32'hafa6404d;
    11'b01001101011: data <= 32'hb7ee4001;
    11'b01001101100: data <= 32'hbc992e75;
    11'b01001101101: data <= 32'hb95bbdf2;
    11'b01001101110: data <= 32'h390dbabd;
    11'b01001101111: data <= 32'h3d883c06;
    11'b01001110000: data <= 32'h3d763e2a;
    11'b01001110001: data <= 32'h3dba35ae;
    11'b01001110010: data <= 32'h3e2db854;
    11'b01001110011: data <= 32'h397d2026;
    11'b01001110100: data <= 32'hbbd9391b;
    11'b01001110101: data <= 32'hbe6fb1e1;
    11'b01001110110: data <= 32'hb439bee1;
    11'b01001110111: data <= 32'h3d56c060;
    11'b01001111000: data <= 32'h3c41bd8a;
    11'b01001111001: data <= 32'hb85eb84b;
    11'b01001111010: data <= 32'hbcbcadfa;
    11'b01001111011: data <= 32'hb49a38c4;
    11'b01001111100: data <= 32'h332e3dbd;
    11'b01001111101: data <= 32'hbb4d3ce1;
    11'b01001111110: data <= 32'hc08eb378;
    11'b01001111111: data <= 32'hbfa3bcad;
    11'b01010000000: data <= 32'hb0e5b405;
    11'b01010000001: data <= 32'h3c6a3d26;
    11'b01010000010: data <= 32'h3ccc3d77;
    11'b01010000011: data <= 32'h3c38329d;
    11'b01010000100: data <= 32'h3c59ab94;
    11'b01010000101: data <= 32'h38ca3cbd;
    11'b01010000110: data <= 32'hb7203fbd;
    11'b01010000111: data <= 32'hb9d93898;
    11'b01010001000: data <= 32'h35ffbe91;
    11'b01010001001: data <= 32'h3dd2c0c6;
    11'b01010001010: data <= 32'h3c06bdbc;
    11'b01010001011: data <= 32'hb17ab72f;
    11'b01010001100: data <= 32'hb18db434;
    11'b01010001101: data <= 32'h3b08af43;
    11'b01010001110: data <= 32'h3ab03649;
    11'b01010001111: data <= 32'hbc733655;
    11'b01010010000: data <= 32'hc1cdb7c9;
    11'b01010010001: data <= 32'hc0d0bc46;
    11'b01010010010: data <= 32'hb64fb609;
    11'b01010010011: data <= 32'h3a3238f3;
    11'b01010010100: data <= 32'h372537d3;
    11'b01010010101: data <= 32'h1ec2b1f0;
    11'b01010010110: data <= 32'h343d3663;
    11'b01010010111: data <= 32'h365f405a;
    11'b01010011000: data <= 32'hb14241a3;
    11'b01010011001: data <= 32'hb8233c33;
    11'b01010011010: data <= 32'h3019bd38;
    11'b01010011011: data <= 32'h3b85bf1f;
    11'b01010011100: data <= 32'h3ac5b87c;
    11'b01010011101: data <= 32'h374e32eb;
    11'b01010011110: data <= 32'h3c1cb3eb;
    11'b01010011111: data <= 32'h3ffbb95d;
    11'b01010100000: data <= 32'h3dabb243;
    11'b01010100001: data <= 32'hbb5333b4;
    11'b01010100010: data <= 32'hc13eb4a5;
    11'b01010100011: data <= 32'hbf88bc4b;
    11'b01010100100: data <= 32'h1c2ebc2d;
    11'b01010100101: data <= 32'h3885b8bf;
    11'b01010100110: data <= 32'hb624b936;
    11'b01010100111: data <= 32'hbb56b9bd;
    11'b01010101000: data <= 32'hb2843725;
    11'b01010101001: data <= 32'h368240a8;
    11'b01010101010: data <= 32'hb1ee4181;
    11'b01010101011: data <= 32'hbc433bc8;
    11'b01010101100: data <= 32'hbb52bb51;
    11'b01010101101: data <= 32'ha8a8ba52;
    11'b01010101110: data <= 32'h3805388c;
    11'b01010101111: data <= 32'h3a6a3aec;
    11'b01010110000: data <= 32'h3e73b32c;
    11'b01010110001: data <= 32'h40c2ba79;
    11'b01010110010: data <= 32'h3e8d2c90;
    11'b01010110011: data <= 32'hb7063bdb;
    11'b01010110100: data <= 32'hbe9c36ae;
    11'b01010110101: data <= 32'hba04bbde;
    11'b01010110110: data <= 32'h3959beba;
    11'b01010110111: data <= 32'h37dbbe1c;
    11'b01010111000: data <= 32'hba7cbd7b;
    11'b01010111001: data <= 32'hbc3abc7f;
    11'b01010111010: data <= 32'h310321ab;
    11'b01010111011: data <= 32'h3ab13e40;
    11'b01010111100: data <= 32'hb4dd3f55;
    11'b01010111101: data <= 32'hbfa2376a;
    11'b01010111110: data <= 32'hc021b943;
    11'b01010111111: data <= 32'hbb57a950;
    11'b01011000000: data <= 32'h2d353c93;
    11'b01011000001: data <= 32'h38703b28;
    11'b01011000010: data <= 32'h3cc0b6f4;
    11'b01011000011: data <= 32'h3f4bb8f1;
    11'b01011000100: data <= 32'h3da03b98;
    11'b01011000101: data <= 32'h288a405a;
    11'b01011000110: data <= 32'hb9203d2c;
    11'b01011000111: data <= 32'h3156b9b2;
    11'b01011001000: data <= 32'h3c06bf06;
    11'b01011001001: data <= 32'h365fbe1d;
    11'b01011001010: data <= 32'hb9b0bce7;
    11'b01011001011: data <= 32'hb5a8bcc7;
    11'b01011001100: data <= 32'h3cd6b92e;
    11'b01011001101: data <= 32'h3e4f367d;
    11'b01011001110: data <= 32'hb45539f8;
    11'b01011001111: data <= 32'hc0bda40a;
    11'b01011010000: data <= 32'hc107b869;
    11'b01011010001: data <= 32'hbc952db4;
    11'b01011010010: data <= 32'hb27d3a4c;
    11'b01011010011: data <= 32'hb17430ad;
    11'b01011010100: data <= 32'h2937bbaa;
    11'b01011010101: data <= 32'h3a19b6b7;
    11'b01011010110: data <= 32'h3bd43efc;
    11'b01011010111: data <= 32'h34c04206;
    11'b01011011000: data <= 32'hb2203f32;
    11'b01011011001: data <= 32'h3390b5d0;
    11'b01011011010: data <= 32'h3920bc95;
    11'b01011011011: data <= 32'h2f68b88f;
    11'b01011011100: data <= 32'hb5c8b5a6;
    11'b01011011101: data <= 32'h3905bbb4;
    11'b01011011110: data <= 32'h408ebcaa;
    11'b01011011111: data <= 32'h4074b652;
    11'b01011100000: data <= 32'h9d0d345b;
    11'b01011100001: data <= 32'hc01b1d69;
    11'b01011100010: data <= 32'hbfa8b73b;
    11'b01011100011: data <= 32'hb89db4aa;
    11'b01011100100: data <= 32'hb30fb1d9;
    11'b01011100101: data <= 32'hbba4bb8c;
    11'b01011100110: data <= 32'hbc4bbe60;
    11'b01011100111: data <= 32'ha5c3b7ea;
    11'b01011101000: data <= 32'h3a4c3f52;
    11'b01011101001: data <= 32'h35a441c4;
    11'b01011101010: data <= 32'hb74a3e60;
    11'b01011101011: data <= 32'hb85ab01c;
    11'b01011101100: data <= 32'hb468b253;
    11'b01011101101: data <= 32'hb5b639dc;
    11'b01011101110: data <= 32'hb1ef38d6;
    11'b01011101111: data <= 32'h3c75b9c3;
    11'b01011110000: data <= 32'h413abd69;
    11'b01011110001: data <= 32'h40bdb679;
    11'b01011110010: data <= 32'h35c339da;
    11'b01011110011: data <= 32'hbc753913;
    11'b01011110100: data <= 32'hb902b30e;
    11'b01011110101: data <= 32'h3620b9c4;
    11'b01011110110: data <= 32'hac27bbee;
    11'b01011110111: data <= 32'hbd9ebe85;
    11'b01011111000: data <= 32'hbdeabfe5;
    11'b01011111001: data <= 32'h290fbaf4;
    11'b01011111010: data <= 32'h3c733c4f;
    11'b01011111011: data <= 32'h35fb3f4c;
    11'b01011111100: data <= 32'hbc3f3a7b;
    11'b01011111101: data <= 32'hbe29ae87;
    11'b01011111110: data <= 32'hbc8a3870;
    11'b01011111111: data <= 32'hba6c3e3f;
    11'b01100000000: data <= 32'hb6d53b93;
    11'b01100000001: data <= 32'h397aba63;
    11'b01100000010: data <= 32'h3fc3bd27;
    11'b01100000011: data <= 32'h3f953303;
    11'b01100000100: data <= 32'h38ea3efe;
    11'b01100000101: data <= 32'haf0e3df8;
    11'b01100000110: data <= 32'h384d2fa9;
    11'b01100000111: data <= 32'h3c2fb9f8;
    11'b01100001000: data <= 32'h1b8bbbbb;
    11'b01100001001: data <= 32'hbda8bd92;
    11'b01100001010: data <= 32'hbc29bf61;
    11'b01100001011: data <= 32'h3b1ebd52;
    11'b01100001100: data <= 32'h3f53ac2a;
    11'b01100001101: data <= 32'h38123806;
    11'b01100001110: data <= 32'hbdb29cc1;
    11'b01100001111: data <= 32'hbfc4b1e6;
    11'b01100010000: data <= 32'hbd303a33;
    11'b01100010001: data <= 32'hbb833de9;
    11'b01100010010: data <= 32'hbbec36d3;
    11'b01100010011: data <= 32'hb72abd26;
    11'b01100010100: data <= 32'h3948bcdb;
    11'b01100010101: data <= 32'h3c863b06;
    11'b01100010110: data <= 32'h39504107;
    11'b01100010111: data <= 32'h36883fd2;
    11'b01100011000: data <= 32'h3b153604;
    11'b01100011001: data <= 32'h3b7fb410;
    11'b01100011010: data <= 32'hb32ca421;
    11'b01100011011: data <= 32'hbccbb528;
    11'b01100011100: data <= 32'hb354bd27;
    11'b01100011101: data <= 32'h3f7bbe80;
    11'b01100011110: data <= 32'h40ebbb54;
    11'b01100011111: data <= 32'h39e2b40d;
    11'b01100100000: data <= 32'hbcb7b453;
    11'b01100100001: data <= 32'hbd5eb160;
    11'b01100100010: data <= 32'hb871383e;
    11'b01100100011: data <= 32'hb94539a5;
    11'b01100100100: data <= 32'hbe34b86f;
    11'b01100100101: data <= 32'hbe64bfac;
    11'b01100100110: data <= 32'hb686bd31;
    11'b01100100111: data <= 32'h38fe3be5;
    11'b01100101000: data <= 32'h38d440c0;
    11'b01100101001: data <= 32'h34603e6d;
    11'b01100101010: data <= 32'h35433598;
    11'b01100101011: data <= 32'h30f837c1;
    11'b01100101100: data <= 32'hb9983d41;
    11'b01100101101: data <= 32'hbc4c3b51;
    11'b01100101110: data <= 32'h33aeb9ad;
    11'b01100101111: data <= 32'h4061bea5;
    11'b01100110000: data <= 32'h40fcbc2c;
    11'b01100110001: data <= 32'h3b13a921;
    11'b01100110010: data <= 32'hb6cf3225;
    11'b01100110011: data <= 32'ha7a22bf3;
    11'b01100110100: data <= 32'h396831f5;
    11'b01100110101: data <= 32'hb0faa9b7;
    11'b01100110110: data <= 32'hbf4cbcdf;
    11'b01100110111: data <= 32'hc037c073;
    11'b01100111000: data <= 32'hb8e3be07;
    11'b01100111001: data <= 32'h39f9363f;
    11'b01100111010: data <= 32'h38da3d2f;
    11'b01100111011: data <= 32'hb3343887;
    11'b01100111100: data <= 32'hb892274d;
    11'b01100111101: data <= 32'hb95e3c2d;
    11'b01100111110: data <= 32'hbc6c4078;
    11'b01100111111: data <= 32'hbcd13e28;
    11'b01101000000: data <= 32'hac4ab85f;
    11'b01101000001: data <= 32'h3dfebe37;
    11'b01101000010: data <= 32'h3f22b84e;
    11'b01101000011: data <= 32'h3a6c3ac4;
    11'b01101000100: data <= 32'h360c3c00;
    11'b01101000101: data <= 32'h3ce1363c;
    11'b01101000110: data <= 32'h3e8c2e8a;
    11'b01101000111: data <= 32'h3217aed8;
    11'b01101001000: data <= 32'hbf0cbbc2;
    11'b01101001001: data <= 32'hbf2abf92;
    11'b01101001010: data <= 32'h2cecbea1;
    11'b01101001011: data <= 32'h3d91b86c;
    11'b01101001100: data <= 32'h39f5aeb2;
    11'b01101001101: data <= 32'hb8cbb877;
    11'b01101001110: data <= 32'hbc18b5d2;
    11'b01101001111: data <= 32'hba9f3ca7;
    11'b01101010000: data <= 32'hbc52408d;
    11'b01101010001: data <= 32'hbdf93cd9;
    11'b01101010010: data <= 32'hbc09bb74;
    11'b01101010011: data <= 32'h30b4bdf1;
    11'b01101010100: data <= 32'h39a52e1a;
    11'b01101010101: data <= 32'h38233e83;
    11'b01101010110: data <= 32'h3a273dd8;
    11'b01101010111: data <= 32'h3ec63837;
    11'b01101011000: data <= 32'h3f0335df;
    11'b01101011001: data <= 32'h2e85395b;
    11'b01101011010: data <= 32'hbe2f312f;
    11'b01101011011: data <= 32'hbc22bc20;
    11'b01101011100: data <= 32'h3c29be68;
    11'b01101011101: data <= 32'h4009bd04;
    11'b01101011110: data <= 32'h3b21bbe8;
    11'b01101011111: data <= 32'hb842bc56;
    11'b01101100000: data <= 32'hb899b83a;
    11'b01101100001: data <= 32'ha8be3b3c;
    11'b01101100010: data <= 32'hb81d3e52;
    11'b01101100011: data <= 32'hbed2347f;
    11'b01101100100: data <= 32'hbffbbe37;
    11'b01101100101: data <= 32'hbc31be17;
    11'b01101100110: data <= 32'hadf1355f;
    11'b01101100111: data <= 32'h33603e77;
    11'b01101101000: data <= 32'h38cd3c4f;
    11'b01101101001: data <= 32'h3cee33d2;
    11'b01101101010: data <= 32'h3c3b3a2b;
    11'b01101101011: data <= 32'hb5a33f51;
    11'b01101101100: data <= 32'hbd9a3e18;
    11'b01101101101: data <= 32'hb79bb05a;
    11'b01101101110: data <= 32'h3ddcbd7a;
    11'b01101101111: data <= 32'h400ebd4a;
    11'b01101110000: data <= 32'h3a90bb19;
    11'b01101110001: data <= 32'had9ab9fc;
    11'b01101110010: data <= 32'h388db57e;
    11'b01101110011: data <= 32'h3d413871;
    11'b01101110100: data <= 32'h351a3a3d;
    11'b01101110101: data <= 32'hbeb4b772;
    11'b01101110110: data <= 32'hc0d7bf6d;
    11'b01101110111: data <= 32'hbd82be36;
    11'b01101111000: data <= 32'hb08b23af;
    11'b01101111001: data <= 32'h30e63996;
    11'b01101111010: data <= 32'h2e81accc;
    11'b01101111011: data <= 32'h3515b68e;
    11'b01101111100: data <= 32'h318f3c06;
    11'b01101111101: data <= 32'hba26414c;
    11'b01101111110: data <= 32'hbd944092;
    11'b01101111111: data <= 32'hb85833c3;
    11'b01110000000: data <= 32'h3b6ebc8e;
    11'b01110000001: data <= 32'h3ce4ba7f;
    11'b01110000010: data <= 32'h36a0a4fb;
    11'b01110000011: data <= 32'h361d2d78;
    11'b01110000100: data <= 32'h3ed00a80;
    11'b01110000101: data <= 32'h40d93605;
    11'b01110000110: data <= 32'h3b5f3822;
    11'b01110000111: data <= 32'hbdc8b5d9;
    11'b01110001000: data <= 32'hc02cbdcc;
    11'b01110001001: data <= 32'hb9e1bd98;
    11'b01110001010: data <= 32'h37dfb8c2;
    11'b01110001011: data <= 32'h34d0b8a3;
    11'b01110001100: data <= 32'hb55bbd6f;
    11'b01110001101: data <= 32'hb4babc62;
    11'b01110001110: data <= 32'hafe03b52;
    11'b01110001111: data <= 32'hb98d4150;
    11'b01110010000: data <= 32'hbda4400f;
    11'b01110010001: data <= 32'hbca5adc2;
    11'b01110010010: data <= 32'hb4b5bc40;
    11'b01110010011: data <= 32'ha4beb06f;
    11'b01110010100: data <= 32'hb23c3b19;
    11'b01110010101: data <= 32'h38343967;
    11'b01110010110: data <= 32'h40442f4b;
    11'b01110010111: data <= 32'h41483684;
    11'b01110011000: data <= 32'h3b763beb;
    11'b01110011001: data <= 32'hbcc7390d;
    11'b01110011010: data <= 32'hbd34b6dd;
    11'b01110011011: data <= 32'h3518bc02;
    11'b01110011100: data <= 32'h3cebbc12;
    11'b01110011101: data <= 32'h3721bda3;
    11'b01110011110: data <= 32'hb75bc006;
    11'b01110011111: data <= 32'hb000bda4;
    11'b01110100000: data <= 32'h383838b3;
    11'b01110100001: data <= 32'h23f23fc2;
    11'b01110100010: data <= 32'hbd1d3c2a;
    11'b01110100011: data <= 32'hbf64ba6b;
    11'b01110100100: data <= 32'hbdb3bc72;
    11'b01110100101: data <= 32'hbbc83418;
    11'b01110100110: data <= 32'hb97a3c80;
    11'b01110100111: data <= 32'h33f136f4;
    11'b01110101000: data <= 32'h3e9cb49d;
    11'b01110101001: data <= 32'h3fae37ad;
    11'b01110101010: data <= 32'h36aa3f5b;
    11'b01110101011: data <= 32'hbc433fad;
    11'b01110101100: data <= 32'hb8f93923;
    11'b01110101101: data <= 32'h3bbdb823;
    11'b01110101110: data <= 32'h3d8dbb7c;
    11'b01110101111: data <= 32'h3483bd28;
    11'b01110110000: data <= 32'hb52fbec4;
    11'b01110110001: data <= 32'h39acbccf;
    11'b01110110010: data <= 32'h3f2f3402;
    11'b01110110011: data <= 32'h3c253c2d;
    11'b01110110100: data <= 32'hbba72e34;
    11'b01110110101: data <= 32'hc02bbd05;
    11'b01110110110: data <= 32'hbeeebc50;
    11'b01110110111: data <= 32'hbc4f32e6;
    11'b01110111000: data <= 32'hba4d3815;
    11'b01110111001: data <= 32'hb412b903;
    11'b01110111010: data <= 32'h3952bc87;
    11'b01110111011: data <= 32'h3aef3657;
    11'b01110111100: data <= 32'hb0c340e0;
    11'b01110111101: data <= 32'hbc1a4151;
    11'b01110111110: data <= 32'hb70b3c77;
    11'b01110111111: data <= 32'h39ccb291;
    11'b01111000000: data <= 32'h3979b64f;
    11'b01111000001: data <= 32'hb4eab5d4;
    11'b01111000010: data <= 32'hb1fcb9c6;
    11'b01111000011: data <= 32'h3e65b9c1;
    11'b01111000100: data <= 32'h41c32bd1;
    11'b01111000101: data <= 32'h3f163885;
    11'b01111000110: data <= 32'hb8b5ad91;
    11'b01111000111: data <= 32'hbebdbbb8;
    11'b01111001000: data <= 32'hbc2fba0f;
    11'b01111001001: data <= 32'hb585ab7f;
    11'b01111001010: data <= 32'hb82eb80d;
    11'b01111001011: data <= 32'hb97dbf89;
    11'b01111001100: data <= 32'hb03cbfef;
    11'b01111001101: data <= 32'h34c92f5e;
    11'b01111001110: data <= 32'hb2b340b1;
    11'b01111001111: data <= 32'hbb3640bc;
    11'b01111010000: data <= 32'hb9d839d3;
    11'b01111010001: data <= 32'hb337b2cb;
    11'b01111010010: data <= 32'hb838345a;
    11'b01111010011: data <= 32'hbc6e3997;
    11'b01111010100: data <= 32'hb4792fd7;
    11'b01111010101: data <= 32'h3f98b744;
    11'b01111010110: data <= 32'h4226a3c1;
    11'b01111010111: data <= 32'h3f1739ce;
    11'b01111011000: data <= 32'hb60d3907;
    11'b01111011001: data <= 32'hbb3023ae;
    11'b01111011010: data <= 32'h307eb0ef;
    11'b01111011011: data <= 32'h3902b2a8;
    11'b01111011100: data <= 32'hb2f4bcb6;
    11'b01111011101: data <= 32'hbb17c10e;
    11'b01111011110: data <= 32'hb405c0ac;
    11'b01111011111: data <= 32'h394db31a;
    11'b01111100000: data <= 32'h37123e72;
    11'b01111100001: data <= 32'hb87c3d10;
    11'b01111100010: data <= 32'hbc76b225;
    11'b01111100011: data <= 32'hbcb2b6be;
    11'b01111100100: data <= 32'hbdee39ba;
    11'b01111100101: data <= 32'hbebf3ccf;
    11'b01111100110: data <= 32'hb8f5317d;
    11'b01111100111: data <= 32'h3d86ba35;
    11'b01111101000: data <= 32'h4085b074;
    11'b01111101001: data <= 32'h3c533d09;
    11'b01111101010: data <= 32'hb6623ed9;
    11'b01111101011: data <= 32'hb1fd3c61;
    11'b01111101100: data <= 32'h3c203775;
    11'b01111101101: data <= 32'h3c4c9fa6;
    11'b01111101110: data <= 32'hb46dbbff;
    11'b01111101111: data <= 32'hbb68c046;
    11'b01111110000: data <= 32'h3437bffb;
    11'b01111110001: data <= 32'h3ed5b6e2;
    11'b01111110010: data <= 32'h3de3398f;
    11'b01111110011: data <= 32'hac462e4c;
    11'b01111110100: data <= 32'hbcbabb77;
    11'b01111110101: data <= 32'hbd9ab81f;
    11'b01111110110: data <= 32'hbe2d3a9a;
    11'b01111110111: data <= 32'hbed23b38;
    11'b01111111000: data <= 32'hbc1bb937;
    11'b01111111001: data <= 32'h3603be7d;
    11'b01111111010: data <= 32'h3c06b6b4;
    11'b01111111011: data <= 32'h33723e93;
    11'b01111111100: data <= 32'hb80b40b1;
    11'b01111111101: data <= 32'h2f913e34;
    11'b01111111110: data <= 32'h3c643a01;
    11'b01111111111: data <= 32'h38fe37b7;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    