module pin_update_vmm_input(
output_real_0_0, output_imag_0_0,
output_real_1_0, output_imag_1_0,
output_real_2_0, output_imag_2_0,
output_real_3_0, output_imag_3_0,
output_real_4_0, output_imag_4_0,
output_real_5_0, output_imag_5_0,
output_real_6_0, output_imag_6_0,
output_real_7_0, output_imag_7_0,
output_real_8_0, output_imag_8_0,
output_real_9_0, output_imag_9_0,
output_real_10_0, output_imag_10_0,
output_real_11_0, output_imag_11_0,
output_real_12_0, output_imag_12_0,
output_real_13_0, output_imag_13_0,
output_real_14_0, output_imag_14_0,
output_real_15_0, output_imag_15_0,
output_real_16_0, output_imag_16_0,
output_real_17_0, output_imag_17_0,
output_real_18_0, output_imag_18_0,
output_real_19_0, output_imag_19_0,
output_real_20_0, output_imag_20_0,
output_real_21_0, output_imag_21_0,
output_real_22_0, output_imag_22_0,
output_real_23_0, output_imag_23_0,
output_real_24_0, output_imag_24_0,
output_real_25_0, output_imag_25_0,
output_real_26_0, output_imag_26_0,
output_real_27_0, output_imag_27_0,
output_real_28_0, output_imag_28_0,
output_real_29_0, output_imag_29_0,
output_real_30_0, output_imag_30_0,
output_real_31_0, output_imag_31_0,
output_real_32_0, output_imag_32_0,
output_real_33_0, output_imag_33_0,
output_real_34_0, output_imag_34_0,
output_real_35_0, output_imag_35_0,
output_real_36_0, output_imag_36_0,
output_real_37_0, output_imag_37_0,
output_real_38_0, output_imag_38_0,
output_real_39_0, output_imag_39_0,
output_real_40_0, output_imag_40_0,
output_real_41_0, output_imag_41_0,
output_real_42_0, output_imag_42_0,
output_real_43_0, output_imag_43_0,
output_real_44_0, output_imag_44_0,
output_real_45_0, output_imag_45_0,
output_real_46_0, output_imag_46_0,
output_real_47_0, output_imag_47_0,
output_real_48_0, output_imag_48_0,
output_real_49_0, output_imag_49_0,
output_real_50_0, output_imag_50_0,
output_real_51_0, output_imag_51_0,
output_real_52_0, output_imag_52_0,
output_real_53_0, output_imag_53_0,
output_real_54_0, output_imag_54_0,
output_real_55_0, output_imag_55_0,
output_real_56_0, output_imag_56_0,
output_real_57_0, output_imag_57_0,
output_real_58_0, output_imag_58_0,
output_real_59_0, output_imag_59_0,
output_real_60_0, output_imag_60_0,
output_real_61_0, output_imag_61_0,
output_real_62_0, output_imag_62_0,
output_real_63_0, output_imag_63_0,

output_real_0_1, output_imag_0_1,
output_real_1_1, output_imag_1_1,
output_real_2_1, output_imag_2_1,
output_real_3_1, output_imag_3_1,
output_real_4_1, output_imag_4_1,
output_real_5_1, output_imag_5_1,
output_real_6_1, output_imag_6_1,
output_real_7_1, output_imag_7_1,
output_real_8_1, output_imag_8_1,
output_real_9_1, output_imag_9_1,
output_real_10_1, output_imag_10_1,
output_real_11_1, output_imag_11_1,
output_real_12_1, output_imag_12_1,
output_real_13_1, output_imag_13_1,
output_real_14_1, output_imag_14_1,
output_real_15_1, output_imag_15_1,
output_real_16_1, output_imag_16_1,
output_real_17_1, output_imag_17_1,
output_real_18_1, output_imag_18_1,
output_real_19_1, output_imag_19_1,
output_real_20_1, output_imag_20_1,
output_real_21_1, output_imag_21_1,
output_real_22_1, output_imag_22_1,
output_real_23_1, output_imag_23_1,
output_real_24_1, output_imag_24_1,
output_real_25_1, output_imag_25_1,
output_real_26_1, output_imag_26_1,
output_real_27_1, output_imag_27_1,
output_real_28_1, output_imag_28_1,
output_real_29_1, output_imag_29_1,
output_real_30_1, output_imag_30_1,
output_real_31_1, output_imag_31_1,
output_real_32_1, output_imag_32_1,
output_real_33_1, output_imag_33_1,
output_real_34_1, output_imag_34_1,
output_real_35_1, output_imag_35_1,
output_real_36_1, output_imag_36_1,
output_real_37_1, output_imag_37_1,
output_real_38_1, output_imag_38_1,
output_real_39_1, output_imag_39_1,
output_real_40_1, output_imag_40_1,
output_real_41_1, output_imag_41_1,
output_real_42_1, output_imag_42_1,
output_real_43_1, output_imag_43_1,
output_real_44_1, output_imag_44_1,
output_real_45_1, output_imag_45_1,
output_real_46_1, output_imag_46_1,
output_real_47_1, output_imag_47_1,
output_real_48_1, output_imag_48_1,
output_real_49_1, output_imag_49_1,
output_real_50_1, output_imag_50_1,
output_real_51_1, output_imag_51_1,
output_real_52_1, output_imag_52_1,
output_real_53_1, output_imag_53_1,
output_real_54_1, output_imag_54_1,
output_real_55_1, output_imag_55_1,
output_real_56_1, output_imag_56_1,
output_real_57_1, output_imag_57_1,
output_real_58_1, output_imag_58_1,
output_real_59_1, output_imag_59_1,
output_real_60_1, output_imag_60_1,
output_real_61_1, output_imag_61_1,
output_real_62_1, output_imag_62_1,
output_real_63_1, output_imag_63_1,

output_real_0_2, output_imag_0_2,
output_real_1_2, output_imag_1_2,
output_real_2_2, output_imag_2_2,
output_real_3_2, output_imag_3_2,
output_real_4_2, output_imag_4_2,
output_real_5_2, output_imag_5_2,
output_real_6_2, output_imag_6_2,
output_real_7_2, output_imag_7_2,
output_real_8_2, output_imag_8_2,
output_real_9_2, output_imag_9_2,
output_real_10_2, output_imag_10_2,
output_real_11_2, output_imag_11_2,
output_real_12_2, output_imag_12_2,
output_real_13_2, output_imag_13_2,
output_real_14_2, output_imag_14_2,
output_real_15_2, output_imag_15_2,
output_real_16_2, output_imag_16_2,
output_real_17_2, output_imag_17_2,
output_real_18_2, output_imag_18_2,
output_real_19_2, output_imag_19_2,
output_real_20_2, output_imag_20_2,
output_real_21_2, output_imag_21_2,
output_real_22_2, output_imag_22_2,
output_real_23_2, output_imag_23_2,
output_real_24_2, output_imag_24_2,
output_real_25_2, output_imag_25_2,
output_real_26_2, output_imag_26_2,
output_real_27_2, output_imag_27_2,
output_real_28_2, output_imag_28_2,
output_real_29_2, output_imag_29_2,
output_real_30_2, output_imag_30_2,
output_real_31_2, output_imag_31_2,
output_real_32_2, output_imag_32_2,
output_real_33_2, output_imag_33_2,
output_real_34_2, output_imag_34_2,
output_real_35_2, output_imag_35_2,
output_real_36_2, output_imag_36_2,
output_real_37_2, output_imag_37_2,
output_real_38_2, output_imag_38_2,
output_real_39_2, output_imag_39_2,
output_real_40_2, output_imag_40_2,
output_real_41_2, output_imag_41_2,
output_real_42_2, output_imag_42_2,
output_real_43_2, output_imag_43_2,
output_real_44_2, output_imag_44_2,
output_real_45_2, output_imag_45_2,
output_real_46_2, output_imag_46_2,
output_real_47_2, output_imag_47_2,
output_real_48_2, output_imag_48_2,
output_real_49_2, output_imag_49_2,
output_real_50_2, output_imag_50_2,
output_real_51_2, output_imag_51_2,
output_real_52_2, output_imag_52_2,
output_real_53_2, output_imag_53_2,
output_real_54_2, output_imag_54_2,
output_real_55_2, output_imag_55_2,
output_real_56_2, output_imag_56_2,
output_real_57_2, output_imag_57_2,
output_real_58_2, output_imag_58_2,
output_real_59_2, output_imag_59_2,
output_real_60_2, output_imag_60_2,
output_real_61_2, output_imag_61_2,
output_real_62_2, output_imag_62_2,
output_real_63_2, output_imag_63_2,

output_real_0_3, output_imag_0_3,
output_real_1_3, output_imag_1_3,
output_real_2_3, output_imag_2_3,
output_real_3_3, output_imag_3_3,
output_real_4_3, output_imag_4_3,
output_real_5_3, output_imag_5_3,
output_real_6_3, output_imag_6_3,
output_real_7_3, output_imag_7_3,
output_real_8_3, output_imag_8_3,
output_real_9_3, output_imag_9_3,
output_real_10_3, output_imag_10_3,
output_real_11_3, output_imag_11_3,
output_real_12_3, output_imag_12_3,
output_real_13_3, output_imag_13_3,
output_real_14_3, output_imag_14_3,
output_real_15_3, output_imag_15_3,
output_real_16_3, output_imag_16_3,
output_real_17_3, output_imag_17_3,
output_real_18_3, output_imag_18_3,
output_real_19_3, output_imag_19_3,
output_real_20_3, output_imag_20_3,
output_real_21_3, output_imag_21_3,
output_real_22_3, output_imag_22_3,
output_real_23_3, output_imag_23_3,
output_real_24_3, output_imag_24_3,
output_real_25_3, output_imag_25_3,
output_real_26_3, output_imag_26_3,
output_real_27_3, output_imag_27_3,
output_real_28_3, output_imag_28_3,
output_real_29_3, output_imag_29_3,
output_real_30_3, output_imag_30_3,
output_real_31_3, output_imag_31_3,
output_real_32_3, output_imag_32_3,
output_real_33_3, output_imag_33_3,
output_real_34_3, output_imag_34_3,
output_real_35_3, output_imag_35_3,
output_real_36_3, output_imag_36_3,
output_real_37_3, output_imag_37_3,
output_real_38_3, output_imag_38_3,
output_real_39_3, output_imag_39_3,
output_real_40_3, output_imag_40_3,
output_real_41_3, output_imag_41_3,
output_real_42_3, output_imag_42_3,
output_real_43_3, output_imag_43_3,
output_real_44_3, output_imag_44_3,
output_real_45_3, output_imag_45_3,
output_real_46_3, output_imag_46_3,
output_real_47_3, output_imag_47_3,
output_real_48_3, output_imag_48_3,
output_real_49_3, output_imag_49_3,
output_real_50_3, output_imag_50_3,
output_real_51_3, output_imag_51_3,
output_real_52_3, output_imag_52_3,
output_real_53_3, output_imag_53_3,
output_real_54_3, output_imag_54_3,
output_real_55_3, output_imag_55_3,
output_real_56_3, output_imag_56_3,
output_real_57_3, output_imag_57_3,
output_real_58_3, output_imag_58_3,
output_real_59_3, output_imag_59_3,
output_real_60_3, output_imag_60_3,
output_real_61_3, output_imag_61_3,
output_real_62_3, output_imag_62_3,
output_real_63_3, output_imag_63_3,

ssb,sdi,vmm_load,CLK,rst
);
input ssb,CLK;
input [27:0] sdi;
input vmm_load;
input rst;
reg [27:0] config0_0;
reg [27:0] config1_0;
reg [27:0] config2_0;
reg [27:0] config3_0;
reg [27:0] config4_0;
reg [27:0] config5_0;
reg [27:0] config6_0;
reg [27:0] config7_0;
reg [27:0] config8_0;
reg [27:0] config9_0;
reg [27:0] config10_0;
reg [27:0] config11_0;
reg [27:0] config12_0;
reg [27:0] config13_0;
reg [27:0] config14_0;
reg [27:0] config15_0;
reg [27:0] config16_0;
reg [27:0] config17_0;
reg [27:0] config18_0;
reg [27:0] config19_0;
reg [27:0] config20_0;
reg [27:0] config21_0;
reg [27:0] config22_0;
reg [27:0] config23_0;
reg [27:0] config24_0;
reg [27:0] config25_0;
reg [27:0] config26_0;
reg [27:0] config27_0;
reg [27:0] config28_0;
reg [27:0] config29_0;
reg [27:0] config30_0;
reg [27:0] config31_0;
reg [27:0] config32_0;
reg [27:0] config33_0;
reg [27:0] config34_0;
reg [27:0] config35_0;
reg [27:0] config36_0;
reg [27:0] config37_0;
reg [27:0] config38_0;
reg [27:0] config39_0;
reg [27:0] config40_0;
reg [27:0] config41_0;
reg [27:0] config42_0;
reg [27:0] config43_0;
reg [27:0] config44_0;
reg [27:0] config45_0;
reg [27:0] config46_0;
reg [27:0] config47_0;
reg [27:0] config48_0;
reg [27:0] config49_0;
reg [27:0] config50_0;
reg [27:0] config51_0;
reg [27:0] config52_0;
reg [27:0] config53_0;
reg [27:0] config54_0;
reg [27:0] config55_0;
reg [27:0] config56_0;
reg [27:0] config57_0;
reg [27:0] config58_0;
reg [27:0] config59_0;
reg [27:0] config60_0;
reg [27:0] config61_0;
reg [27:0] config62_0;
reg [27:0] config63_0;

reg [27:0] config0_1;
reg [27:0] config1_1;
reg [27:0] config2_1;
reg [27:0] config3_1;
reg [27:0] config4_1;
reg [27:0] config5_1;
reg [27:0] config6_1;
reg [27:0] config7_1;
reg [27:0] config8_1;
reg [27:0] config9_1;
reg [27:0] config10_1;
reg [27:0] config11_1;
reg [27:0] config12_1;
reg [27:0] config13_1;
reg [27:0] config14_1;
reg [27:0] config15_1;
reg [27:0] config16_1;
reg [27:0] config17_1;
reg [27:0] config18_1;
reg [27:0] config19_1;
reg [27:0] config20_1;
reg [27:0] config21_1;
reg [27:0] config22_1;
reg [27:0] config23_1;
reg [27:0] config24_1;
reg [27:0] config25_1;
reg [27:0] config26_1;
reg [27:0] config27_1;
reg [27:0] config28_1;
reg [27:0] config29_1;
reg [27:0] config30_1;
reg [27:0] config31_1;
reg [27:0] config32_1;
reg [27:0] config33_1;
reg [27:0] config34_1;
reg [27:0] config35_1;
reg [27:0] config36_1;
reg [27:0] config37_1;
reg [27:0] config38_1;
reg [27:0] config39_1;
reg [27:0] config40_1;
reg [27:0] config41_1;
reg [27:0] config42_1;
reg [27:0] config43_1;
reg [27:0] config44_1;
reg [27:0] config45_1;
reg [27:0] config46_1;
reg [27:0] config47_1;
reg [27:0] config48_1;
reg [27:0] config49_1;
reg [27:0] config50_1;
reg [27:0] config51_1;
reg [27:0] config52_1;
reg [27:0] config53_1;
reg [27:0] config54_1;
reg [27:0] config55_1;
reg [27:0] config56_1;
reg [27:0] config57_1;
reg [27:0] config58_1;
reg [27:0] config59_1;
reg [27:0] config60_1;
reg [27:0] config61_1;
reg [27:0] config62_1;
reg [27:0] config63_1;

reg [27:0] config0_2;
reg [27:0] config1_2;
reg [27:0] config2_2;
reg [27:0] config3_2;
reg [27:0] config4_2;
reg [27:0] config5_2;
reg [27:0] config6_2;
reg [27:0] config7_2;
reg [27:0] config8_2;
reg [27:0] config9_2;
reg [27:0] config10_2;
reg [27:0] config11_2;
reg [27:0] config12_2;
reg [27:0] config13_2;
reg [27:0] config14_2;
reg [27:0] config15_2;
reg [27:0] config16_2;
reg [27:0] config17_2;
reg [27:0] config18_2;
reg [27:0] config19_2;
reg [27:0] config20_2;
reg [27:0] config21_2;
reg [27:0] config22_2;
reg [27:0] config23_2;
reg [27:0] config24_2;
reg [27:0] config25_2;
reg [27:0] config26_2;
reg [27:0] config27_2;
reg [27:0] config28_2;
reg [27:0] config29_2;
reg [27:0] config30_2;
reg [27:0] config31_2;
reg [27:0] config32_2;
reg [27:0] config33_2;
reg [27:0] config34_2;
reg [27:0] config35_2;
reg [27:0] config36_2;
reg [27:0] config37_2;
reg [27:0] config38_2;
reg [27:0] config39_2;
reg [27:0] config40_2;
reg [27:0] config41_2;
reg [27:0] config42_2;
reg [27:0] config43_2;
reg [27:0] config44_2;
reg [27:0] config45_2;
reg [27:0] config46_2;
reg [27:0] config47_2;
reg [27:0] config48_2;
reg [27:0] config49_2;
reg [27:0] config50_2;
reg [27:0] config51_2;
reg [27:0] config52_2;
reg [27:0] config53_2;
reg [27:0] config54_2;
reg [27:0] config55_2;
reg [27:0] config56_2;
reg [27:0] config57_2;
reg [27:0] config58_2;
reg [27:0] config59_2;
reg [27:0] config60_2;
reg [27:0] config61_2;
reg [27:0] config62_2;
reg [27:0] config63_2;

reg [27:0] config0_3;
reg [27:0] config1_3;
reg [27:0] config2_3;
reg [27:0] config3_3;
reg [27:0] config4_3;
reg [27:0] config5_3;
reg [27:0] config6_3;
reg [27:0] config7_3;
reg [27:0] config8_3;
reg [27:0] config9_3;
reg [27:0] config10_3;
reg [27:0] config11_3;
reg [27:0] config12_3;
reg [27:0] config13_3;
reg [27:0] config14_3;
reg [27:0] config15_3;
reg [27:0] config16_3;
reg [27:0] config17_3;
reg [27:0] config18_3;
reg [27:0] config19_3;
reg [27:0] config20_3;
reg [27:0] config21_3;
reg [27:0] config22_3;
reg [27:0] config23_3;
reg [27:0] config24_3;
reg [27:0] config25_3;
reg [27:0] config26_3;
reg [27:0] config27_3;
reg [27:0] config28_3;
reg [27:0] config29_3;
reg [27:0] config30_3;
reg [27:0] config31_3;
reg [27:0] config32_3;
reg [27:0] config33_3;
reg [27:0] config34_3;
reg [27:0] config35_3;
reg [27:0] config36_3;
reg [27:0] config37_3;
reg [27:0] config38_3;
reg [27:0] config39_3;
reg [27:0] config40_3;
reg [27:0] config41_3;
reg [27:0] config42_3;
reg [27:0] config43_3;
reg [27:0] config44_3;
reg [27:0] config45_3;
reg [27:0] config46_3;
reg [27:0] config47_3;
reg [27:0] config48_3;
reg [27:0] config49_3;
reg [27:0] config50_3;
reg [27:0] config51_3;
reg [27:0] config52_3;
reg [27:0] config53_3;
reg [27:0] config54_3;
reg [27:0] config55_3;
reg [27:0] config56_3;
reg [27:0] config57_3;
reg [27:0] config58_3;
reg [27:0] config59_3;
reg [27:0] config60_3;
reg [27:0] config61_3;
reg [27:0] config62_3;
reg [27:0] config63_3;

output [9:0] output_real_0_0;
output [9:0] output_imag_0_0;
output [9:0] output_real_1_0;
output [9:0] output_imag_1_0;
output [9:0] output_real_2_0;
output [9:0] output_imag_2_0;
output [9:0] output_real_3_0;
output [9:0] output_imag_3_0;
output [9:0] output_real_4_0;
output [9:0] output_imag_4_0;
output [9:0] output_real_5_0;
output [9:0] output_imag_5_0;
output [9:0] output_real_6_0;
output [9:0] output_imag_6_0;
output [9:0] output_real_7_0;
output [9:0] output_imag_7_0;
output [9:0] output_real_8_0;
output [9:0] output_imag_8_0;
output [9:0] output_real_9_0;
output [9:0] output_imag_9_0;
output [9:0] output_real_10_0;
output [9:0] output_imag_10_0;
output [9:0] output_real_11_0;
output [9:0] output_imag_11_0;
output [9:0] output_real_12_0;
output [9:0] output_imag_12_0;
output [9:0] output_real_13_0;
output [9:0] output_imag_13_0;
output [9:0] output_real_14_0;
output [9:0] output_imag_14_0;
output [9:0] output_real_15_0;
output [9:0] output_imag_15_0;
output [9:0] output_real_16_0;
output [9:0] output_imag_16_0;
output [9:0] output_real_17_0;
output [9:0] output_imag_17_0;
output [9:0] output_real_18_0;
output [9:0] output_imag_18_0;
output [9:0] output_real_19_0;
output [9:0] output_imag_19_0;
output [9:0] output_real_20_0;
output [9:0] output_imag_20_0;
output [9:0] output_real_21_0;
output [9:0] output_imag_21_0;
output [9:0] output_real_22_0;
output [9:0] output_imag_22_0;
output [9:0] output_real_23_0;
output [9:0] output_imag_23_0;
output [9:0] output_real_24_0;
output [9:0] output_imag_24_0;
output [9:0] output_real_25_0;
output [9:0] output_imag_25_0;
output [9:0] output_real_26_0;
output [9:0] output_imag_26_0;
output [9:0] output_real_27_0;
output [9:0] output_imag_27_0;
output [9:0] output_real_28_0;
output [9:0] output_imag_28_0;
output [9:0] output_real_29_0;
output [9:0] output_imag_29_0;
output [9:0] output_real_30_0;
output [9:0] output_imag_30_0;
output [9:0] output_real_31_0;
output [9:0] output_imag_31_0;
output [9:0] output_real_32_0;
output [9:0] output_imag_32_0;
output [9:0] output_real_33_0;
output [9:0] output_imag_33_0;
output [9:0] output_real_34_0;
output [9:0] output_imag_34_0;
output [9:0] output_real_35_0;
output [9:0] output_imag_35_0;
output [9:0] output_real_36_0;
output [9:0] output_imag_36_0;
output [9:0] output_real_37_0;
output [9:0] output_imag_37_0;
output [9:0] output_real_38_0;
output [9:0] output_imag_38_0;
output [9:0] output_real_39_0;
output [9:0] output_imag_39_0;
output [9:0] output_real_40_0;
output [9:0] output_imag_40_0;
output [9:0] output_real_41_0;
output [9:0] output_imag_41_0;
output [9:0] output_real_42_0;
output [9:0] output_imag_42_0;
output [9:0] output_real_43_0;
output [9:0] output_imag_43_0;
output [9:0] output_real_44_0;
output [9:0] output_imag_44_0;
output [9:0] output_real_45_0;
output [9:0] output_imag_45_0;
output [9:0] output_real_46_0;
output [9:0] output_imag_46_0;
output [9:0] output_real_47_0;
output [9:0] output_imag_47_0;
output [9:0] output_real_48_0;
output [9:0] output_imag_48_0;
output [9:0] output_real_49_0;
output [9:0] output_imag_49_0;
output [9:0] output_real_50_0;
output [9:0] output_imag_50_0;
output [9:0] output_real_51_0;
output [9:0] output_imag_51_0;
output [9:0] output_real_52_0;
output [9:0] output_imag_52_0;
output [9:0] output_real_53_0;
output [9:0] output_imag_53_0;
output [9:0] output_real_54_0;
output [9:0] output_imag_54_0;
output [9:0] output_real_55_0;
output [9:0] output_imag_55_0;
output [9:0] output_real_56_0;
output [9:0] output_imag_56_0;
output [9:0] output_real_57_0;
output [9:0] output_imag_57_0;
output [9:0] output_real_58_0;
output [9:0] output_imag_58_0;
output [9:0] output_real_59_0;
output [9:0] output_imag_59_0;
output [9:0] output_real_60_0;
output [9:0] output_imag_60_0;
output [9:0] output_real_61_0;
output [9:0] output_imag_61_0;
output [9:0] output_real_62_0;
output [9:0] output_imag_62_0;
output [9:0] output_real_63_0;
output [9:0] output_imag_63_0;

output [9:0] output_real_0_1;
output [9:0] output_imag_0_1;
output [9:0] output_real_1_1;
output [9:0] output_imag_1_1;
output [9:0] output_real_2_1;
output [9:0] output_imag_2_1;
output [9:0] output_real_3_1;
output [9:0] output_imag_3_1;
output [9:0] output_real_4_1;
output [9:0] output_imag_4_1;
output [9:0] output_real_5_1;
output [9:0] output_imag_5_1;
output [9:0] output_real_6_1;
output [9:0] output_imag_6_1;
output [9:0] output_real_7_1;
output [9:0] output_imag_7_1;
output [9:0] output_real_8_1;
output [9:0] output_imag_8_1;
output [9:0] output_real_9_1;
output [9:0] output_imag_9_1;
output [9:0] output_real_10_1;
output [9:0] output_imag_10_1;
output [9:0] output_real_11_1;
output [9:0] output_imag_11_1;
output [9:0] output_real_12_1;
output [9:0] output_imag_12_1;
output [9:0] output_real_13_1;
output [9:0] output_imag_13_1;
output [9:0] output_real_14_1;
output [9:0] output_imag_14_1;
output [9:0] output_real_15_1;
output [9:0] output_imag_15_1;
output [9:0] output_real_16_1;
output [9:0] output_imag_16_1;
output [9:0] output_real_17_1;
output [9:0] output_imag_17_1;
output [9:0] output_real_18_1;
output [9:0] output_imag_18_1;
output [9:0] output_real_19_1;
output [9:0] output_imag_19_1;
output [9:0] output_real_20_1;
output [9:0] output_imag_20_1;
output [9:0] output_real_21_1;
output [9:0] output_imag_21_1;
output [9:0] output_real_22_1;
output [9:0] output_imag_22_1;
output [9:0] output_real_23_1;
output [9:0] output_imag_23_1;
output [9:0] output_real_24_1;
output [9:0] output_imag_24_1;
output [9:0] output_real_25_1;
output [9:0] output_imag_25_1;
output [9:0] output_real_26_1;
output [9:0] output_imag_26_1;
output [9:0] output_real_27_1;
output [9:0] output_imag_27_1;
output [9:0] output_real_28_1;
output [9:0] output_imag_28_1;
output [9:0] output_real_29_1;
output [9:0] output_imag_29_1;
output [9:0] output_real_30_1;
output [9:0] output_imag_30_1;
output [9:0] output_real_31_1;
output [9:0] output_imag_31_1;
output [9:0] output_real_32_1;
output [9:0] output_imag_32_1;
output [9:0] output_real_33_1;
output [9:0] output_imag_33_1;
output [9:0] output_real_34_1;
output [9:0] output_imag_34_1;
output [9:0] output_real_35_1;
output [9:0] output_imag_35_1;
output [9:0] output_real_36_1;
output [9:0] output_imag_36_1;
output [9:0] output_real_37_1;
output [9:0] output_imag_37_1;
output [9:0] output_real_38_1;
output [9:0] output_imag_38_1;
output [9:0] output_real_39_1;
output [9:0] output_imag_39_1;
output [9:0] output_real_40_1;
output [9:0] output_imag_40_1;
output [9:0] output_real_41_1;
output [9:0] output_imag_41_1;
output [9:0] output_real_42_1;
output [9:0] output_imag_42_1;
output [9:0] output_real_43_1;
output [9:0] output_imag_43_1;
output [9:0] output_real_44_1;
output [9:0] output_imag_44_1;
output [9:0] output_real_45_1;
output [9:0] output_imag_45_1;
output [9:0] output_real_46_1;
output [9:0] output_imag_46_1;
output [9:0] output_real_47_1;
output [9:0] output_imag_47_1;
output [9:0] output_real_48_1;
output [9:0] output_imag_48_1;
output [9:0] output_real_49_1;
output [9:0] output_imag_49_1;
output [9:0] output_real_50_1;
output [9:0] output_imag_50_1;
output [9:0] output_real_51_1;
output [9:0] output_imag_51_1;
output [9:0] output_real_52_1;
output [9:0] output_imag_52_1;
output [9:0] output_real_53_1;
output [9:0] output_imag_53_1;
output [9:0] output_real_54_1;
output [9:0] output_imag_54_1;
output [9:0] output_real_55_1;
output [9:0] output_imag_55_1;
output [9:0] output_real_56_1;
output [9:0] output_imag_56_1;
output [9:0] output_real_57_1;
output [9:0] output_imag_57_1;
output [9:0] output_real_58_1;
output [9:0] output_imag_58_1;
output [9:0] output_real_59_1;
output [9:0] output_imag_59_1;
output [9:0] output_real_60_1;
output [9:0] output_imag_60_1;
output [9:0] output_real_61_1;
output [9:0] output_imag_61_1;
output [9:0] output_real_62_1;
output [9:0] output_imag_62_1;
output [9:0] output_real_63_1;
output [9:0] output_imag_63_1;

output [9:0] output_real_0_2;
output [9:0] output_imag_0_2;
output [9:0] output_real_1_2;
output [9:0] output_imag_1_2;
output [9:0] output_real_2_2;
output [9:0] output_imag_2_2;
output [9:0] output_real_3_2;
output [9:0] output_imag_3_2;
output [9:0] output_real_4_2;
output [9:0] output_imag_4_2;
output [9:0] output_real_5_2;
output [9:0] output_imag_5_2;
output [9:0] output_real_6_2;
output [9:0] output_imag_6_2;
output [9:0] output_real_7_2;
output [9:0] output_imag_7_2;
output [9:0] output_real_8_2;
output [9:0] output_imag_8_2;
output [9:0] output_real_9_2;
output [9:0] output_imag_9_2;
output [9:0] output_real_10_2;
output [9:0] output_imag_10_2;
output [9:0] output_real_11_2;
output [9:0] output_imag_11_2;
output [9:0] output_real_12_2;
output [9:0] output_imag_12_2;
output [9:0] output_real_13_2;
output [9:0] output_imag_13_2;
output [9:0] output_real_14_2;
output [9:0] output_imag_14_2;
output [9:0] output_real_15_2;
output [9:0] output_imag_15_2;
output [9:0] output_real_16_2;
output [9:0] output_imag_16_2;
output [9:0] output_real_17_2;
output [9:0] output_imag_17_2;
output [9:0] output_real_18_2;
output [9:0] output_imag_18_2;
output [9:0] output_real_19_2;
output [9:0] output_imag_19_2;
output [9:0] output_real_20_2;
output [9:0] output_imag_20_2;
output [9:0] output_real_21_2;
output [9:0] output_imag_21_2;
output [9:0] output_real_22_2;
output [9:0] output_imag_22_2;
output [9:0] output_real_23_2;
output [9:0] output_imag_23_2;
output [9:0] output_real_24_2;
output [9:0] output_imag_24_2;
output [9:0] output_real_25_2;
output [9:0] output_imag_25_2;
output [9:0] output_real_26_2;
output [9:0] output_imag_26_2;
output [9:0] output_real_27_2;
output [9:0] output_imag_27_2;
output [9:0] output_real_28_2;
output [9:0] output_imag_28_2;
output [9:0] output_real_29_2;
output [9:0] output_imag_29_2;
output [9:0] output_real_30_2;
output [9:0] output_imag_30_2;
output [9:0] output_real_31_2;
output [9:0] output_imag_31_2;
output [9:0] output_real_32_2;
output [9:0] output_imag_32_2;
output [9:0] output_real_33_2;
output [9:0] output_imag_33_2;
output [9:0] output_real_34_2;
output [9:0] output_imag_34_2;
output [9:0] output_real_35_2;
output [9:0] output_imag_35_2;
output [9:0] output_real_36_2;
output [9:0] output_imag_36_2;
output [9:0] output_real_37_2;
output [9:0] output_imag_37_2;
output [9:0] output_real_38_2;
output [9:0] output_imag_38_2;
output [9:0] output_real_39_2;
output [9:0] output_imag_39_2;
output [9:0] output_real_40_2;
output [9:0] output_imag_40_2;
output [9:0] output_real_41_2;
output [9:0] output_imag_41_2;
output [9:0] output_real_42_2;
output [9:0] output_imag_42_2;
output [9:0] output_real_43_2;
output [9:0] output_imag_43_2;
output [9:0] output_real_44_2;
output [9:0] output_imag_44_2;
output [9:0] output_real_45_2;
output [9:0] output_imag_45_2;
output [9:0] output_real_46_2;
output [9:0] output_imag_46_2;
output [9:0] output_real_47_2;
output [9:0] output_imag_47_2;
output [9:0] output_real_48_2;
output [9:0] output_imag_48_2;
output [9:0] output_real_49_2;
output [9:0] output_imag_49_2;
output [9:0] output_real_50_2;
output [9:0] output_imag_50_2;
output [9:0] output_real_51_2;
output [9:0] output_imag_51_2;
output [9:0] output_real_52_2;
output [9:0] output_imag_52_2;
output [9:0] output_real_53_2;
output [9:0] output_imag_53_2;
output [9:0] output_real_54_2;
output [9:0] output_imag_54_2;
output [9:0] output_real_55_2;
output [9:0] output_imag_55_2;
output [9:0] output_real_56_2;
output [9:0] output_imag_56_2;
output [9:0] output_real_57_2;
output [9:0] output_imag_57_2;
output [9:0] output_real_58_2;
output [9:0] output_imag_58_2;
output [9:0] output_real_59_2;
output [9:0] output_imag_59_2;
output [9:0] output_real_60_2;
output [9:0] output_imag_60_2;
output [9:0] output_real_61_2;
output [9:0] output_imag_61_2;
output [9:0] output_real_62_2;
output [9:0] output_imag_62_2;
output [9:0] output_real_63_2;
output [9:0] output_imag_63_2;

output [9:0] output_real_0_3;
output [9:0] output_imag_0_3;
output [9:0] output_real_1_3;
output [9:0] output_imag_1_3;
output [9:0] output_real_2_3;
output [9:0] output_imag_2_3;
output [9:0] output_real_3_3;
output [9:0] output_imag_3_3;
output [9:0] output_real_4_3;
output [9:0] output_imag_4_3;
output [9:0] output_real_5_3;
output [9:0] output_imag_5_3;
output [9:0] output_real_6_3;
output [9:0] output_imag_6_3;
output [9:0] output_real_7_3;
output [9:0] output_imag_7_3;
output [9:0] output_real_8_3;
output [9:0] output_imag_8_3;
output [9:0] output_real_9_3;
output [9:0] output_imag_9_3;
output [9:0] output_real_10_3;
output [9:0] output_imag_10_3;
output [9:0] output_real_11_3;
output [9:0] output_imag_11_3;
output [9:0] output_real_12_3;
output [9:0] output_imag_12_3;
output [9:0] output_real_13_3;
output [9:0] output_imag_13_3;
output [9:0] output_real_14_3;
output [9:0] output_imag_14_3;
output [9:0] output_real_15_3;
output [9:0] output_imag_15_3;
output [9:0] output_real_16_3;
output [9:0] output_imag_16_3;
output [9:0] output_real_17_3;
output [9:0] output_imag_17_3;
output [9:0] output_real_18_3;
output [9:0] output_imag_18_3;
output [9:0] output_real_19_3;
output [9:0] output_imag_19_3;
output [9:0] output_real_20_3;
output [9:0] output_imag_20_3;
output [9:0] output_real_21_3;
output [9:0] output_imag_21_3;
output [9:0] output_real_22_3;
output [9:0] output_imag_22_3;
output [9:0] output_real_23_3;
output [9:0] output_imag_23_3;
output [9:0] output_real_24_3;
output [9:0] output_imag_24_3;
output [9:0] output_real_25_3;
output [9:0] output_imag_25_3;
output [9:0] output_real_26_3;
output [9:0] output_imag_26_3;
output [9:0] output_real_27_3;
output [9:0] output_imag_27_3;
output [9:0] output_real_28_3;
output [9:0] output_imag_28_3;
output [9:0] output_real_29_3;
output [9:0] output_imag_29_3;
output [9:0] output_real_30_3;
output [9:0] output_imag_30_3;
output [9:0] output_real_31_3;
output [9:0] output_imag_31_3;
output [9:0] output_real_32_3;
output [9:0] output_imag_32_3;
output [9:0] output_real_33_3;
output [9:0] output_imag_33_3;
output [9:0] output_real_34_3;
output [9:0] output_imag_34_3;
output [9:0] output_real_35_3;
output [9:0] output_imag_35_3;
output [9:0] output_real_36_3;
output [9:0] output_imag_36_3;
output [9:0] output_real_37_3;
output [9:0] output_imag_37_3;
output [9:0] output_real_38_3;
output [9:0] output_imag_38_3;
output [9:0] output_real_39_3;
output [9:0] output_imag_39_3;
output [9:0] output_real_40_3;
output [9:0] output_imag_40_3;
output [9:0] output_real_41_3;
output [9:0] output_imag_41_3;
output [9:0] output_real_42_3;
output [9:0] output_imag_42_3;
output [9:0] output_real_43_3;
output [9:0] output_imag_43_3;
output [9:0] output_real_44_3;
output [9:0] output_imag_44_3;
output [9:0] output_real_45_3;
output [9:0] output_imag_45_3;
output [9:0] output_real_46_3;
output [9:0] output_imag_46_3;
output [9:0] output_real_47_3;
output [9:0] output_imag_47_3;
output [9:0] output_real_48_3;
output [9:0] output_imag_48_3;
output [9:0] output_real_49_3;
output [9:0] output_imag_49_3;
output [9:0] output_real_50_3;
output [9:0] output_imag_50_3;
output [9:0] output_real_51_3;
output [9:0] output_imag_51_3;
output [9:0] output_real_52_3;
output [9:0] output_imag_52_3;
output [9:0] output_real_53_3;
output [9:0] output_imag_53_3;
output [9:0] output_real_54_3;
output [9:0] output_imag_54_3;
output [9:0] output_real_55_3;
output [9:0] output_imag_55_3;
output [9:0] output_real_56_3;
output [9:0] output_imag_56_3;
output [9:0] output_real_57_3;
output [9:0] output_imag_57_3;
output [9:0] output_real_58_3;
output [9:0] output_imag_58_3;
output [9:0] output_real_59_3;
output [9:0] output_imag_59_3;
output [9:0] output_real_60_3;
output [9:0] output_imag_60_3;
output [9:0] output_real_61_3;
output [9:0] output_imag_61_3;
output [9:0] output_real_62_3;
output [9:0] output_imag_62_3;
output [9:0] output_real_63_3;
output [9:0] output_imag_63_3;


always @(posedge CLK or posedge rst) begin
        if(rst==1'b1) begin
                config0_0 <= 28'b0;
                config1_0 <= 28'b0;
                config2_0 <= 28'b0;
                config3_0 <= 28'b0;
                config4_0 <= 28'b0;
                config5_0 <= 28'b0;
                config6_0 <= 28'b0;
                config7_0 <= 28'b0;
                config8_0 <= 28'b0;
                config9_0 <= 28'b0;
                config10_0 <= 28'b0;
                config11_0 <= 28'b0;
                config12_0 <= 28'b0;
                config13_0 <= 28'b0;
                config14_0 <= 28'b0;
                config15_0 <= 28'b0;
                config16_0 <= 28'b0;
                config17_0 <= 28'b0;
                config18_0 <= 28'b0;
                config19_0 <= 28'b0;
                config20_0 <= 28'b0;
                config21_0 <= 28'b0;
                config22_0 <= 28'b0;
                config23_0 <= 28'b0;
                config24_0 <= 28'b0;
                config25_0 <= 28'b0;
                config26_0 <= 28'b0;
                config27_0 <= 28'b0;
                config28_0 <= 28'b0;
                config29_0 <= 28'b0;
                config30_0 <= 28'b0;
                config31_0 <= 28'b0;
                config32_0 <= 28'b0;
                config33_0 <= 28'b0;
                config34_0 <= 28'b0;
                config35_0 <= 28'b0;
                config36_0 <= 28'b0;
                config37_0 <= 28'b0;
                config38_0 <= 28'b0;
                config39_0 <= 28'b0;
                config40_0 <= 28'b0;
                config41_0 <= 28'b0;
                config42_0 <= 28'b0;
                config43_0 <= 28'b0;
                config44_0 <= 28'b0;
                config45_0 <= 28'b0;
                config46_0 <= 28'b0;
                config47_0 <= 28'b0;
                config48_0 <= 28'b0;
                config49_0 <= 28'b0;
                config50_0 <= 28'b0;
                config51_0 <= 28'b0;
                config52_0 <= 28'b0;
                config53_0 <= 28'b0;
                config54_0 <= 28'b0;
                config55_0 <= 28'b0;
                config56_0 <= 28'b0;
                config57_0 <= 28'b0;
                config58_0 <= 28'b0;
                config59_0 <= 28'b0;
                config60_0 <= 28'b0;
                config61_0 <= 28'b0;
                config62_0 <= 28'b0;
                config63_0 <= 28'b0;

                config0_1 <= 28'b0;
                config1_1 <= 28'b0;
                config2_1 <= 28'b0;
                config3_1 <= 28'b0;
                config4_1 <= 28'b0;
                config5_1 <= 28'b0;
                config6_1 <= 28'b0;
                config7_1 <= 28'b0;
                config8_1 <= 28'b0;
                config9_1 <= 28'b0;
                config10_1 <= 28'b0;
                config11_1 <= 28'b0;
                config12_1 <= 28'b0;
                config13_1 <= 28'b0;
                config14_1 <= 28'b0;
                config15_1 <= 28'b0;
                config16_1 <= 28'b0;
                config17_1 <= 28'b0;
                config18_1 <= 28'b0;
                config19_1 <= 28'b0;
                config20_1 <= 28'b0;
                config21_1 <= 28'b0;
                config22_1 <= 28'b0;
                config23_1 <= 28'b0;
                config24_1 <= 28'b0;
                config25_1 <= 28'b0;
                config26_1 <= 28'b0;
                config27_1 <= 28'b0;
                config28_1 <= 28'b0;
                config29_1 <= 28'b0;
                config30_1 <= 28'b0;
                config31_1 <= 28'b0;
                config32_1 <= 28'b0;
                config33_1 <= 28'b0;
                config34_1 <= 28'b0;
                config35_1 <= 28'b0;
                config36_1 <= 28'b0;
                config37_1 <= 28'b0;
                config38_1 <= 28'b0;
                config39_1 <= 28'b0;
                config40_1 <= 28'b0;
                config41_1 <= 28'b0;
                config42_1 <= 28'b0;
                config43_1 <= 28'b0;
                config44_1 <= 28'b0;
                config45_1 <= 28'b0;
                config46_1 <= 28'b0;
                config47_1 <= 28'b0;
                config48_1 <= 28'b0;
                config49_1 <= 28'b0;
                config50_1 <= 28'b0;
                config51_1 <= 28'b0;
                config52_1 <= 28'b0;
                config53_1 <= 28'b0;
                config54_1 <= 28'b0;
                config55_1 <= 28'b0;
                config56_1 <= 28'b0;
                config57_1 <= 28'b0;
                config58_1 <= 28'b0;
                config59_1 <= 28'b0;
                config60_1 <= 28'b0;
                config61_1 <= 28'b0;
                config62_1 <= 28'b0;
                config63_1 <= 28'b0;

                config0_2 <= 28'b0;
                config1_2 <= 28'b0;
                config2_2 <= 28'b0;
                config3_2 <= 28'b0;
                config4_2 <= 28'b0;
                config5_2 <= 28'b0;
                config6_2 <= 28'b0;
                config7_2 <= 28'b0;
                config8_2 <= 28'b0;
                config9_2 <= 28'b0;
                config10_2 <= 28'b0;
                config11_2 <= 28'b0;
                config12_2 <= 28'b0;
                config13_2 <= 28'b0;
                config14_2 <= 28'b0;
                config15_2 <= 28'b0;
                config16_2 <= 28'b0;
                config17_2 <= 28'b0;
                config18_2 <= 28'b0;
                config19_2 <= 28'b0;
                config20_2 <= 28'b0;
                config21_2 <= 28'b0;
                config22_2 <= 28'b0;
                config23_2 <= 28'b0;
                config24_2 <= 28'b0;
                config25_2 <= 28'b0;
                config26_2 <= 28'b0;
                config27_2 <= 28'b0;
                config28_2 <= 28'b0;
                config29_2 <= 28'b0;
                config30_2 <= 28'b0;
                config31_2 <= 28'b0;
                config32_2 <= 28'b0;
                config33_2 <= 28'b0;
                config34_2 <= 28'b0;
                config35_2 <= 28'b0;
                config36_2 <= 28'b0;
                config37_2 <= 28'b0;
                config38_2 <= 28'b0;
                config39_2 <= 28'b0;
                config40_2 <= 28'b0;
                config41_2 <= 28'b0;
                config42_2 <= 28'b0;
                config43_2 <= 28'b0;
                config44_2 <= 28'b0;
                config45_2 <= 28'b0;
                config46_2 <= 28'b0;
                config47_2 <= 28'b0;
                config48_2 <= 28'b0;
                config49_2 <= 28'b0;
                config50_2 <= 28'b0;
                config51_2 <= 28'b0;
                config52_2 <= 28'b0;
                config53_2 <= 28'b0;
                config54_2 <= 28'b0;
                config55_2 <= 28'b0;
                config56_2 <= 28'b0;
                config57_2 <= 28'b0;
                config58_2 <= 28'b0;
                config59_2 <= 28'b0;
                config60_2 <= 28'b0;
                config61_2 <= 28'b0;
                config62_2 <= 28'b0;
                config63_2 <= 28'b0;

                config0_3 <= 28'b0;
                config1_3 <= 28'b0;
                config2_3 <= 28'b0;
                config3_3 <= 28'b0;
                config4_3 <= 28'b0;
                config5_3 <= 28'b0;
                config6_3 <= 28'b0;
                config7_3 <= 28'b0;
                config8_3 <= 28'b0;
                config9_3 <= 28'b0;
                config10_3 <= 28'b0;
                config11_3 <= 28'b0;
                config12_3 <= 28'b0;
                config13_3 <= 28'b0;
                config14_3 <= 28'b0;
                config15_3 <= 28'b0;
                config16_3 <= 28'b0;
                config17_3 <= 28'b0;
                config18_3 <= 28'b0;
                config19_3 <= 28'b0;
                config20_3 <= 28'b0;
                config21_3 <= 28'b0;
                config22_3 <= 28'b0;
                config23_3 <= 28'b0;
                config24_3 <= 28'b0;
                config25_3 <= 28'b0;
                config26_3 <= 28'b0;
                config27_3 <= 28'b0;
                config28_3 <= 28'b0;
                config29_3 <= 28'b0;
                config30_3 <= 28'b0;
                config31_3 <= 28'b0;
                config32_3 <= 28'b0;
                config33_3 <= 28'b0;
                config34_3 <= 28'b0;
                config35_3 <= 28'b0;
                config36_3 <= 28'b0;
                config37_3 <= 28'b0;
                config38_3 <= 28'b0;
                config39_3 <= 28'b0;
                config40_3 <= 28'b0;
                config41_3 <= 28'b0;
                config42_3 <= 28'b0;
                config43_3 <= 28'b0;
                config44_3 <= 28'b0;
                config45_3 <= 28'b0;
                config46_3 <= 28'b0;
                config47_3 <= 28'b0;
                config48_3 <= 28'b0;
                config49_3 <= 28'b0;
                config50_3 <= 28'b0;
                config51_3 <= 28'b0;
                config52_3 <= 28'b0;
                config53_3 <= 28'b0;
                config54_3 <= 28'b0;
                config55_3 <= 28'b0;
                config56_3 <= 28'b0;
                config57_3 <= 28'b0;
                config58_3 <= 28'b0;
                config59_3 <= 28'b0;
                config60_3 <= 28'b0;
                config61_3 <= 28'b0;
                config62_3 <= 28'b0;
                config63_3 <= 28'b0;
				


        end
        else begin
                if(ssb == 1'b1) begin
	                case (sdi[7:0])
		                8'd0: config0_0 <= sdi[27:8];
		                8'd1: config1_0 <= sdi[27:8];
		                8'd2: config2_0 <= sdi[27:8];
		                8'd3: config3_0 <= sdi[27:8];
		                8'd4: config4_0 <= sdi[27:8];
		                8'd5: config5_0 <= sdi[27:8];
		                8'd6: config6_0 <= sdi[27:8];
		                8'd7: config7_0 <= sdi[27:8];
		                8'd8: config8_0 <= sdi[27:8];
		                8'd9: config9_0 <= sdi[27:8];
		                8'd10: config10_0 <= sdi[27:8];
		                8'd11: config11_0 <= sdi[27:8];
		                8'd12: config12_0 <= sdi[27:8];
		                8'd13: config13_0 <= sdi[27:8];
		                8'd14: config14_0 <= sdi[27:8];
		                8'd15: config15_0 <= sdi[27:8];
		                8'd16: config16_0 <= sdi[27:8];
		                8'd17: config17_0 <= sdi[27:8];
		                8'd18: config18_0 <= sdi[27:8];
		                8'd19: config19_0 <= sdi[27:8];
		                8'd20: config20_0 <= sdi[27:8];
		                8'd21: config21_0 <= sdi[27:8];
		                8'd22: config22_0 <= sdi[27:8];
		                8'd23: config23_0 <= sdi[27:8];
		                8'd24: config24_0 <= sdi[27:8];
		                8'd25: config25_0 <= sdi[27:8];
		                8'd26: config26_0 <= sdi[27:8];
		                8'd27: config27_0 <= sdi[27:8];
		                8'd28: config28_0 <= sdi[27:8];
		                8'd29: config29_0 <= sdi[27:8];
		                8'd30: config30_0 <= sdi[27:8];
		                8'd31: config31_0 <= sdi[27:8];
		                8'd32: config32_0 <= sdi[27:8];
		                8'd33: config33_0 <= sdi[27:8];
		                8'd34: config34_0 <= sdi[27:8];
		                8'd35: config35_0 <= sdi[27:8];
		                8'd36: config36_0 <= sdi[27:8];
		                8'd37: config37_0 <= sdi[27:8];
		                8'd38: config38_0 <= sdi[27:8];
		                8'd39: config39_0 <= sdi[27:8];
		                8'd40: config40_0 <= sdi[27:8];
		                8'd41: config41_0 <= sdi[27:8];
		                8'd42: config42_0 <= sdi[27:8];
		                8'd43: config43_0 <= sdi[27:8];
		                8'd44: config44_0 <= sdi[27:8];
		                8'd45: config45_0 <= sdi[27:8];
		                8'd46: config46_0 <= sdi[27:8];
		                8'd47: config47_0 <= sdi[27:8];
		                8'd48: config48_0 <= sdi[27:8];
		                8'd49: config49_0 <= sdi[27:8];
		                8'd50: config50_0 <= sdi[27:8];
		                8'd51: config51_0 <= sdi[27:8];
		                8'd52: config52_0 <= sdi[27:8];
		                8'd53: config53_0 <= sdi[27:8];
		                8'd54: config54_0 <= sdi[27:8];
		                8'd55: config55_0 <= sdi[27:8];
		                8'd56: config56_0 <= sdi[27:8];
		                8'd57: config57_0 <= sdi[27:8];
		                8'd58: config58_0 <= sdi[27:8];
		                8'd59: config59_0 <= sdi[27:8];
		                8'd60: config60_0 <= sdi[27:8];
		                8'd61: config61_0 <= sdi[27:8];
		                8'd62: config62_0 <= sdi[27:8];
		                8'd63: config63_0 <= sdi[27:8];

		                8'd64: config0_1 <= sdi[27:8];
		                8'd65: config1_1 <= sdi[27:8];
		                8'd66: config2_1 <= sdi[27:8];
		                8'd67: config3_1 <= sdi[27:8];
		                8'd68: config4_1 <= sdi[27:8];
		                8'd69: config5_1 <= sdi[27:8];
		                8'd70: config6_1 <= sdi[27:8];
		                8'd71: config7_1 <= sdi[27:8];
		                8'd72: config8_1 <= sdi[27:8];
		                8'd73: config9_1 <= sdi[27:8];
		                8'd74: config10_1 <= sdi[27:8];
		                8'd75: config11_1 <= sdi[27:8];
		                8'd76: config12_1 <= sdi[27:8];
		                8'd77: config13_1 <= sdi[27:8];
		                8'd78: config14_1 <= sdi[27:8];
		                8'd79: config15_1 <= sdi[27:8];
		                8'd80: config16_1 <= sdi[27:8];
		                8'd81: config17_1 <= sdi[27:8];
		                8'd82: config18_1 <= sdi[27:8];
		                8'd83: config19_1 <= sdi[27:8];
		                8'd84: config20_1 <= sdi[27:8];
		                8'd85: config21_1 <= sdi[27:8];
		                8'd86: config22_1 <= sdi[27:8];
		                8'd87: config23_1 <= sdi[27:8];
		                8'd88: config24_1 <= sdi[27:8];
		                8'd89: config25_1 <= sdi[27:8];
		                8'd90: config26_1 <= sdi[27:8];
		                8'd91: config27_1 <= sdi[27:8];
		                8'd92: config28_1 <= sdi[27:8];
		                8'd93: config29_1 <= sdi[27:8];
		                8'd94: config30_1 <= sdi[27:8];
		                8'd95: config31_1 <= sdi[27:8];
		                8'd96: config32_1 <= sdi[27:8];
		                8'd97: config33_1 <= sdi[27:8];
		                8'd98: config34_1 <= sdi[27:8];
		                8'd99: config35_1 <= sdi[27:8];
		                8'd100: config36_1 <= sdi[27:8];
		                8'd101: config37_1 <= sdi[27:8];
		                8'd102: config38_1 <= sdi[27:8];
		                8'd103: config39_1 <= sdi[27:8];
		                8'd104: config40_1 <= sdi[27:8];
		                8'd105: config41_1 <= sdi[27:8];
		                8'd106: config42_1 <= sdi[27:8];
		                8'd107: config43_1 <= sdi[27:8];
		                8'd108: config44_1 <= sdi[27:8];
		                8'd109: config45_1 <= sdi[27:8];
		                8'd110: config46_1 <= sdi[27:8];
		                8'd111: config47_1 <= sdi[27:8];
		                8'd112: config48_1 <= sdi[27:8];
		                8'd113: config49_1 <= sdi[27:8];
		                8'd114: config50_1 <= sdi[27:8];
		                8'd115: config51_1 <= sdi[27:8];
		                8'd116: config52_1 <= sdi[27:8];
		                8'd117: config53_1 <= sdi[27:8];
		                8'd118: config54_1 <= sdi[27:8];
		                8'd119: config55_1 <= sdi[27:8];
		                8'd120: config56_1 <= sdi[27:8];
		                8'd121: config57_1 <= sdi[27:8];
		                8'd122: config58_1 <= sdi[27:8];
		                8'd123: config59_1 <= sdi[27:8];
		                8'd124: config60_1 <= sdi[27:8];
		                8'd125: config61_1 <= sdi[27:8];
		                8'd126: config62_1 <= sdi[27:8];
		                8'd127: config63_1 <= sdi[27:8];

		                8'd128: config0_2 <= sdi[27:8];
		                8'd129: config1_2 <= sdi[27:8];
		                8'd130: config2_2 <= sdi[27:8];
		                8'd131: config3_2 <= sdi[27:8];
		                8'd132: config4_2 <= sdi[27:8];
		                8'd133: config5_2 <= sdi[27:8];
		                8'd134: config6_2 <= sdi[27:8];
		                8'd135: config7_2 <= sdi[27:8];
		                8'd136: config8_2 <= sdi[27:8];
		                8'd137: config9_2 <= sdi[27:8];
		                8'd138: config10_2 <= sdi[27:8];
		                8'd139: config11_2 <= sdi[27:8];
		                8'd140: config12_2 <= sdi[27:8];
		                8'd141: config13_2 <= sdi[27:8];
		                8'd142: config14_2 <= sdi[27:8];
		                8'd143: config15_2 <= sdi[27:8];
		                8'd144: config16_2 <= sdi[27:8];
		                8'd145: config17_2 <= sdi[27:8];
		                8'd146: config18_2 <= sdi[27:8];
		                8'd147: config19_2 <= sdi[27:8];
		                8'd148: config20_2 <= sdi[27:8];
		                8'd149: config21_2 <= sdi[27:8];
		                8'd150: config22_2 <= sdi[27:8];
		                8'd151: config23_2 <= sdi[27:8];
		                8'd152: config24_2 <= sdi[27:8];
		                8'd153: config25_2 <= sdi[27:8];
		                8'd154: config26_2 <= sdi[27:8];
		                8'd155: config27_2 <= sdi[27:8];
		                8'd156: config28_2 <= sdi[27:8];
		                8'd157: config29_2 <= sdi[27:8];
		                8'd158: config30_2 <= sdi[27:8];
		                8'd159: config31_2 <= sdi[27:8];
		                8'd160: config32_2 <= sdi[27:8];
		                8'd161: config33_2 <= sdi[27:8];
		                8'd162: config34_2 <= sdi[27:8];
		                8'd163: config35_2 <= sdi[27:8];
		                8'd164: config36_2 <= sdi[27:8];
		                8'd165: config37_2 <= sdi[27:8];
		                8'd166: config38_2 <= sdi[27:8];
		                8'd167: config39_2 <= sdi[27:8];
		                8'd168: config40_2 <= sdi[27:8];
		                8'd169: config41_2 <= sdi[27:8];
		                8'd170: config42_2 <= sdi[27:8];
		                8'd171: config43_2 <= sdi[27:8];
		                8'd172: config44_2 <= sdi[27:8];
		                8'd173: config45_2 <= sdi[27:8];
		                8'd174: config46_2 <= sdi[27:8];
		                8'd175: config47_2 <= sdi[27:8];
		                8'd176: config48_2 <= sdi[27:8];
		                8'd177: config49_2 <= sdi[27:8];
		                8'd178: config50_2 <= sdi[27:8];
		                8'd179: config51_2 <= sdi[27:8];
		                8'd180: config52_2 <= sdi[27:8];
		                8'd181: config53_2 <= sdi[27:8];
		                8'd182: config54_2 <= sdi[27:8];
		                8'd183: config55_2 <= sdi[27:8];
		                8'd184: config56_2 <= sdi[27:8];
		                8'd185: config57_2 <= sdi[27:8];
		                8'd186: config58_2 <= sdi[27:8];
		                8'd187: config59_2 <= sdi[27:8];
		                8'd188: config60_2 <= sdi[27:8];
		                8'd189: config61_2 <= sdi[27:8];
		                8'd190: config62_2 <= sdi[27:8];
		                8'd191: config63_2 <= sdi[27:8];

		                8'd192: config0_3 <= sdi[27:8];
		                8'd193: config1_3 <= sdi[27:8];
		                8'd194: config2_3 <= sdi[27:8];
		                8'd195: config3_3 <= sdi[27:8];
		                8'd196: config4_3 <= sdi[27:8];
		                8'd197: config5_3 <= sdi[27:8];
		                8'd198: config6_3 <= sdi[27:8];
		                8'd199: config7_3 <= sdi[27:8];
		                8'd200: config8_3 <= sdi[27:8];
		                8'd201: config9_3 <= sdi[27:8];
		                8'd202: config10_3 <= sdi[27:8];
		                8'd203: config11_3 <= sdi[27:8];
		                8'd204: config12_3 <= sdi[27:8];
		                8'd205: config13_3 <= sdi[27:8];
		                8'd206: config14_3 <= sdi[27:8];
		                8'd207: config15_3 <= sdi[27:8];
		                8'd208: config16_3 <= sdi[27:8];
		                8'd209: config17_3 <= sdi[27:8];
		                8'd210: config18_3 <= sdi[27:8];
		                8'd211: config19_3 <= sdi[27:8];
		                8'd212: config20_3 <= sdi[27:8];
		                8'd213: config21_3 <= sdi[27:8];
		                8'd214: config22_3 <= sdi[27:8];
		                8'd215: config23_3 <= sdi[27:8];
		                8'd216: config24_3 <= sdi[27:8];
		                8'd217: config25_3 <= sdi[27:8];
		                8'd218: config26_3 <= sdi[27:8];
		                8'd219: config27_3 <= sdi[27:8];
		                8'd220: config28_3 <= sdi[27:8];
		                8'd221: config29_3 <= sdi[27:8];
		                8'd222: config30_3 <= sdi[27:8];
		                8'd223: config31_3 <= sdi[27:8];
		                8'd224: config32_3 <= sdi[27:8];
		                8'd225: config33_3 <= sdi[27:8];
		                8'd226: config34_3 <= sdi[27:8];
		                8'd227: config35_3 <= sdi[27:8];
		                8'd228: config36_3 <= sdi[27:8];
		                8'd229: config37_3 <= sdi[27:8];
		                8'd230: config38_3 <= sdi[27:8];
		                8'd231: config39_3 <= sdi[27:8];
		                8'd232: config40_3 <= sdi[27:8];
		                8'd233: config41_3 <= sdi[27:8];
		                8'd234: config42_3 <= sdi[27:8];
		                8'd235: config43_3 <= sdi[27:8];
		                8'd236: config44_3 <= sdi[27:8];
		                8'd237: config45_3 <= sdi[27:8];
		                8'd238: config46_3 <= sdi[27:8];
		                8'd239: config47_3 <= sdi[27:8];
		                8'd240: config48_3 <= sdi[27:8];
		                8'd241: config49_3 <= sdi[27:8];
		                8'd242: config50_3 <= sdi[27:8];
		                8'd243: config51_3 <= sdi[27:8];
		                8'd244: config52_3 <= sdi[27:8];
		                8'd245: config53_3 <= sdi[27:8];
		                8'd246: config54_3 <= sdi[27:8];
		                8'd247: config55_3 <= sdi[27:8];
		                8'd248: config56_3 <= sdi[27:8];
		                8'd249: config57_3 <= sdi[27:8];
		                8'd250: config58_3 <= sdi[27:8];
		                8'd251: config59_3 <= sdi[27:8];
		                8'd252: config60_3 <= sdi[27:8];
		                8'd253: config61_3 <= sdi[27:8];
		                8'd254: config62_3 <= sdi[27:8];
		                8'd255: config63_3 <= sdi[27:8];
                    endcase                   
                end	
                else begin
	                        config0_0 <= config0_0;
	                        config1_0 <= config1_0;
	                        config2_0 <= config2_0;
	                        config3_0 <= config3_0;
	                        config4_0 <= config4_0;
	                        config5_0 <= config5_0;
	                        config6_0 <= config6_0;
	                        config7_0 <= config7_0;
	                        config8_0 <= config8_0;
	                        config9_0 <= config9_0;
	                        config10_0 <= config10_0;
	                        config11_0 <= config11_0;
	                        config12_0 <= config12_0;
	                        config13_0 <= config13_0;
	                        config14_0 <= config14_0;
	                        config15_0 <= config15_0;
	                        config16_0 <= config16_0;
	                        config17_0 <= config17_0;
	                        config18_0 <= config18_0;
	                        config19_0 <= config19_0;
	                        config20_0 <= config20_0;
	                        config21_0 <= config21_0;
	                        config22_0 <= config22_0;
	                        config23_0 <= config23_0;
	                        config24_0 <= config24_0;
	                        config25_0 <= config25_0;
	                        config26_0 <= config26_0;
	                        config27_0 <= config27_0;
	                        config28_0 <= config28_0;
	                        config29_0 <= config29_0;
	                        config30_0 <= config30_0;
	                        config31_0 <= config31_0;
	                        config32_0 <= config32_0;
	                        config33_0 <= config33_0;
	                        config34_0 <= config34_0;
	                        config35_0 <= config35_0;
	                        config36_0 <= config36_0;
	                        config37_0 <= config37_0;
	                        config38_0 <= config38_0;
	                        config39_0 <= config39_0;
	                        config40_0 <= config40_0;
	                        config41_0 <= config41_0;
	                        config42_0 <= config42_0;
	                        config43_0 <= config43_0;
	                        config44_0 <= config44_0;
	                        config45_0 <= config45_0;
	                        config46_0 <= config46_0;
	                        config47_0 <= config47_0;
	                        config48_0 <= config48_0;
	                        config49_0 <= config49_0;
	                        config50_0 <= config50_0;
	                        config51_0 <= config51_0;
	                        config52_0 <= config52_0;
	                        config53_0 <= config53_0;
	                        config54_0 <= config54_0;
	                        config55_0 <= config55_0;
	                        config56_0 <= config56_0;
	                        config57_0 <= config57_0;
	                        config58_0 <= config58_0;
	                        config59_0 <= config59_0;
	                        config60_0 <= config60_0;
	                        config61_0 <= config61_0;
	                        config62_0 <= config62_0;
	                        config63_0 <= config63_0;

	                        config0_1 <= config0_1;
	                        config1_1 <= config1_1;
	                        config2_1 <= config2_1;
	                        config3_1 <= config3_1;
	                        config4_1 <= config4_1;
	                        config5_1 <= config5_1;
	                        config6_1 <= config6_1;
	                        config7_1 <= config7_1;
	                        config8_1 <= config8_1;
	                        config9_1 <= config9_1;
	                        config10_1 <= config10_1;
	                        config11_1 <= config11_1;
	                        config12_1 <= config12_1;
	                        config13_1 <= config13_1;
	                        config14_1 <= config14_1;
	                        config15_1 <= config15_1;
	                        config16_1 <= config16_1;
	                        config17_1 <= config17_1;
	                        config18_1 <= config18_1;
	                        config19_1 <= config19_1;
	                        config20_1 <= config20_1;
	                        config21_1 <= config21_1;
	                        config22_1 <= config22_1;
	                        config23_1 <= config23_1;
	                        config24_1 <= config24_1;
	                        config25_1 <= config25_1;
	                        config26_1 <= config26_1;
	                        config27_1 <= config27_1;
	                        config28_1 <= config28_1;
	                        config29_1 <= config29_1;
	                        config30_1 <= config30_1;
	                        config31_1 <= config31_1;
	                        config32_1 <= config32_1;
	                        config33_1 <= config33_1;
	                        config34_1 <= config34_1;
	                        config35_1 <= config35_1;
	                        config36_1 <= config36_1;
	                        config37_1 <= config37_1;
	                        config38_1 <= config38_1;
	                        config39_1 <= config39_1;
	                        config40_1 <= config40_1;
	                        config41_1 <= config41_1;
	                        config42_1 <= config42_1;
	                        config43_1 <= config43_1;
	                        config44_1 <= config44_1;
	                        config45_1 <= config45_1;
	                        config46_1 <= config46_1;
	                        config47_1 <= config47_1;
	                        config48_1 <= config48_1;
	                        config49_1 <= config49_1;
	                        config50_1 <= config50_1;
	                        config51_1 <= config51_1;
	                        config52_1 <= config52_1;
	                        config53_1 <= config53_1;
	                        config54_1 <= config54_1;
	                        config55_1 <= config55_1;
	                        config56_1 <= config56_1;
	                        config57_1 <= config57_1;
	                        config58_1 <= config58_1;
	                        config59_1 <= config59_1;
	                        config60_1 <= config60_1;
	                        config61_1 <= config61_1;
	                        config62_1 <= config62_1;
	                        config63_1 <= config63_1;

	                        config0_2 <= config0_2;
	                        config1_2 <= config1_2;
	                        config2_2 <= config2_2;
	                        config3_2 <= config3_2;
	                        config4_2 <= config4_2;
	                        config5_2 <= config5_2;
	                        config6_2 <= config6_2;
	                        config7_2 <= config7_2;
	                        config8_2 <= config8_2;
	                        config9_2 <= config9_2;
	                        config10_2 <= config10_2;
	                        config11_2 <= config11_2;
	                        config12_2 <= config12_2;
	                        config13_2 <= config13_2;
	                        config14_2 <= config14_2;
	                        config15_2 <= config15_2;
	                        config16_2 <= config16_2;
	                        config17_2 <= config17_2;
	                        config18_2 <= config18_2;
	                        config19_2 <= config19_2;
	                        config20_2 <= config20_2;
	                        config21_2 <= config21_2;
	                        config22_2 <= config22_2;
	                        config23_2 <= config23_2;
	                        config24_2 <= config24_2;
	                        config25_2 <= config25_2;
	                        config26_2 <= config26_2;
	                        config27_2 <= config27_2;
	                        config28_2 <= config28_2;
	                        config29_2 <= config29_2;
	                        config30_2 <= config30_2;
	                        config31_2 <= config31_2;
	                        config32_2 <= config32_2;
	                        config33_2 <= config33_2;
	                        config34_2 <= config34_2;
	                        config35_2 <= config35_2;
	                        config36_2 <= config36_2;
	                        config37_2 <= config37_2;
	                        config38_2 <= config38_2;
	                        config39_2 <= config39_2;
	                        config40_2 <= config40_2;
	                        config41_2 <= config41_2;
	                        config42_2 <= config42_2;
	                        config43_2 <= config43_2;
	                        config44_2 <= config44_2;
	                        config45_2 <= config45_2;
	                        config46_2 <= config46_2;
	                        config47_2 <= config47_2;
	                        config48_2 <= config48_2;
	                        config49_2 <= config49_2;
	                        config50_2 <= config50_2;
	                        config51_2 <= config51_2;
	                        config52_2 <= config52_2;
	                        config53_2 <= config53_2;
	                        config54_2 <= config54_2;
	                        config55_2 <= config55_2;
	                        config56_2 <= config56_2;
	                        config57_2 <= config57_2;
	                        config58_2 <= config58_2;
	                        config59_2 <= config59_2;
	                        config60_2 <= config60_2;
	                        config61_2 <= config61_2;
	                        config62_2 <= config62_2;
	                        config63_2 <= config63_2;

	                        config0_3 <= config0_3;
	                        config1_3 <= config1_3;
	                        config2_3 <= config2_3;
	                        config3_3 <= config3_3;
	                        config4_3 <= config4_3;
	                        config5_3 <= config5_3;
	                        config6_3 <= config6_3;
	                        config7_3 <= config7_3;
	                        config8_3 <= config8_3;
	                        config9_3 <= config9_3;
	                        config10_3 <= config10_3;
	                        config11_3 <= config11_3;
	                        config12_3 <= config12_3;
	                        config13_3 <= config13_3;
	                        config14_3 <= config14_3;
	                        config15_3 <= config15_3;
	                        config16_3 <= config16_3;
	                        config17_3 <= config17_3;
	                        config18_3 <= config18_3;
	                        config19_3 <= config19_3;
	                        config20_3 <= config20_3;
	                        config21_3 <= config21_3;
	                        config22_3 <= config22_3;
	                        config23_3 <= config23_3;
	                        config24_3 <= config24_3;
	                        config25_3 <= config25_3;
	                        config26_3 <= config26_3;
	                        config27_3 <= config27_3;
	                        config28_3 <= config28_3;
	                        config29_3 <= config29_3;
	                        config30_3 <= config30_3;
	                        config31_3 <= config31_3;
	                        config32_3 <= config32_3;
	                        config33_3 <= config33_3;
	                        config34_3 <= config34_3;
	                        config35_3 <= config35_3;
	                        config36_3 <= config36_3;
	                        config37_3 <= config37_3;
	                        config38_3 <= config38_3;
	                        config39_3 <= config39_3;
	                        config40_3 <= config40_3;
	                        config41_3 <= config41_3;
	                        config42_3 <= config42_3;
	                        config43_3 <= config43_3;
	                        config44_3 <= config44_3;
	                        config45_3 <= config45_3;
	                        config46_3 <= config46_3;
	                        config47_3 <= config47_3;
	                        config48_3 <= config48_3;
	                        config49_3 <= config49_3;
	                        config50_3 <= config50_3;
	                        config51_3 <= config51_3;
	                        config52_3 <= config52_3;
	                        config53_3 <= config53_3;
	                        config54_3 <= config54_3;
	                        config55_3 <= config55_3;
	                        config56_3 <= config56_3;
	                        config57_3 <= config57_3;
	                        config58_3 <= config58_3;
	                        config59_3 <= config59_3;
	                        config60_3 <= config60_3;
	                        config61_3 <= config61_3;
	                        config62_3 <= config62_3;
	                        config63_3 <= config63_3;

	
                end
        end
end
reg [9:0] output_real_0_0_pipe;
reg [9:0] output_imag_0_0_pipe;
reg [9:0] output_real_1_0_pipe;
reg [9:0] output_imag_1_0_pipe;
reg [9:0] output_real_2_0_pipe;
reg [9:0] output_imag_2_0_pipe;
reg [9:0] output_real_3_0_pipe;
reg [9:0] output_imag_3_0_pipe;
reg [9:0] output_real_4_0_pipe;
reg [9:0] output_imag_4_0_pipe;
reg [9:0] output_real_5_0_pipe;
reg [9:0] output_imag_5_0_pipe;
reg [9:0] output_real_6_0_pipe;
reg [9:0] output_imag_6_0_pipe;
reg [9:0] output_real_7_0_pipe;
reg [9:0] output_imag_7_0_pipe;
reg [9:0] output_real_8_0_pipe;
reg [9:0] output_imag_8_0_pipe;
reg [9:0] output_real_9_0_pipe;
reg [9:0] output_imag_9_0_pipe;
reg [9:0] output_real_10_0_pipe;
reg [9:0] output_imag_10_0_pipe;
reg [9:0] output_real_11_0_pipe;
reg [9:0] output_imag_11_0_pipe;
reg [9:0] output_real_12_0_pipe;
reg [9:0] output_imag_12_0_pipe;
reg [9:0] output_real_13_0_pipe;
reg [9:0] output_imag_13_0_pipe;
reg [9:0] output_real_14_0_pipe;
reg [9:0] output_imag_14_0_pipe;
reg [9:0] output_real_15_0_pipe;
reg [9:0] output_imag_15_0_pipe;
reg [9:0] output_real_16_0_pipe;
reg [9:0] output_imag_16_0_pipe;
reg [9:0] output_real_17_0_pipe;
reg [9:0] output_imag_17_0_pipe;
reg [9:0] output_real_18_0_pipe;
reg [9:0] output_imag_18_0_pipe;
reg [9:0] output_real_19_0_pipe;
reg [9:0] output_imag_19_0_pipe;
reg [9:0] output_real_20_0_pipe;
reg [9:0] output_imag_20_0_pipe;
reg [9:0] output_real_21_0_pipe;
reg [9:0] output_imag_21_0_pipe;
reg [9:0] output_real_22_0_pipe;
reg [9:0] output_imag_22_0_pipe;
reg [9:0] output_real_23_0_pipe;
reg [9:0] output_imag_23_0_pipe;
reg [9:0] output_real_24_0_pipe;
reg [9:0] output_imag_24_0_pipe;
reg [9:0] output_real_25_0_pipe;
reg [9:0] output_imag_25_0_pipe;
reg [9:0] output_real_26_0_pipe;
reg [9:0] output_imag_26_0_pipe;
reg [9:0] output_real_27_0_pipe;
reg [9:0] output_imag_27_0_pipe;
reg [9:0] output_real_28_0_pipe;
reg [9:0] output_imag_28_0_pipe;
reg [9:0] output_real_29_0_pipe;
reg [9:0] output_imag_29_0_pipe;
reg [9:0] output_real_30_0_pipe;
reg [9:0] output_imag_30_0_pipe;
reg [9:0] output_real_31_0_pipe;
reg [9:0] output_imag_31_0_pipe;
reg [9:0] output_real_32_0_pipe;
reg [9:0] output_imag_32_0_pipe;
reg [9:0] output_real_33_0_pipe;
reg [9:0] output_imag_33_0_pipe;
reg [9:0] output_real_34_0_pipe;
reg [9:0] output_imag_34_0_pipe;
reg [9:0] output_real_35_0_pipe;
reg [9:0] output_imag_35_0_pipe;
reg [9:0] output_real_36_0_pipe;
reg [9:0] output_imag_36_0_pipe;
reg [9:0] output_real_37_0_pipe;
reg [9:0] output_imag_37_0_pipe;
reg [9:0] output_real_38_0_pipe;
reg [9:0] output_imag_38_0_pipe;
reg [9:0] output_real_39_0_pipe;
reg [9:0] output_imag_39_0_pipe;
reg [9:0] output_real_40_0_pipe;
reg [9:0] output_imag_40_0_pipe;
reg [9:0] output_real_41_0_pipe;
reg [9:0] output_imag_41_0_pipe;
reg [9:0] output_real_42_0_pipe;
reg [9:0] output_imag_42_0_pipe;
reg [9:0] output_real_43_0_pipe;
reg [9:0] output_imag_43_0_pipe;
reg [9:0] output_real_44_0_pipe;
reg [9:0] output_imag_44_0_pipe;
reg [9:0] output_real_45_0_pipe;
reg [9:0] output_imag_45_0_pipe;
reg [9:0] output_real_46_0_pipe;
reg [9:0] output_imag_46_0_pipe;
reg [9:0] output_real_47_0_pipe;
reg [9:0] output_imag_47_0_pipe;
reg [9:0] output_real_48_0_pipe;
reg [9:0] output_imag_48_0_pipe;
reg [9:0] output_real_49_0_pipe;
reg [9:0] output_imag_49_0_pipe;
reg [9:0] output_real_50_0_pipe;
reg [9:0] output_imag_50_0_pipe;
reg [9:0] output_real_51_0_pipe;
reg [9:0] output_imag_51_0_pipe;
reg [9:0] output_real_52_0_pipe;
reg [9:0] output_imag_52_0_pipe;
reg [9:0] output_real_53_0_pipe;
reg [9:0] output_imag_53_0_pipe;
reg [9:0] output_real_54_0_pipe;
reg [9:0] output_imag_54_0_pipe;
reg [9:0] output_real_55_0_pipe;
reg [9:0] output_imag_55_0_pipe;
reg [9:0] output_real_56_0_pipe;
reg [9:0] output_imag_56_0_pipe;
reg [9:0] output_real_57_0_pipe;
reg [9:0] output_imag_57_0_pipe;
reg [9:0] output_real_58_0_pipe;
reg [9:0] output_imag_58_0_pipe;
reg [9:0] output_real_59_0_pipe;
reg [9:0] output_imag_59_0_pipe;
reg [9:0] output_real_60_0_pipe;
reg [9:0] output_imag_60_0_pipe;
reg [9:0] output_real_61_0_pipe;
reg [9:0] output_imag_61_0_pipe;
reg [9:0] output_real_62_0_pipe;
reg [9:0] output_imag_62_0_pipe;
reg [9:0] output_real_63_0_pipe;
reg [9:0] output_imag_63_0_pipe;
reg [9:0] output_real_0_1_pipe;
reg [9:0] output_imag_0_1_pipe;
reg [9:0] output_real_1_1_pipe;
reg [9:0] output_imag_1_1_pipe;
reg [9:0] output_real_2_1_pipe;
reg [9:0] output_imag_2_1_pipe;
reg [9:0] output_real_3_1_pipe;
reg [9:0] output_imag_3_1_pipe;
reg [9:0] output_real_4_1_pipe;
reg [9:0] output_imag_4_1_pipe;
reg [9:0] output_real_5_1_pipe;
reg [9:0] output_imag_5_1_pipe;
reg [9:0] output_real_6_1_pipe;
reg [9:0] output_imag_6_1_pipe;
reg [9:0] output_real_7_1_pipe;
reg [9:0] output_imag_7_1_pipe;
reg [9:0] output_real_8_1_pipe;
reg [9:0] output_imag_8_1_pipe;
reg [9:0] output_real_9_1_pipe;
reg [9:0] output_imag_9_1_pipe;
reg [9:0] output_real_10_1_pipe;
reg [9:0] output_imag_10_1_pipe;
reg [9:0] output_real_11_1_pipe;
reg [9:0] output_imag_11_1_pipe;
reg [9:0] output_real_12_1_pipe;
reg [9:0] output_imag_12_1_pipe;
reg [9:0] output_real_13_1_pipe;
reg [9:0] output_imag_13_1_pipe;
reg [9:0] output_real_14_1_pipe;
reg [9:0] output_imag_14_1_pipe;
reg [9:0] output_real_15_1_pipe;
reg [9:0] output_imag_15_1_pipe;
reg [9:0] output_real_16_1_pipe;
reg [9:0] output_imag_16_1_pipe;
reg [9:0] output_real_17_1_pipe;
reg [9:0] output_imag_17_1_pipe;
reg [9:0] output_real_18_1_pipe;
reg [9:0] output_imag_18_1_pipe;
reg [9:0] output_real_19_1_pipe;
reg [9:0] output_imag_19_1_pipe;
reg [9:0] output_real_20_1_pipe;
reg [9:0] output_imag_20_1_pipe;
reg [9:0] output_real_21_1_pipe;
reg [9:0] output_imag_21_1_pipe;
reg [9:0] output_real_22_1_pipe;
reg [9:0] output_imag_22_1_pipe;
reg [9:0] output_real_23_1_pipe;
reg [9:0] output_imag_23_1_pipe;
reg [9:0] output_real_24_1_pipe;
reg [9:0] output_imag_24_1_pipe;
reg [9:0] output_real_25_1_pipe;
reg [9:0] output_imag_25_1_pipe;
reg [9:0] output_real_26_1_pipe;
reg [9:0] output_imag_26_1_pipe;
reg [9:0] output_real_27_1_pipe;
reg [9:0] output_imag_27_1_pipe;
reg [9:0] output_real_28_1_pipe;
reg [9:0] output_imag_28_1_pipe;
reg [9:0] output_real_29_1_pipe;
reg [9:0] output_imag_29_1_pipe;
reg [9:0] output_real_30_1_pipe;
reg [9:0] output_imag_30_1_pipe;
reg [9:0] output_real_31_1_pipe;
reg [9:0] output_imag_31_1_pipe;
reg [9:0] output_real_32_1_pipe;
reg [9:0] output_imag_32_1_pipe;
reg [9:0] output_real_33_1_pipe;
reg [9:0] output_imag_33_1_pipe;
reg [9:0] output_real_34_1_pipe;
reg [9:0] output_imag_34_1_pipe;
reg [9:0] output_real_35_1_pipe;
reg [9:0] output_imag_35_1_pipe;
reg [9:0] output_real_36_1_pipe;
reg [9:0] output_imag_36_1_pipe;
reg [9:0] output_real_37_1_pipe;
reg [9:0] output_imag_37_1_pipe;
reg [9:0] output_real_38_1_pipe;
reg [9:0] output_imag_38_1_pipe;
reg [9:0] output_real_39_1_pipe;
reg [9:0] output_imag_39_1_pipe;
reg [9:0] output_real_40_1_pipe;
reg [9:0] output_imag_40_1_pipe;
reg [9:0] output_real_41_1_pipe;
reg [9:0] output_imag_41_1_pipe;
reg [9:0] output_real_42_1_pipe;
reg [9:0] output_imag_42_1_pipe;
reg [9:0] output_real_43_1_pipe;
reg [9:0] output_imag_43_1_pipe;
reg [9:0] output_real_44_1_pipe;
reg [9:0] output_imag_44_1_pipe;
reg [9:0] output_real_45_1_pipe;
reg [9:0] output_imag_45_1_pipe;
reg [9:0] output_real_46_1_pipe;
reg [9:0] output_imag_46_1_pipe;
reg [9:0] output_real_47_1_pipe;
reg [9:0] output_imag_47_1_pipe;
reg [9:0] output_real_48_1_pipe;
reg [9:0] output_imag_48_1_pipe;
reg [9:0] output_real_49_1_pipe;
reg [9:0] output_imag_49_1_pipe;
reg [9:0] output_real_50_1_pipe;
reg [9:0] output_imag_50_1_pipe;
reg [9:0] output_real_51_1_pipe;
reg [9:0] output_imag_51_1_pipe;
reg [9:0] output_real_52_1_pipe;
reg [9:0] output_imag_52_1_pipe;
reg [9:0] output_real_53_1_pipe;
reg [9:0] output_imag_53_1_pipe;
reg [9:0] output_real_54_1_pipe;
reg [9:0] output_imag_54_1_pipe;
reg [9:0] output_real_55_1_pipe;
reg [9:0] output_imag_55_1_pipe;
reg [9:0] output_real_56_1_pipe;
reg [9:0] output_imag_56_1_pipe;
reg [9:0] output_real_57_1_pipe;
reg [9:0] output_imag_57_1_pipe;
reg [9:0] output_real_58_1_pipe;
reg [9:0] output_imag_58_1_pipe;
reg [9:0] output_real_59_1_pipe;
reg [9:0] output_imag_59_1_pipe;
reg [9:0] output_real_60_1_pipe;
reg [9:0] output_imag_60_1_pipe;
reg [9:0] output_real_61_1_pipe;
reg [9:0] output_imag_61_1_pipe;
reg [9:0] output_real_62_1_pipe;
reg [9:0] output_imag_62_1_pipe;
reg [9:0] output_real_63_1_pipe;
reg [9:0] output_imag_63_1_pipe;
reg [9:0] output_real_0_2_pipe;
reg [9:0] output_imag_0_2_pipe;
reg [9:0] output_real_1_2_pipe;
reg [9:0] output_imag_1_2_pipe;
reg [9:0] output_real_2_2_pipe;
reg [9:0] output_imag_2_2_pipe;
reg [9:0] output_real_3_2_pipe;
reg [9:0] output_imag_3_2_pipe;
reg [9:0] output_real_4_2_pipe;
reg [9:0] output_imag_4_2_pipe;
reg [9:0] output_real_5_2_pipe;
reg [9:0] output_imag_5_2_pipe;
reg [9:0] output_real_6_2_pipe;
reg [9:0] output_imag_6_2_pipe;
reg [9:0] output_real_7_2_pipe;
reg [9:0] output_imag_7_2_pipe;
reg [9:0] output_real_8_2_pipe;
reg [9:0] output_imag_8_2_pipe;
reg [9:0] output_real_9_2_pipe;
reg [9:0] output_imag_9_2_pipe;
reg [9:0] output_real_10_2_pipe;
reg [9:0] output_imag_10_2_pipe;
reg [9:0] output_real_11_2_pipe;
reg [9:0] output_imag_11_2_pipe;
reg [9:0] output_real_12_2_pipe;
reg [9:0] output_imag_12_2_pipe;
reg [9:0] output_real_13_2_pipe;
reg [9:0] output_imag_13_2_pipe;
reg [9:0] output_real_14_2_pipe;
reg [9:0] output_imag_14_2_pipe;
reg [9:0] output_real_15_2_pipe;
reg [9:0] output_imag_15_2_pipe;
reg [9:0] output_real_16_2_pipe;
reg [9:0] output_imag_16_2_pipe;
reg [9:0] output_real_17_2_pipe;
reg [9:0] output_imag_17_2_pipe;
reg [9:0] output_real_18_2_pipe;
reg [9:0] output_imag_18_2_pipe;
reg [9:0] output_real_19_2_pipe;
reg [9:0] output_imag_19_2_pipe;
reg [9:0] output_real_20_2_pipe;
reg [9:0] output_imag_20_2_pipe;
reg [9:0] output_real_21_2_pipe;
reg [9:0] output_imag_21_2_pipe;
reg [9:0] output_real_22_2_pipe;
reg [9:0] output_imag_22_2_pipe;
reg [9:0] output_real_23_2_pipe;
reg [9:0] output_imag_23_2_pipe;
reg [9:0] output_real_24_2_pipe;
reg [9:0] output_imag_24_2_pipe;
reg [9:0] output_real_25_2_pipe;
reg [9:0] output_imag_25_2_pipe;
reg [9:0] output_real_26_2_pipe;
reg [9:0] output_imag_26_2_pipe;
reg [9:0] output_real_27_2_pipe;
reg [9:0] output_imag_27_2_pipe;
reg [9:0] output_real_28_2_pipe;
reg [9:0] output_imag_28_2_pipe;
reg [9:0] output_real_29_2_pipe;
reg [9:0] output_imag_29_2_pipe;
reg [9:0] output_real_30_2_pipe;
reg [9:0] output_imag_30_2_pipe;
reg [9:0] output_real_31_2_pipe;
reg [9:0] output_imag_31_2_pipe;
reg [9:0] output_real_32_2_pipe;
reg [9:0] output_imag_32_2_pipe;
reg [9:0] output_real_33_2_pipe;
reg [9:0] output_imag_33_2_pipe;
reg [9:0] output_real_34_2_pipe;
reg [9:0] output_imag_34_2_pipe;
reg [9:0] output_real_35_2_pipe;
reg [9:0] output_imag_35_2_pipe;
reg [9:0] output_real_36_2_pipe;
reg [9:0] output_imag_36_2_pipe;
reg [9:0] output_real_37_2_pipe;
reg [9:0] output_imag_37_2_pipe;
reg [9:0] output_real_38_2_pipe;
reg [9:0] output_imag_38_2_pipe;
reg [9:0] output_real_39_2_pipe;
reg [9:0] output_imag_39_2_pipe;
reg [9:0] output_real_40_2_pipe;
reg [9:0] output_imag_40_2_pipe;
reg [9:0] output_real_41_2_pipe;
reg [9:0] output_imag_41_2_pipe;
reg [9:0] output_real_42_2_pipe;
reg [9:0] output_imag_42_2_pipe;
reg [9:0] output_real_43_2_pipe;
reg [9:0] output_imag_43_2_pipe;
reg [9:0] output_real_44_2_pipe;
reg [9:0] output_imag_44_2_pipe;
reg [9:0] output_real_45_2_pipe;
reg [9:0] output_imag_45_2_pipe;
reg [9:0] output_real_46_2_pipe;
reg [9:0] output_imag_46_2_pipe;
reg [9:0] output_real_47_2_pipe;
reg [9:0] output_imag_47_2_pipe;
reg [9:0] output_real_48_2_pipe;
reg [9:0] output_imag_48_2_pipe;
reg [9:0] output_real_49_2_pipe;
reg [9:0] output_imag_49_2_pipe;
reg [9:0] output_real_50_2_pipe;
reg [9:0] output_imag_50_2_pipe;
reg [9:0] output_real_51_2_pipe;
reg [9:0] output_imag_51_2_pipe;
reg [9:0] output_real_52_2_pipe;
reg [9:0] output_imag_52_2_pipe;
reg [9:0] output_real_53_2_pipe;
reg [9:0] output_imag_53_2_pipe;
reg [9:0] output_real_54_2_pipe;
reg [9:0] output_imag_54_2_pipe;
reg [9:0] output_real_55_2_pipe;
reg [9:0] output_imag_55_2_pipe;
reg [9:0] output_real_56_2_pipe;
reg [9:0] output_imag_56_2_pipe;
reg [9:0] output_real_57_2_pipe;
reg [9:0] output_imag_57_2_pipe;
reg [9:0] output_real_58_2_pipe;
reg [9:0] output_imag_58_2_pipe;
reg [9:0] output_real_59_2_pipe;
reg [9:0] output_imag_59_2_pipe;
reg [9:0] output_real_60_2_pipe;
reg [9:0] output_imag_60_2_pipe;
reg [9:0] output_real_61_2_pipe;
reg [9:0] output_imag_61_2_pipe;
reg [9:0] output_real_62_2_pipe;
reg [9:0] output_imag_62_2_pipe;
reg [9:0] output_real_63_2_pipe;
reg [9:0] output_imag_63_2_pipe;
reg [9:0] output_real_0_3_pipe;
reg [9:0] output_imag_0_3_pipe;
reg [9:0] output_real_1_3_pipe;
reg [9:0] output_imag_1_3_pipe;
reg [9:0] output_real_2_3_pipe;
reg [9:0] output_imag_2_3_pipe;
reg [9:0] output_real_3_3_pipe;
reg [9:0] output_imag_3_3_pipe;
reg [9:0] output_real_4_3_pipe;
reg [9:0] output_imag_4_3_pipe;
reg [9:0] output_real_5_3_pipe;
reg [9:0] output_imag_5_3_pipe;
reg [9:0] output_real_6_3_pipe;
reg [9:0] output_imag_6_3_pipe;
reg [9:0] output_real_7_3_pipe;
reg [9:0] output_imag_7_3_pipe;
reg [9:0] output_real_8_3_pipe;
reg [9:0] output_imag_8_3_pipe;
reg [9:0] output_real_9_3_pipe;
reg [9:0] output_imag_9_3_pipe;
reg [9:0] output_real_10_3_pipe;
reg [9:0] output_imag_10_3_pipe;
reg [9:0] output_real_11_3_pipe;
reg [9:0] output_imag_11_3_pipe;
reg [9:0] output_real_12_3_pipe;
reg [9:0] output_imag_12_3_pipe;
reg [9:0] output_real_13_3_pipe;
reg [9:0] output_imag_13_3_pipe;
reg [9:0] output_real_14_3_pipe;
reg [9:0] output_imag_14_3_pipe;
reg [9:0] output_real_15_3_pipe;
reg [9:0] output_imag_15_3_pipe;
reg [9:0] output_real_16_3_pipe;
reg [9:0] output_imag_16_3_pipe;
reg [9:0] output_real_17_3_pipe;
reg [9:0] output_imag_17_3_pipe;
reg [9:0] output_real_18_3_pipe;
reg [9:0] output_imag_18_3_pipe;
reg [9:0] output_real_19_3_pipe;
reg [9:0] output_imag_19_3_pipe;
reg [9:0] output_real_20_3_pipe;
reg [9:0] output_imag_20_3_pipe;
reg [9:0] output_real_21_3_pipe;
reg [9:0] output_imag_21_3_pipe;
reg [9:0] output_real_22_3_pipe;
reg [9:0] output_imag_22_3_pipe;
reg [9:0] output_real_23_3_pipe;
reg [9:0] output_imag_23_3_pipe;
reg [9:0] output_real_24_3_pipe;
reg [9:0] output_imag_24_3_pipe;
reg [9:0] output_real_25_3_pipe;
reg [9:0] output_imag_25_3_pipe;
reg [9:0] output_real_26_3_pipe;
reg [9:0] output_imag_26_3_pipe;
reg [9:0] output_real_27_3_pipe;
reg [9:0] output_imag_27_3_pipe;
reg [9:0] output_real_28_3_pipe;
reg [9:0] output_imag_28_3_pipe;
reg [9:0] output_real_29_3_pipe;
reg [9:0] output_imag_29_3_pipe;
reg [9:0] output_real_30_3_pipe;
reg [9:0] output_imag_30_3_pipe;
reg [9:0] output_real_31_3_pipe;
reg [9:0] output_imag_31_3_pipe;
reg [9:0] output_real_32_3_pipe;
reg [9:0] output_imag_32_3_pipe;
reg [9:0] output_real_33_3_pipe;
reg [9:0] output_imag_33_3_pipe;
reg [9:0] output_real_34_3_pipe;
reg [9:0] output_imag_34_3_pipe;
reg [9:0] output_real_35_3_pipe;
reg [9:0] output_imag_35_3_pipe;
reg [9:0] output_real_36_3_pipe;
reg [9:0] output_imag_36_3_pipe;
reg [9:0] output_real_37_3_pipe;
reg [9:0] output_imag_37_3_pipe;
reg [9:0] output_real_38_3_pipe;
reg [9:0] output_imag_38_3_pipe;
reg [9:0] output_real_39_3_pipe;
reg [9:0] output_imag_39_3_pipe;
reg [9:0] output_real_40_3_pipe;
reg [9:0] output_imag_40_3_pipe;
reg [9:0] output_real_41_3_pipe;
reg [9:0] output_imag_41_3_pipe;
reg [9:0] output_real_42_3_pipe;
reg [9:0] output_imag_42_3_pipe;
reg [9:0] output_real_43_3_pipe;
reg [9:0] output_imag_43_3_pipe;
reg [9:0] output_real_44_3_pipe;
reg [9:0] output_imag_44_3_pipe;
reg [9:0] output_real_45_3_pipe;
reg [9:0] output_imag_45_3_pipe;
reg [9:0] output_real_46_3_pipe;
reg [9:0] output_imag_46_3_pipe;
reg [9:0] output_real_47_3_pipe;
reg [9:0] output_imag_47_3_pipe;
reg [9:0] output_real_48_3_pipe;
reg [9:0] output_imag_48_3_pipe;
reg [9:0] output_real_49_3_pipe;
reg [9:0] output_imag_49_3_pipe;
reg [9:0] output_real_50_3_pipe;
reg [9:0] output_imag_50_3_pipe;
reg [9:0] output_real_51_3_pipe;
reg [9:0] output_imag_51_3_pipe;
reg [9:0] output_real_52_3_pipe;
reg [9:0] output_imag_52_3_pipe;
reg [9:0] output_real_53_3_pipe;
reg [9:0] output_imag_53_3_pipe;
reg [9:0] output_real_54_3_pipe;
reg [9:0] output_imag_54_3_pipe;
reg [9:0] output_real_55_3_pipe;
reg [9:0] output_imag_55_3_pipe;
reg [9:0] output_real_56_3_pipe;
reg [9:0] output_imag_56_3_pipe;
reg [9:0] output_real_57_3_pipe;
reg [9:0] output_imag_57_3_pipe;
reg [9:0] output_real_58_3_pipe;
reg [9:0] output_imag_58_3_pipe;
reg [9:0] output_real_59_3_pipe;
reg [9:0] output_imag_59_3_pipe;
reg [9:0] output_real_60_3_pipe;
reg [9:0] output_imag_60_3_pipe;
reg [9:0] output_real_61_3_pipe;
reg [9:0] output_imag_61_3_pipe;
reg [9:0] output_real_62_3_pipe;
reg [9:0] output_imag_62_3_pipe;
reg [9:0] output_real_63_3_pipe;
reg [9:0] output_imag_63_3_pipe;

always @(posedge CLK or posedge rst) begin
        if(rst==1'b1) begin

                output_real_0_0_pipe <= 10'd0;
                output_imag_0_0_pipe <= 10'd0;
                output_real_1_0_pipe <= 10'd0;
                output_imag_1_0_pipe <= 10'd0;
                output_real_2_0_pipe <= 10'd0;
                output_imag_2_0_pipe <= 10'd0;
                output_real_3_0_pipe <= 10'd0;
                output_imag_3_0_pipe <= 10'd0;
                output_real_4_0_pipe <= 10'd0;
                output_imag_4_0_pipe <= 10'd0;
                output_real_5_0_pipe <= 10'd0;
                output_imag_5_0_pipe <= 10'd0;
                output_real_6_0_pipe <= 10'd0;
                output_imag_6_0_pipe <= 10'd0;
                output_real_7_0_pipe <= 10'd0;
                output_imag_7_0_pipe <= 10'd0;
                output_real_8_0_pipe <= 10'd0;
                output_imag_8_0_pipe <= 10'd0;
                output_real_9_0_pipe <= 10'd0;
                output_imag_9_0_pipe <= 10'd0;
                output_real_10_0_pipe <= 10'd0;
                output_imag_10_0_pipe <= 10'd0;
                output_real_11_0_pipe <= 10'd0;
                output_imag_11_0_pipe <= 10'd0;
                output_real_12_0_pipe <= 10'd0;
                output_imag_12_0_pipe <= 10'd0;
                output_real_13_0_pipe <= 10'd0;
                output_imag_13_0_pipe <= 10'd0;
                output_real_14_0_pipe <= 10'd0;
                output_imag_14_0_pipe <= 10'd0;
                output_real_15_0_pipe <= 10'd0;
                output_imag_15_0_pipe <= 10'd0;
                output_real_16_0_pipe <= 10'd0;
                output_imag_16_0_pipe <= 10'd0;
                output_real_17_0_pipe <= 10'd0;
                output_imag_17_0_pipe <= 10'd0;
                output_real_18_0_pipe <= 10'd0;
                output_imag_18_0_pipe <= 10'd0;
                output_real_19_0_pipe <= 10'd0;
                output_imag_19_0_pipe <= 10'd0;
                output_real_20_0_pipe <= 10'd0;
                output_imag_20_0_pipe <= 10'd0;
                output_real_21_0_pipe <= 10'd0;
                output_imag_21_0_pipe <= 10'd0;
                output_real_22_0_pipe <= 10'd0;
                output_imag_22_0_pipe <= 10'd0;
                output_real_23_0_pipe <= 10'd0;
                output_imag_23_0_pipe <= 10'd0;
                output_real_24_0_pipe <= 10'd0;
                output_imag_24_0_pipe <= 10'd0;
                output_real_25_0_pipe <= 10'd0;
                output_imag_25_0_pipe <= 10'd0;
                output_real_26_0_pipe <= 10'd0;
                output_imag_26_0_pipe <= 10'd0;
                output_real_27_0_pipe <= 10'd0;
                output_imag_27_0_pipe <= 10'd0;
                output_real_28_0_pipe <= 10'd0;
                output_imag_28_0_pipe <= 10'd0;
                output_real_29_0_pipe <= 10'd0;
                output_imag_29_0_pipe <= 10'd0;
                output_real_30_0_pipe <= 10'd0;
                output_imag_30_0_pipe <= 10'd0;
                output_real_31_0_pipe <= 10'd0;
                output_imag_31_0_pipe <= 10'd0;
                output_real_32_0_pipe <= 10'd0;
                output_imag_32_0_pipe <= 10'd0;
                output_real_33_0_pipe <= 10'd0;
                output_imag_33_0_pipe <= 10'd0;
                output_real_34_0_pipe <= 10'd0;
                output_imag_34_0_pipe <= 10'd0;
                output_real_35_0_pipe <= 10'd0;
                output_imag_35_0_pipe <= 10'd0;
                output_real_36_0_pipe <= 10'd0;
                output_imag_36_0_pipe <= 10'd0;
                output_real_37_0_pipe <= 10'd0;
                output_imag_37_0_pipe <= 10'd0;
                output_real_38_0_pipe <= 10'd0;
                output_imag_38_0_pipe <= 10'd0;
                output_real_39_0_pipe <= 10'd0;
                output_imag_39_0_pipe <= 10'd0;
                output_real_40_0_pipe <= 10'd0;
                output_imag_40_0_pipe <= 10'd0;
                output_real_41_0_pipe <= 10'd0;
                output_imag_41_0_pipe <= 10'd0;
                output_real_42_0_pipe <= 10'd0;
                output_imag_42_0_pipe <= 10'd0;
                output_real_43_0_pipe <= 10'd0;
                output_imag_43_0_pipe <= 10'd0;
                output_real_44_0_pipe <= 10'd0;
                output_imag_44_0_pipe <= 10'd0;
                output_real_45_0_pipe <= 10'd0;
                output_imag_45_0_pipe <= 10'd0;
                output_real_46_0_pipe <= 10'd0;
                output_imag_46_0_pipe <= 10'd0;
                output_real_47_0_pipe <= 10'd0;
                output_imag_47_0_pipe <= 10'd0;
                output_real_48_0_pipe <= 10'd0;
                output_imag_48_0_pipe <= 10'd0;
                output_real_49_0_pipe <= 10'd0;
                output_imag_49_0_pipe <= 10'd0;
                output_real_50_0_pipe <= 10'd0;
                output_imag_50_0_pipe <= 10'd0;
                output_real_51_0_pipe <= 10'd0;
                output_imag_51_0_pipe <= 10'd0;
                output_real_52_0_pipe <= 10'd0;
                output_imag_52_0_pipe <= 10'd0;
                output_real_53_0_pipe <= 10'd0;
                output_imag_53_0_pipe <= 10'd0;
                output_real_54_0_pipe <= 10'd0;
                output_imag_54_0_pipe <= 10'd0;
                output_real_55_0_pipe <= 10'd0;
                output_imag_55_0_pipe <= 10'd0;
                output_real_56_0_pipe <= 10'd0;
                output_imag_56_0_pipe <= 10'd0;
                output_real_57_0_pipe <= 10'd0;
                output_imag_57_0_pipe <= 10'd0;
                output_real_58_0_pipe <= 10'd0;
                output_imag_58_0_pipe <= 10'd0;
                output_real_59_0_pipe <= 10'd0;
                output_imag_59_0_pipe <= 10'd0;
                output_real_60_0_pipe <= 10'd0;
                output_imag_60_0_pipe <= 10'd0;
                output_real_61_0_pipe <= 10'd0;
                output_imag_61_0_pipe <= 10'd0;
                output_real_62_0_pipe <= 10'd0;
                output_imag_62_0_pipe <= 10'd0;
                output_real_63_0_pipe <= 10'd0;
                output_imag_63_0_pipe <= 10'd0;
                output_real_0_1_pipe <= 10'd0;
                output_imag_0_1_pipe <= 10'd0;
                output_real_1_1_pipe <= 10'd0;
                output_imag_1_1_pipe <= 10'd0;
                output_real_2_1_pipe <= 10'd0;
                output_imag_2_1_pipe <= 10'd0;
                output_real_3_1_pipe <= 10'd0;
                output_imag_3_1_pipe <= 10'd0;
                output_real_4_1_pipe <= 10'd0;
                output_imag_4_1_pipe <= 10'd0;
                output_real_5_1_pipe <= 10'd0;
                output_imag_5_1_pipe <= 10'd0;
                output_real_6_1_pipe <= 10'd0;
                output_imag_6_1_pipe <= 10'd0;
                output_real_7_1_pipe <= 10'd0;
                output_imag_7_1_pipe <= 10'd0;
                output_real_8_1_pipe <= 10'd0;
                output_imag_8_1_pipe <= 10'd0;
                output_real_9_1_pipe <= 10'd0;
                output_imag_9_1_pipe <= 10'd0;
                output_real_10_1_pipe <= 10'd0;
                output_imag_10_1_pipe <= 10'd0;
                output_real_11_1_pipe <= 10'd0;
                output_imag_11_1_pipe <= 10'd0;
                output_real_12_1_pipe <= 10'd0;
                output_imag_12_1_pipe <= 10'd0;
                output_real_13_1_pipe <= 10'd0;
                output_imag_13_1_pipe <= 10'd0;
                output_real_14_1_pipe <= 10'd0;
                output_imag_14_1_pipe <= 10'd0;
                output_real_15_1_pipe <= 10'd0;
                output_imag_15_1_pipe <= 10'd0;
                output_real_16_1_pipe <= 10'd0;
                output_imag_16_1_pipe <= 10'd0;
                output_real_17_1_pipe <= 10'd0;
                output_imag_17_1_pipe <= 10'd0;
                output_real_18_1_pipe <= 10'd0;
                output_imag_18_1_pipe <= 10'd0;
                output_real_19_1_pipe <= 10'd0;
                output_imag_19_1_pipe <= 10'd0;
                output_real_20_1_pipe <= 10'd0;
                output_imag_20_1_pipe <= 10'd0;
                output_real_21_1_pipe <= 10'd0;
                output_imag_21_1_pipe <= 10'd0;
                output_real_22_1_pipe <= 10'd0;
                output_imag_22_1_pipe <= 10'd0;
                output_real_23_1_pipe <= 10'd0;
                output_imag_23_1_pipe <= 10'd0;
                output_real_24_1_pipe <= 10'd0;
                output_imag_24_1_pipe <= 10'd0;
                output_real_25_1_pipe <= 10'd0;
                output_imag_25_1_pipe <= 10'd0;
                output_real_26_1_pipe <= 10'd0;
                output_imag_26_1_pipe <= 10'd0;
                output_real_27_1_pipe <= 10'd0;
                output_imag_27_1_pipe <= 10'd0;
                output_real_28_1_pipe <= 10'd0;
                output_imag_28_1_pipe <= 10'd0;
                output_real_29_1_pipe <= 10'd0;
                output_imag_29_1_pipe <= 10'd0;
                output_real_30_1_pipe <= 10'd0;
                output_imag_30_1_pipe <= 10'd0;
                output_real_31_1_pipe <= 10'd0;
                output_imag_31_1_pipe <= 10'd0;
                output_real_32_1_pipe <= 10'd0;
                output_imag_32_1_pipe <= 10'd0;
                output_real_33_1_pipe <= 10'd0;
                output_imag_33_1_pipe <= 10'd0;
                output_real_34_1_pipe <= 10'd0;
                output_imag_34_1_pipe <= 10'd0;
                output_real_35_1_pipe <= 10'd0;
                output_imag_35_1_pipe <= 10'd0;
                output_real_36_1_pipe <= 10'd0;
                output_imag_36_1_pipe <= 10'd0;
                output_real_37_1_pipe <= 10'd0;
                output_imag_37_1_pipe <= 10'd0;
                output_real_38_1_pipe <= 10'd0;
                output_imag_38_1_pipe <= 10'd0;
                output_real_39_1_pipe <= 10'd0;
                output_imag_39_1_pipe <= 10'd0;
                output_real_40_1_pipe <= 10'd0;
                output_imag_40_1_pipe <= 10'd0;
                output_real_41_1_pipe <= 10'd0;
                output_imag_41_1_pipe <= 10'd0;
                output_real_42_1_pipe <= 10'd0;
                output_imag_42_1_pipe <= 10'd0;
                output_real_43_1_pipe <= 10'd0;
                output_imag_43_1_pipe <= 10'd0;
                output_real_44_1_pipe <= 10'd0;
                output_imag_44_1_pipe <= 10'd0;
                output_real_45_1_pipe <= 10'd0;
                output_imag_45_1_pipe <= 10'd0;
                output_real_46_1_pipe <= 10'd0;
                output_imag_46_1_pipe <= 10'd0;
                output_real_47_1_pipe <= 10'd0;
                output_imag_47_1_pipe <= 10'd0;
                output_real_48_1_pipe <= 10'd0;
                output_imag_48_1_pipe <= 10'd0;
                output_real_49_1_pipe <= 10'd0;
                output_imag_49_1_pipe <= 10'd0;
                output_real_50_1_pipe <= 10'd0;
                output_imag_50_1_pipe <= 10'd0;
                output_real_51_1_pipe <= 10'd0;
                output_imag_51_1_pipe <= 10'd0;
                output_real_52_1_pipe <= 10'd0;
                output_imag_52_1_pipe <= 10'd0;
                output_real_53_1_pipe <= 10'd0;
                output_imag_53_1_pipe <= 10'd0;
                output_real_54_1_pipe <= 10'd0;
                output_imag_54_1_pipe <= 10'd0;
                output_real_55_1_pipe <= 10'd0;
                output_imag_55_1_pipe <= 10'd0;
                output_real_56_1_pipe <= 10'd0;
                output_imag_56_1_pipe <= 10'd0;
                output_real_57_1_pipe <= 10'd0;
                output_imag_57_1_pipe <= 10'd0;
                output_real_58_1_pipe <= 10'd0;
                output_imag_58_1_pipe <= 10'd0;
                output_real_59_1_pipe <= 10'd0;
                output_imag_59_1_pipe <= 10'd0;
                output_real_60_1_pipe <= 10'd0;
                output_imag_60_1_pipe <= 10'd0;
                output_real_61_1_pipe <= 10'd0;
                output_imag_61_1_pipe <= 10'd0;
                output_real_62_1_pipe <= 10'd0;
                output_imag_62_1_pipe <= 10'd0;
                output_real_63_1_pipe <= 10'd0;
                output_imag_63_1_pipe <= 10'd0;
                output_real_0_2_pipe <= 10'd0;
                output_imag_0_2_pipe <= 10'd0;
                output_real_1_2_pipe <= 10'd0;
                output_imag_1_2_pipe <= 10'd0;
                output_real_2_2_pipe <= 10'd0;
                output_imag_2_2_pipe <= 10'd0;
                output_real_3_2_pipe <= 10'd0;
                output_imag_3_2_pipe <= 10'd0;
                output_real_4_2_pipe <= 10'd0;
                output_imag_4_2_pipe <= 10'd0;
                output_real_5_2_pipe <= 10'd0;
                output_imag_5_2_pipe <= 10'd0;
                output_real_6_2_pipe <= 10'd0;
                output_imag_6_2_pipe <= 10'd0;
                output_real_7_2_pipe <= 10'd0;
                output_imag_7_2_pipe <= 10'd0;
                output_real_8_2_pipe <= 10'd0;
                output_imag_8_2_pipe <= 10'd0;
                output_real_9_2_pipe <= 10'd0;
                output_imag_9_2_pipe <= 10'd0;
                output_real_10_2_pipe <= 10'd0;
                output_imag_10_2_pipe <= 10'd0;
                output_real_11_2_pipe <= 10'd0;
                output_imag_11_2_pipe <= 10'd0;
                output_real_12_2_pipe <= 10'd0;
                output_imag_12_2_pipe <= 10'd0;
                output_real_13_2_pipe <= 10'd0;
                output_imag_13_2_pipe <= 10'd0;
                output_real_14_2_pipe <= 10'd0;
                output_imag_14_2_pipe <= 10'd0;
                output_real_15_2_pipe <= 10'd0;
                output_imag_15_2_pipe <= 10'd0;
                output_real_16_2_pipe <= 10'd0;
                output_imag_16_2_pipe <= 10'd0;
                output_real_17_2_pipe <= 10'd0;
                output_imag_17_2_pipe <= 10'd0;
                output_real_18_2_pipe <= 10'd0;
                output_imag_18_2_pipe <= 10'd0;
                output_real_19_2_pipe <= 10'd0;
                output_imag_19_2_pipe <= 10'd0;
                output_real_20_2_pipe <= 10'd0;
                output_imag_20_2_pipe <= 10'd0;
                output_real_21_2_pipe <= 10'd0;
                output_imag_21_2_pipe <= 10'd0;
                output_real_22_2_pipe <= 10'd0;
                output_imag_22_2_pipe <= 10'd0;
                output_real_23_2_pipe <= 10'd0;
                output_imag_23_2_pipe <= 10'd0;
                output_real_24_2_pipe <= 10'd0;
                output_imag_24_2_pipe <= 10'd0;
                output_real_25_2_pipe <= 10'd0;
                output_imag_25_2_pipe <= 10'd0;
                output_real_26_2_pipe <= 10'd0;
                output_imag_26_2_pipe <= 10'd0;
                output_real_27_2_pipe <= 10'd0;
                output_imag_27_2_pipe <= 10'd0;
                output_real_28_2_pipe <= 10'd0;
                output_imag_28_2_pipe <= 10'd0;
                output_real_29_2_pipe <= 10'd0;
                output_imag_29_2_pipe <= 10'd0;
                output_real_30_2_pipe <= 10'd0;
                output_imag_30_2_pipe <= 10'd0;
                output_real_31_2_pipe <= 10'd0;
                output_imag_31_2_pipe <= 10'd0;
                output_real_32_2_pipe <= 10'd0;
                output_imag_32_2_pipe <= 10'd0;
                output_real_33_2_pipe <= 10'd0;
                output_imag_33_2_pipe <= 10'd0;
                output_real_34_2_pipe <= 10'd0;
                output_imag_34_2_pipe <= 10'd0;
                output_real_35_2_pipe <= 10'd0;
                output_imag_35_2_pipe <= 10'd0;
                output_real_36_2_pipe <= 10'd0;
                output_imag_36_2_pipe <= 10'd0;
                output_real_37_2_pipe <= 10'd0;
                output_imag_37_2_pipe <= 10'd0;
                output_real_38_2_pipe <= 10'd0;
                output_imag_38_2_pipe <= 10'd0;
                output_real_39_2_pipe <= 10'd0;
                output_imag_39_2_pipe <= 10'd0;
                output_real_40_2_pipe <= 10'd0;
                output_imag_40_2_pipe <= 10'd0;
                output_real_41_2_pipe <= 10'd0;
                output_imag_41_2_pipe <= 10'd0;
                output_real_42_2_pipe <= 10'd0;
                output_imag_42_2_pipe <= 10'd0;
                output_real_43_2_pipe <= 10'd0;
                output_imag_43_2_pipe <= 10'd0;
                output_real_44_2_pipe <= 10'd0;
                output_imag_44_2_pipe <= 10'd0;
                output_real_45_2_pipe <= 10'd0;
                output_imag_45_2_pipe <= 10'd0;
                output_real_46_2_pipe <= 10'd0;
                output_imag_46_2_pipe <= 10'd0;
                output_real_47_2_pipe <= 10'd0;
                output_imag_47_2_pipe <= 10'd0;
                output_real_48_2_pipe <= 10'd0;
                output_imag_48_2_pipe <= 10'd0;
                output_real_49_2_pipe <= 10'd0;
                output_imag_49_2_pipe <= 10'd0;
                output_real_50_2_pipe <= 10'd0;
                output_imag_50_2_pipe <= 10'd0;
                output_real_51_2_pipe <= 10'd0;
                output_imag_51_2_pipe <= 10'd0;
                output_real_52_2_pipe <= 10'd0;
                output_imag_52_2_pipe <= 10'd0;
                output_real_53_2_pipe <= 10'd0;
                output_imag_53_2_pipe <= 10'd0;
                output_real_54_2_pipe <= 10'd0;
                output_imag_54_2_pipe <= 10'd0;
                output_real_55_2_pipe <= 10'd0;
                output_imag_55_2_pipe <= 10'd0;
                output_real_56_2_pipe <= 10'd0;
                output_imag_56_2_pipe <= 10'd0;
                output_real_57_2_pipe <= 10'd0;
                output_imag_57_2_pipe <= 10'd0;
                output_real_58_2_pipe <= 10'd0;
                output_imag_58_2_pipe <= 10'd0;
                output_real_59_2_pipe <= 10'd0;
                output_imag_59_2_pipe <= 10'd0;
                output_real_60_2_pipe <= 10'd0;
                output_imag_60_2_pipe <= 10'd0;
                output_real_61_2_pipe <= 10'd0;
                output_imag_61_2_pipe <= 10'd0;
                output_real_62_2_pipe <= 10'd0;
                output_imag_62_2_pipe <= 10'd0;
                output_real_63_2_pipe <= 10'd0;
                output_imag_63_2_pipe <= 10'd0;
                output_real_0_3_pipe <= 10'd0;
                output_imag_0_3_pipe <= 10'd0;
                output_real_1_3_pipe <= 10'd0;
                output_imag_1_3_pipe <= 10'd0;
                output_real_2_3_pipe <= 10'd0;
                output_imag_2_3_pipe <= 10'd0;
                output_real_3_3_pipe <= 10'd0;
                output_imag_3_3_pipe <= 10'd0;
                output_real_4_3_pipe <= 10'd0;
                output_imag_4_3_pipe <= 10'd0;
                output_real_5_3_pipe <= 10'd0;
                output_imag_5_3_pipe <= 10'd0;
                output_real_6_3_pipe <= 10'd0;
                output_imag_6_3_pipe <= 10'd0;
                output_real_7_3_pipe <= 10'd0;
                output_imag_7_3_pipe <= 10'd0;
                output_real_8_3_pipe <= 10'd0;
                output_imag_8_3_pipe <= 10'd0;
                output_real_9_3_pipe <= 10'd0;
                output_imag_9_3_pipe <= 10'd0;
                output_real_10_3_pipe <= 10'd0;
                output_imag_10_3_pipe <= 10'd0;
                output_real_11_3_pipe <= 10'd0;
                output_imag_11_3_pipe <= 10'd0;
                output_real_12_3_pipe <= 10'd0;
                output_imag_12_3_pipe <= 10'd0;
                output_real_13_3_pipe <= 10'd0;
                output_imag_13_3_pipe <= 10'd0;
                output_real_14_3_pipe <= 10'd0;
                output_imag_14_3_pipe <= 10'd0;
                output_real_15_3_pipe <= 10'd0;
                output_imag_15_3_pipe <= 10'd0;
                output_real_16_3_pipe <= 10'd0;
                output_imag_16_3_pipe <= 10'd0;
                output_real_17_3_pipe <= 10'd0;
                output_imag_17_3_pipe <= 10'd0;
                output_real_18_3_pipe <= 10'd0;
                output_imag_18_3_pipe <= 10'd0;
                output_real_19_3_pipe <= 10'd0;
                output_imag_19_3_pipe <= 10'd0;
                output_real_20_3_pipe <= 10'd0;
                output_imag_20_3_pipe <= 10'd0;
                output_real_21_3_pipe <= 10'd0;
                output_imag_21_3_pipe <= 10'd0;
                output_real_22_3_pipe <= 10'd0;
                output_imag_22_3_pipe <= 10'd0;
                output_real_23_3_pipe <= 10'd0;
                output_imag_23_3_pipe <= 10'd0;
                output_real_24_3_pipe <= 10'd0;
                output_imag_24_3_pipe <= 10'd0;
                output_real_25_3_pipe <= 10'd0;
                output_imag_25_3_pipe <= 10'd0;
                output_real_26_3_pipe <= 10'd0;
                output_imag_26_3_pipe <= 10'd0;
                output_real_27_3_pipe <= 10'd0;
                output_imag_27_3_pipe <= 10'd0;
                output_real_28_3_pipe <= 10'd0;
                output_imag_28_3_pipe <= 10'd0;
                output_real_29_3_pipe <= 10'd0;
                output_imag_29_3_pipe <= 10'd0;
                output_real_30_3_pipe <= 10'd0;
                output_imag_30_3_pipe <= 10'd0;
                output_real_31_3_pipe <= 10'd0;
                output_imag_31_3_pipe <= 10'd0;
                output_real_32_3_pipe <= 10'd0;
                output_imag_32_3_pipe <= 10'd0;
                output_real_33_3_pipe <= 10'd0;
                output_imag_33_3_pipe <= 10'd0;
                output_real_34_3_pipe <= 10'd0;
                output_imag_34_3_pipe <= 10'd0;
                output_real_35_3_pipe <= 10'd0;
                output_imag_35_3_pipe <= 10'd0;
                output_real_36_3_pipe <= 10'd0;
                output_imag_36_3_pipe <= 10'd0;
                output_real_37_3_pipe <= 10'd0;
                output_imag_37_3_pipe <= 10'd0;
                output_real_38_3_pipe <= 10'd0;
                output_imag_38_3_pipe <= 10'd0;
                output_real_39_3_pipe <= 10'd0;
                output_imag_39_3_pipe <= 10'd0;
                output_real_40_3_pipe <= 10'd0;
                output_imag_40_3_pipe <= 10'd0;
                output_real_41_3_pipe <= 10'd0;
                output_imag_41_3_pipe <= 10'd0;
                output_real_42_3_pipe <= 10'd0;
                output_imag_42_3_pipe <= 10'd0;
                output_real_43_3_pipe <= 10'd0;
                output_imag_43_3_pipe <= 10'd0;
                output_real_44_3_pipe <= 10'd0;
                output_imag_44_3_pipe <= 10'd0;
                output_real_45_3_pipe <= 10'd0;
                output_imag_45_3_pipe <= 10'd0;
                output_real_46_3_pipe <= 10'd0;
                output_imag_46_3_pipe <= 10'd0;
                output_real_47_3_pipe <= 10'd0;
                output_imag_47_3_pipe <= 10'd0;
                output_real_48_3_pipe <= 10'd0;
                output_imag_48_3_pipe <= 10'd0;
                output_real_49_3_pipe <= 10'd0;
                output_imag_49_3_pipe <= 10'd0;
                output_real_50_3_pipe <= 10'd0;
                output_imag_50_3_pipe <= 10'd0;
                output_real_51_3_pipe <= 10'd0;
                output_imag_51_3_pipe <= 10'd0;
                output_real_52_3_pipe <= 10'd0;
                output_imag_52_3_pipe <= 10'd0;
                output_real_53_3_pipe <= 10'd0;
                output_imag_53_3_pipe <= 10'd0;
                output_real_54_3_pipe <= 10'd0;
                output_imag_54_3_pipe <= 10'd0;
                output_real_55_3_pipe <= 10'd0;
                output_imag_55_3_pipe <= 10'd0;
                output_real_56_3_pipe <= 10'd0;
                output_imag_56_3_pipe <= 10'd0;
                output_real_57_3_pipe <= 10'd0;
                output_imag_57_3_pipe <= 10'd0;
                output_real_58_3_pipe <= 10'd0;
                output_imag_58_3_pipe <= 10'd0;
                output_real_59_3_pipe <= 10'd0;
                output_imag_59_3_pipe <= 10'd0;
                output_real_60_3_pipe <= 10'd0;
                output_imag_60_3_pipe <= 10'd0;
                output_real_61_3_pipe <= 10'd0;
                output_imag_61_3_pipe <= 10'd0;
                output_real_62_3_pipe <= 10'd0;
                output_imag_62_3_pipe <= 10'd0;
                output_real_63_3_pipe <= 10'd0;
                output_imag_63_3_pipe <= 10'd0;

        end
        else begin
        if (vmm_load == 1'b1) begin
                output_real_0_0_pipe <= config0_0[19:10];
                output_imag_0_0_pipe <= config0_0[9:0];
                output_real_1_0_pipe <= config1_0[19:10];
                output_imag_1_0_pipe <= config1_0[9:0];
                output_real_2_0_pipe <= config2_0[19:10];
                output_imag_2_0_pipe <= config2_0[9:0];
                output_real_3_0_pipe <= config3_0[19:10];
                output_imag_3_0_pipe <= config3_0[9:0];
                output_real_4_0_pipe <= config4_0[19:10];
                output_imag_4_0_pipe <= config4_0[9:0];
                output_real_5_0_pipe <= config5_0[19:10];
                output_imag_5_0_pipe <= config5_0[9:0];
                output_real_6_0_pipe <= config6_0[19:10];
                output_imag_6_0_pipe <= config6_0[9:0];
                output_real_7_0_pipe <= config7_0[19:10];
                output_imag_7_0_pipe <= config7_0[9:0];
                output_real_8_0_pipe <= config8_0[19:10];
                output_imag_8_0_pipe <= config8_0[9:0];
                output_real_9_0_pipe <= config9_0[19:10];
                output_imag_9_0_pipe <= config9_0[9:0];
                output_real_10_0_pipe <= config10_0[19:10];
                output_imag_10_0_pipe <= config10_0[9:0];
                output_real_11_0_pipe <= config11_0[19:10];
                output_imag_11_0_pipe <= config11_0[9:0];
                output_real_12_0_pipe <= config12_0[19:10];
                output_imag_12_0_pipe <= config12_0[9:0];
                output_real_13_0_pipe <= config13_0[19:10];
                output_imag_13_0_pipe <= config13_0[9:0];
                output_real_14_0_pipe <= config14_0[19:10];
                output_imag_14_0_pipe <= config14_0[9:0];
                output_real_15_0_pipe <= config15_0[19:10];
                output_imag_15_0_pipe <= config15_0[9:0];
                output_real_16_0_pipe <= config16_0[19:10];
                output_imag_16_0_pipe <= config16_0[9:0];
                output_real_17_0_pipe <= config17_0[19:10];
                output_imag_17_0_pipe <= config17_0[9:0];
                output_real_18_0_pipe <= config18_0[19:10];
                output_imag_18_0_pipe <= config18_0[9:0];
                output_real_19_0_pipe <= config19_0[19:10];
                output_imag_19_0_pipe <= config19_0[9:0];
                output_real_20_0_pipe <= config20_0[19:10];
                output_imag_20_0_pipe <= config20_0[9:0];
                output_real_21_0_pipe <= config21_0[19:10];
                output_imag_21_0_pipe <= config21_0[9:0];
                output_real_22_0_pipe <= config22_0[19:10];
                output_imag_22_0_pipe <= config22_0[9:0];
                output_real_23_0_pipe <= config23_0[19:10];
                output_imag_23_0_pipe <= config23_0[9:0];
                output_real_24_0_pipe <= config24_0[19:10];
                output_imag_24_0_pipe <= config24_0[9:0];
                output_real_25_0_pipe <= config25_0[19:10];
                output_imag_25_0_pipe <= config25_0[9:0];
                output_real_26_0_pipe <= config26_0[19:10];
                output_imag_26_0_pipe <= config26_0[9:0];
                output_real_27_0_pipe <= config27_0[19:10];
                output_imag_27_0_pipe <= config27_0[9:0];
                output_real_28_0_pipe <= config28_0[19:10];
                output_imag_28_0_pipe <= config28_0[9:0];
                output_real_29_0_pipe <= config29_0[19:10];
                output_imag_29_0_pipe <= config29_0[9:0];
                output_real_30_0_pipe <= config30_0[19:10];
                output_imag_30_0_pipe <= config30_0[9:0];
                output_real_31_0_pipe <= config31_0[19:10];
                output_imag_31_0_pipe <= config31_0[9:0];
                output_real_32_0_pipe <= config32_0[19:10];
                output_imag_32_0_pipe <= config32_0[9:0];
                output_real_33_0_pipe <= config33_0[19:10];
                output_imag_33_0_pipe <= config33_0[9:0];
                output_real_34_0_pipe <= config34_0[19:10];
                output_imag_34_0_pipe <= config34_0[9:0];
                output_real_35_0_pipe <= config35_0[19:10];
                output_imag_35_0_pipe <= config35_0[9:0];
                output_real_36_0_pipe <= config36_0[19:10];
                output_imag_36_0_pipe <= config36_0[9:0];
                output_real_37_0_pipe <= config37_0[19:10];
                output_imag_37_0_pipe <= config37_0[9:0];
                output_real_38_0_pipe <= config38_0[19:10];
                output_imag_38_0_pipe <= config38_0[9:0];
                output_real_39_0_pipe <= config39_0[19:10];
                output_imag_39_0_pipe <= config39_0[9:0];
                output_real_40_0_pipe <= config40_0[19:10];
                output_imag_40_0_pipe <= config40_0[9:0];
                output_real_41_0_pipe <= config41_0[19:10];
                output_imag_41_0_pipe <= config41_0[9:0];
                output_real_42_0_pipe <= config42_0[19:10];
                output_imag_42_0_pipe <= config42_0[9:0];
                output_real_43_0_pipe <= config43_0[19:10];
                output_imag_43_0_pipe <= config43_0[9:0];
                output_real_44_0_pipe <= config44_0[19:10];
                output_imag_44_0_pipe <= config44_0[9:0];
                output_real_45_0_pipe <= config45_0[19:10];
                output_imag_45_0_pipe <= config45_0[9:0];
                output_real_46_0_pipe <= config46_0[19:10];
                output_imag_46_0_pipe <= config46_0[9:0];
                output_real_47_0_pipe <= config47_0[19:10];
                output_imag_47_0_pipe <= config47_0[9:0];
                output_real_48_0_pipe <= config48_0[19:10];
                output_imag_48_0_pipe <= config48_0[9:0];
                output_real_49_0_pipe <= config49_0[19:10];
                output_imag_49_0_pipe <= config49_0[9:0];
                output_real_50_0_pipe <= config50_0[19:10];
                output_imag_50_0_pipe <= config50_0[9:0];
                output_real_51_0_pipe <= config51_0[19:10];
                output_imag_51_0_pipe <= config51_0[9:0];
                output_real_52_0_pipe <= config52_0[19:10];
                output_imag_52_0_pipe <= config52_0[9:0];
                output_real_53_0_pipe <= config53_0[19:10];
                output_imag_53_0_pipe <= config53_0[9:0];
                output_real_54_0_pipe <= config54_0[19:10];
                output_imag_54_0_pipe <= config54_0[9:0];
                output_real_55_0_pipe <= config55_0[19:10];
                output_imag_55_0_pipe <= config55_0[9:0];
                output_real_56_0_pipe <= config56_0[19:10];
                output_imag_56_0_pipe <= config56_0[9:0];
                output_real_57_0_pipe <= config57_0[19:10];
                output_imag_57_0_pipe <= config57_0[9:0];
                output_real_58_0_pipe <= config58_0[19:10];
                output_imag_58_0_pipe <= config58_0[9:0];
                output_real_59_0_pipe <= config59_0[19:10];
                output_imag_59_0_pipe <= config59_0[9:0];
                output_real_60_0_pipe <= config60_0[19:10];
                output_imag_60_0_pipe <= config60_0[9:0];
                output_real_61_0_pipe <= config61_0[19:10];
                output_imag_61_0_pipe <= config61_0[9:0];
                output_real_62_0_pipe <= config62_0[19:10];
                output_imag_62_0_pipe <= config62_0[9:0];
                output_real_63_0_pipe <= config63_0[19:10];
                output_imag_63_0_pipe <= config63_0[9:0];
                output_real_0_1_pipe <= config0_1[19:10];
                output_imag_0_1_pipe <= config0_1[9:0];
                output_real_1_1_pipe <= config1_1[19:10];
                output_imag_1_1_pipe <= config1_1[9:0];
                output_real_2_1_pipe <= config2_1[19:10];
                output_imag_2_1_pipe <= config2_1[9:0];
                output_real_3_1_pipe <= config3_1[19:10];
                output_imag_3_1_pipe <= config3_1[9:0];
                output_real_4_1_pipe <= config4_1[19:10];
                output_imag_4_1_pipe <= config4_1[9:0];
                output_real_5_1_pipe <= config5_1[19:10];
                output_imag_5_1_pipe <= config5_1[9:0];
                output_real_6_1_pipe <= config6_1[19:10];
                output_imag_6_1_pipe <= config6_1[9:0];
                output_real_7_1_pipe <= config7_1[19:10];
                output_imag_7_1_pipe <= config7_1[9:0];
                output_real_8_1_pipe <= config8_1[19:10];
                output_imag_8_1_pipe <= config8_1[9:0];
                output_real_9_1_pipe <= config9_1[19:10];
                output_imag_9_1_pipe <= config9_1[9:0];
                output_real_10_1_pipe <= config10_1[19:10];
                output_imag_10_1_pipe <= config10_1[9:0];
                output_real_11_1_pipe <= config11_1[19:10];
                output_imag_11_1_pipe <= config11_1[9:0];
                output_real_12_1_pipe <= config12_1[19:10];
                output_imag_12_1_pipe <= config12_1[9:0];
                output_real_13_1_pipe <= config13_1[19:10];
                output_imag_13_1_pipe <= config13_1[9:0];
                output_real_14_1_pipe <= config14_1[19:10];
                output_imag_14_1_pipe <= config14_1[9:0];
                output_real_15_1_pipe <= config15_1[19:10];
                output_imag_15_1_pipe <= config15_1[9:0];
                output_real_16_1_pipe <= config16_1[19:10];
                output_imag_16_1_pipe <= config16_1[9:0];
                output_real_17_1_pipe <= config17_1[19:10];
                output_imag_17_1_pipe <= config17_1[9:0];
                output_real_18_1_pipe <= config18_1[19:10];
                output_imag_18_1_pipe <= config18_1[9:0];
                output_real_19_1_pipe <= config19_1[19:10];
                output_imag_19_1_pipe <= config19_1[9:0];
                output_real_20_1_pipe <= config20_1[19:10];
                output_imag_20_1_pipe <= config20_1[9:0];
                output_real_21_1_pipe <= config21_1[19:10];
                output_imag_21_1_pipe <= config21_1[9:0];
                output_real_22_1_pipe <= config22_1[19:10];
                output_imag_22_1_pipe <= config22_1[9:0];
                output_real_23_1_pipe <= config23_1[19:10];
                output_imag_23_1_pipe <= config23_1[9:0];
                output_real_24_1_pipe <= config24_1[19:10];
                output_imag_24_1_pipe <= config24_1[9:0];
                output_real_25_1_pipe <= config25_1[19:10];
                output_imag_25_1_pipe <= config25_1[9:0];
                output_real_26_1_pipe <= config26_1[19:10];
                output_imag_26_1_pipe <= config26_1[9:0];
                output_real_27_1_pipe <= config27_1[19:10];
                output_imag_27_1_pipe <= config27_1[9:0];
                output_real_28_1_pipe <= config28_1[19:10];
                output_imag_28_1_pipe <= config28_1[9:0];
                output_real_29_1_pipe <= config29_1[19:10];
                output_imag_29_1_pipe <= config29_1[9:0];
                output_real_30_1_pipe <= config30_1[19:10];
                output_imag_30_1_pipe <= config30_1[9:0];
                output_real_31_1_pipe <= config31_1[19:10];
                output_imag_31_1_pipe <= config31_1[9:0];
                output_real_32_1_pipe <= config32_1[19:10];
                output_imag_32_1_pipe <= config32_1[9:0];
                output_real_33_1_pipe <= config33_1[19:10];
                output_imag_33_1_pipe <= config33_1[9:0];
                output_real_34_1_pipe <= config34_1[19:10];
                output_imag_34_1_pipe <= config34_1[9:0];
                output_real_35_1_pipe <= config35_1[19:10];
                output_imag_35_1_pipe <= config35_1[9:0];
                output_real_36_1_pipe <= config36_1[19:10];
                output_imag_36_1_pipe <= config36_1[9:0];
                output_real_37_1_pipe <= config37_1[19:10];
                output_imag_37_1_pipe <= config37_1[9:0];
                output_real_38_1_pipe <= config38_1[19:10];
                output_imag_38_1_pipe <= config38_1[9:0];
                output_real_39_1_pipe <= config39_1[19:10];
                output_imag_39_1_pipe <= config39_1[9:0];
                output_real_40_1_pipe <= config40_1[19:10];
                output_imag_40_1_pipe <= config40_1[9:0];
                output_real_41_1_pipe <= config41_1[19:10];
                output_imag_41_1_pipe <= config41_1[9:0];
                output_real_42_1_pipe <= config42_1[19:10];
                output_imag_42_1_pipe <= config42_1[9:0];
                output_real_43_1_pipe <= config43_1[19:10];
                output_imag_43_1_pipe <= config43_1[9:0];
                output_real_44_1_pipe <= config44_1[19:10];
                output_imag_44_1_pipe <= config44_1[9:0];
                output_real_45_1_pipe <= config45_1[19:10];
                output_imag_45_1_pipe <= config45_1[9:0];
                output_real_46_1_pipe <= config46_1[19:10];
                output_imag_46_1_pipe <= config46_1[9:0];
                output_real_47_1_pipe <= config47_1[19:10];
                output_imag_47_1_pipe <= config47_1[9:0];
                output_real_48_1_pipe <= config48_1[19:10];
                output_imag_48_1_pipe <= config48_1[9:0];
                output_real_49_1_pipe <= config49_1[19:10];
                output_imag_49_1_pipe <= config49_1[9:0];
                output_real_50_1_pipe <= config50_1[19:10];
                output_imag_50_1_pipe <= config50_1[9:0];
                output_real_51_1_pipe <= config51_1[19:10];
                output_imag_51_1_pipe <= config51_1[9:0];
                output_real_52_1_pipe <= config52_1[19:10];
                output_imag_52_1_pipe <= config52_1[9:0];
                output_real_53_1_pipe <= config53_1[19:10];
                output_imag_53_1_pipe <= config53_1[9:0];
                output_real_54_1_pipe <= config54_1[19:10];
                output_imag_54_1_pipe <= config54_1[9:0];
                output_real_55_1_pipe <= config55_1[19:10];
                output_imag_55_1_pipe <= config55_1[9:0];
                output_real_56_1_pipe <= config56_1[19:10];
                output_imag_56_1_pipe <= config56_1[9:0];
                output_real_57_1_pipe <= config57_1[19:10];
                output_imag_57_1_pipe <= config57_1[9:0];
                output_real_58_1_pipe <= config58_1[19:10];
                output_imag_58_1_pipe <= config58_1[9:0];
                output_real_59_1_pipe <= config59_1[19:10];
                output_imag_59_1_pipe <= config59_1[9:0];
                output_real_60_1_pipe <= config60_1[19:10];
                output_imag_60_1_pipe <= config60_1[9:0];
                output_real_61_1_pipe <= config61_1[19:10];
                output_imag_61_1_pipe <= config61_1[9:0];
                output_real_62_1_pipe <= config62_1[19:10];
                output_imag_62_1_pipe <= config62_1[9:0];
                output_real_63_1_pipe <= config63_1[19:10];
                output_imag_63_1_pipe <= config63_1[9:0];
                output_real_0_2_pipe <= config0_2[19:10];
                output_imag_0_2_pipe <= config0_2[9:0];
                output_real_1_2_pipe <= config1_2[19:10];
                output_imag_1_2_pipe <= config1_2[9:0];
                output_real_2_2_pipe <= config2_2[19:10];
                output_imag_2_2_pipe <= config2_2[9:0];
                output_real_3_2_pipe <= config3_2[19:10];
                output_imag_3_2_pipe <= config3_2[9:0];
                output_real_4_2_pipe <= config4_2[19:10];
                output_imag_4_2_pipe <= config4_2[9:0];
                output_real_5_2_pipe <= config5_2[19:10];
                output_imag_5_2_pipe <= config5_2[9:0];
                output_real_6_2_pipe <= config6_2[19:10];
                output_imag_6_2_pipe <= config6_2[9:0];
                output_real_7_2_pipe <= config7_2[19:10];
                output_imag_7_2_pipe <= config7_2[9:0];
                output_real_8_2_pipe <= config8_2[19:10];
                output_imag_8_2_pipe <= config8_2[9:0];
                output_real_9_2_pipe <= config9_2[19:10];
                output_imag_9_2_pipe <= config9_2[9:0];
                output_real_10_2_pipe <= config10_2[19:10];
                output_imag_10_2_pipe <= config10_2[9:0];
                output_real_11_2_pipe <= config11_2[19:10];
                output_imag_11_2_pipe <= config11_2[9:0];
                output_real_12_2_pipe <= config12_2[19:10];
                output_imag_12_2_pipe <= config12_2[9:0];
                output_real_13_2_pipe <= config13_2[19:10];
                output_imag_13_2_pipe <= config13_2[9:0];
                output_real_14_2_pipe <= config14_2[19:10];
                output_imag_14_2_pipe <= config14_2[9:0];
                output_real_15_2_pipe <= config15_2[19:10];
                output_imag_15_2_pipe <= config15_2[9:0];
                output_real_16_2_pipe <= config16_2[19:10];
                output_imag_16_2_pipe <= config16_2[9:0];
                output_real_17_2_pipe <= config17_2[19:10];
                output_imag_17_2_pipe <= config17_2[9:0];
                output_real_18_2_pipe <= config18_2[19:10];
                output_imag_18_2_pipe <= config18_2[9:0];
                output_real_19_2_pipe <= config19_2[19:10];
                output_imag_19_2_pipe <= config19_2[9:0];
                output_real_20_2_pipe <= config20_2[19:10];
                output_imag_20_2_pipe <= config20_2[9:0];
                output_real_21_2_pipe <= config21_2[19:10];
                output_imag_21_2_pipe <= config21_2[9:0];
                output_real_22_2_pipe <= config22_2[19:10];
                output_imag_22_2_pipe <= config22_2[9:0];
                output_real_23_2_pipe <= config23_2[19:10];
                output_imag_23_2_pipe <= config23_2[9:0];
                output_real_24_2_pipe <= config24_2[19:10];
                output_imag_24_2_pipe <= config24_2[9:0];
                output_real_25_2_pipe <= config25_2[19:10];
                output_imag_25_2_pipe <= config25_2[9:0];
                output_real_26_2_pipe <= config26_2[19:10];
                output_imag_26_2_pipe <= config26_2[9:0];
                output_real_27_2_pipe <= config27_2[19:10];
                output_imag_27_2_pipe <= config27_2[9:0];
                output_real_28_2_pipe <= config28_2[19:10];
                output_imag_28_2_pipe <= config28_2[9:0];
                output_real_29_2_pipe <= config29_2[19:10];
                output_imag_29_2_pipe <= config29_2[9:0];
                output_real_30_2_pipe <= config30_2[19:10];
                output_imag_30_2_pipe <= config30_2[9:0];
                output_real_31_2_pipe <= config31_2[19:10];
                output_imag_31_2_pipe <= config31_2[9:0];
                output_real_32_2_pipe <= config32_2[19:10];
                output_imag_32_2_pipe <= config32_2[9:0];
                output_real_33_2_pipe <= config33_2[19:10];
                output_imag_33_2_pipe <= config33_2[9:0];
                output_real_34_2_pipe <= config34_2[19:10];
                output_imag_34_2_pipe <= config34_2[9:0];
                output_real_35_2_pipe <= config35_2[19:10];
                output_imag_35_2_pipe <= config35_2[9:0];
                output_real_36_2_pipe <= config36_2[19:10];
                output_imag_36_2_pipe <= config36_2[9:0];
                output_real_37_2_pipe <= config37_2[19:10];
                output_imag_37_2_pipe <= config37_2[9:0];
                output_real_38_2_pipe <= config38_2[19:10];
                output_imag_38_2_pipe <= config38_2[9:0];
                output_real_39_2_pipe <= config39_2[19:10];
                output_imag_39_2_pipe <= config39_2[9:0];
                output_real_40_2_pipe <= config40_2[19:10];
                output_imag_40_2_pipe <= config40_2[9:0];
                output_real_41_2_pipe <= config41_2[19:10];
                output_imag_41_2_pipe <= config41_2[9:0];
                output_real_42_2_pipe <= config42_2[19:10];
                output_imag_42_2_pipe <= config42_2[9:0];
                output_real_43_2_pipe <= config43_2[19:10];
                output_imag_43_2_pipe <= config43_2[9:0];
                output_real_44_2_pipe <= config44_2[19:10];
                output_imag_44_2_pipe <= config44_2[9:0];
                output_real_45_2_pipe <= config45_2[19:10];
                output_imag_45_2_pipe <= config45_2[9:0];
                output_real_46_2_pipe <= config46_2[19:10];
                output_imag_46_2_pipe <= config46_2[9:0];
                output_real_47_2_pipe <= config47_2[19:10];
                output_imag_47_2_pipe <= config47_2[9:0];
                output_real_48_2_pipe <= config48_2[19:10];
                output_imag_48_2_pipe <= config48_2[9:0];
                output_real_49_2_pipe <= config49_2[19:10];
                output_imag_49_2_pipe <= config49_2[9:0];
                output_real_50_2_pipe <= config50_2[19:10];
                output_imag_50_2_pipe <= config50_2[9:0];
                output_real_51_2_pipe <= config51_2[19:10];
                output_imag_51_2_pipe <= config51_2[9:0];
                output_real_52_2_pipe <= config52_2[19:10];
                output_imag_52_2_pipe <= config52_2[9:0];
                output_real_53_2_pipe <= config53_2[19:10];
                output_imag_53_2_pipe <= config53_2[9:0];
                output_real_54_2_pipe <= config54_2[19:10];
                output_imag_54_2_pipe <= config54_2[9:0];
                output_real_55_2_pipe <= config55_2[19:10];
                output_imag_55_2_pipe <= config55_2[9:0];
                output_real_56_2_pipe <= config56_2[19:10];
                output_imag_56_2_pipe <= config56_2[9:0];
                output_real_57_2_pipe <= config57_2[19:10];
                output_imag_57_2_pipe <= config57_2[9:0];
                output_real_58_2_pipe <= config58_2[19:10];
                output_imag_58_2_pipe <= config58_2[9:0];
                output_real_59_2_pipe <= config59_2[19:10];
                output_imag_59_2_pipe <= config59_2[9:0];
                output_real_60_2_pipe <= config60_2[19:10];
                output_imag_60_2_pipe <= config60_2[9:0];
                output_real_61_2_pipe <= config61_2[19:10];
                output_imag_61_2_pipe <= config61_2[9:0];
                output_real_62_2_pipe <= config62_2[19:10];
                output_imag_62_2_pipe <= config62_2[9:0];
                output_real_63_2_pipe <= config63_2[19:10];
                output_imag_63_2_pipe <= config63_2[9:0];
                output_real_0_3_pipe <= config0_3[19:10];
                output_imag_0_3_pipe <= config0_3[9:0];
                output_real_1_3_pipe <= config1_3[19:10];
                output_imag_1_3_pipe <= config1_3[9:0];
                output_real_2_3_pipe <= config2_3[19:10];
                output_imag_2_3_pipe <= config2_3[9:0];
                output_real_3_3_pipe <= config3_3[19:10];
                output_imag_3_3_pipe <= config3_3[9:0];
                output_real_4_3_pipe <= config4_3[19:10];
                output_imag_4_3_pipe <= config4_3[9:0];
                output_real_5_3_pipe <= config5_3[19:10];
                output_imag_5_3_pipe <= config5_3[9:0];
                output_real_6_3_pipe <= config6_3[19:10];
                output_imag_6_3_pipe <= config6_3[9:0];
                output_real_7_3_pipe <= config7_3[19:10];
                output_imag_7_3_pipe <= config7_3[9:0];
                output_real_8_3_pipe <= config8_3[19:10];
                output_imag_8_3_pipe <= config8_3[9:0];
                output_real_9_3_pipe <= config9_3[19:10];
                output_imag_9_3_pipe <= config9_3[9:0];
                output_real_10_3_pipe <= config10_3[19:10];
                output_imag_10_3_pipe <= config10_3[9:0];
                output_real_11_3_pipe <= config11_3[19:10];
                output_imag_11_3_pipe <= config11_3[9:0];
                output_real_12_3_pipe <= config12_3[19:10];
                output_imag_12_3_pipe <= config12_3[9:0];
                output_real_13_3_pipe <= config13_3[19:10];
                output_imag_13_3_pipe <= config13_3[9:0];
                output_real_14_3_pipe <= config14_3[19:10];
                output_imag_14_3_pipe <= config14_3[9:0];
                output_real_15_3_pipe <= config15_3[19:10];
                output_imag_15_3_pipe <= config15_3[9:0];
                output_real_16_3_pipe <= config16_3[19:10];
                output_imag_16_3_pipe <= config16_3[9:0];
                output_real_17_3_pipe <= config17_3[19:10];
                output_imag_17_3_pipe <= config17_3[9:0];
                output_real_18_3_pipe <= config18_3[19:10];
                output_imag_18_3_pipe <= config18_3[9:0];
                output_real_19_3_pipe <= config19_3[19:10];
                output_imag_19_3_pipe <= config19_3[9:0];
                output_real_20_3_pipe <= config20_3[19:10];
                output_imag_20_3_pipe <= config20_3[9:0];
                output_real_21_3_pipe <= config21_3[19:10];
                output_imag_21_3_pipe <= config21_3[9:0];
                output_real_22_3_pipe <= config22_3[19:10];
                output_imag_22_3_pipe <= config22_3[9:0];
                output_real_23_3_pipe <= config23_3[19:10];
                output_imag_23_3_pipe <= config23_3[9:0];
                output_real_24_3_pipe <= config24_3[19:10];
                output_imag_24_3_pipe <= config24_3[9:0];
                output_real_25_3_pipe <= config25_3[19:10];
                output_imag_25_3_pipe <= config25_3[9:0];
                output_real_26_3_pipe <= config26_3[19:10];
                output_imag_26_3_pipe <= config26_3[9:0];
                output_real_27_3_pipe <= config27_3[19:10];
                output_imag_27_3_pipe <= config27_3[9:0];
                output_real_28_3_pipe <= config28_3[19:10];
                output_imag_28_3_pipe <= config28_3[9:0];
                output_real_29_3_pipe <= config29_3[19:10];
                output_imag_29_3_pipe <= config29_3[9:0];
                output_real_30_3_pipe <= config30_3[19:10];
                output_imag_30_3_pipe <= config30_3[9:0];
                output_real_31_3_pipe <= config31_3[19:10];
                output_imag_31_3_pipe <= config31_3[9:0];
                output_real_32_3_pipe <= config32_3[19:10];
                output_imag_32_3_pipe <= config32_3[9:0];
                output_real_33_3_pipe <= config33_3[19:10];
                output_imag_33_3_pipe <= config33_3[9:0];
                output_real_34_3_pipe <= config34_3[19:10];
                output_imag_34_3_pipe <= config34_3[9:0];
                output_real_35_3_pipe <= config35_3[19:10];
                output_imag_35_3_pipe <= config35_3[9:0];
                output_real_36_3_pipe <= config36_3[19:10];
                output_imag_36_3_pipe <= config36_3[9:0];
                output_real_37_3_pipe <= config37_3[19:10];
                output_imag_37_3_pipe <= config37_3[9:0];
                output_real_38_3_pipe <= config38_3[19:10];
                output_imag_38_3_pipe <= config38_3[9:0];
                output_real_39_3_pipe <= config39_3[19:10];
                output_imag_39_3_pipe <= config39_3[9:0];
                output_real_40_3_pipe <= config40_3[19:10];
                output_imag_40_3_pipe <= config40_3[9:0];
                output_real_41_3_pipe <= config41_3[19:10];
                output_imag_41_3_pipe <= config41_3[9:0];
                output_real_42_3_pipe <= config42_3[19:10];
                output_imag_42_3_pipe <= config42_3[9:0];
                output_real_43_3_pipe <= config43_3[19:10];
                output_imag_43_3_pipe <= config43_3[9:0];
                output_real_44_3_pipe <= config44_3[19:10];
                output_imag_44_3_pipe <= config44_3[9:0];
                output_real_45_3_pipe <= config45_3[19:10];
                output_imag_45_3_pipe <= config45_3[9:0];
                output_real_46_3_pipe <= config46_3[19:10];
                output_imag_46_3_pipe <= config46_3[9:0];
                output_real_47_3_pipe <= config47_3[19:10];
                output_imag_47_3_pipe <= config47_3[9:0];
                output_real_48_3_pipe <= config48_3[19:10];
                output_imag_48_3_pipe <= config48_3[9:0];
                output_real_49_3_pipe <= config49_3[19:10];
                output_imag_49_3_pipe <= config49_3[9:0];
                output_real_50_3_pipe <= config50_3[19:10];
                output_imag_50_3_pipe <= config50_3[9:0];
                output_real_51_3_pipe <= config51_3[19:10];
                output_imag_51_3_pipe <= config51_3[9:0];
                output_real_52_3_pipe <= config52_3[19:10];
                output_imag_52_3_pipe <= config52_3[9:0];
                output_real_53_3_pipe <= config53_3[19:10];
                output_imag_53_3_pipe <= config53_3[9:0];
                output_real_54_3_pipe <= config54_3[19:10];
                output_imag_54_3_pipe <= config54_3[9:0];
                output_real_55_3_pipe <= config55_3[19:10];
                output_imag_55_3_pipe <= config55_3[9:0];
                output_real_56_3_pipe <= config56_3[19:10];
                output_imag_56_3_pipe <= config56_3[9:0];
                output_real_57_3_pipe <= config57_3[19:10];
                output_imag_57_3_pipe <= config57_3[9:0];
                output_real_58_3_pipe <= config58_3[19:10];
                output_imag_58_3_pipe <= config58_3[9:0];
                output_real_59_3_pipe <= config59_3[19:10];
                output_imag_59_3_pipe <= config59_3[9:0];
                output_real_60_3_pipe <= config60_3[19:10];
                output_imag_60_3_pipe <= config60_3[9:0];
                output_real_61_3_pipe <= config61_3[19:10];
                output_imag_61_3_pipe <= config61_3[9:0];
                output_real_62_3_pipe <= config62_3[19:10];
                output_imag_62_3_pipe <= config62_3[9:0];
                output_real_63_3_pipe <= config63_3[19:10];
                output_imag_63_3_pipe <= config63_3[9:0];

        end
        else begin
		output_real_0_0_pipe <= output_real_0_0_pipe;
                output_imag_0_0_pipe <= output_imag_0_0_pipe;
		output_real_1_0_pipe <= output_real_1_0_pipe;
                output_imag_1_0_pipe <= output_imag_1_0_pipe;
		output_real_2_0_pipe <= output_real_2_0_pipe;
                output_imag_2_0_pipe <= output_imag_2_0_pipe;
		output_real_3_0_pipe <= output_real_3_0_pipe;
                output_imag_3_0_pipe <= output_imag_3_0_pipe;
		output_real_4_0_pipe <= output_real_4_0_pipe;
                output_imag_4_0_pipe <= output_imag_4_0_pipe;
		output_real_5_0_pipe <= output_real_5_0_pipe;
                output_imag_5_0_pipe <= output_imag_5_0_pipe;
		output_real_6_0_pipe <= output_real_6_0_pipe;
                output_imag_6_0_pipe <= output_imag_6_0_pipe;
		output_real_7_0_pipe <= output_real_7_0_pipe;
                output_imag_7_0_pipe <= output_imag_7_0_pipe;
		output_real_8_0_pipe <= output_real_8_0_pipe;
                output_imag_8_0_pipe <= output_imag_8_0_pipe;
		output_real_9_0_pipe <= output_real_9_0_pipe;
                output_imag_9_0_pipe <= output_imag_9_0_pipe;
		output_real_10_0_pipe <= output_real_10_0_pipe;
                output_imag_10_0_pipe <= output_imag_10_0_pipe;
		output_real_11_0_pipe <= output_real_11_0_pipe;
                output_imag_11_0_pipe <= output_imag_11_0_pipe;
		output_real_12_0_pipe <= output_real_12_0_pipe;
                output_imag_12_0_pipe <= output_imag_12_0_pipe;
		output_real_13_0_pipe <= output_real_13_0_pipe;
                output_imag_13_0_pipe <= output_imag_13_0_pipe;
		output_real_14_0_pipe <= output_real_14_0_pipe;
                output_imag_14_0_pipe <= output_imag_14_0_pipe;
		output_real_15_0_pipe <= output_real_15_0_pipe;
                output_imag_15_0_pipe <= output_imag_15_0_pipe;
		output_real_16_0_pipe <= output_real_16_0_pipe;
                output_imag_16_0_pipe <= output_imag_16_0_pipe;
		output_real_17_0_pipe <= output_real_17_0_pipe;
                output_imag_17_0_pipe <= output_imag_17_0_pipe;
		output_real_18_0_pipe <= output_real_18_0_pipe;
                output_imag_18_0_pipe <= output_imag_18_0_pipe;
		output_real_19_0_pipe <= output_real_19_0_pipe;
                output_imag_19_0_pipe <= output_imag_19_0_pipe;
		output_real_20_0_pipe <= output_real_20_0_pipe;
                output_imag_20_0_pipe <= output_imag_20_0_pipe;
		output_real_21_0_pipe <= output_real_21_0_pipe;
                output_imag_21_0_pipe <= output_imag_21_0_pipe;
		output_real_22_0_pipe <= output_real_22_0_pipe;
                output_imag_22_0_pipe <= output_imag_22_0_pipe;
		output_real_23_0_pipe <= output_real_23_0_pipe;
                output_imag_23_0_pipe <= output_imag_23_0_pipe;
		output_real_24_0_pipe <= output_real_24_0_pipe;
                output_imag_24_0_pipe <= output_imag_24_0_pipe;
		output_real_25_0_pipe <= output_real_25_0_pipe;
                output_imag_25_0_pipe <= output_imag_25_0_pipe;
		output_real_26_0_pipe <= output_real_26_0_pipe;
                output_imag_26_0_pipe <= output_imag_26_0_pipe;
		output_real_27_0_pipe <= output_real_27_0_pipe;
                output_imag_27_0_pipe <= output_imag_27_0_pipe;
		output_real_28_0_pipe <= output_real_28_0_pipe;
                output_imag_28_0_pipe <= output_imag_28_0_pipe;
		output_real_29_0_pipe <= output_real_29_0_pipe;
                output_imag_29_0_pipe <= output_imag_29_0_pipe;
		output_real_30_0_pipe <= output_real_30_0_pipe;
                output_imag_30_0_pipe <= output_imag_30_0_pipe;
		output_real_31_0_pipe <= output_real_31_0_pipe;
                output_imag_31_0_pipe <= output_imag_31_0_pipe;
		output_real_32_0_pipe <= output_real_32_0_pipe;
                output_imag_32_0_pipe <= output_imag_32_0_pipe;
		output_real_33_0_pipe <= output_real_33_0_pipe;
                output_imag_33_0_pipe <= output_imag_33_0_pipe;
		output_real_34_0_pipe <= output_real_34_0_pipe;
                output_imag_34_0_pipe <= output_imag_34_0_pipe;
		output_real_35_0_pipe <= output_real_35_0_pipe;
                output_imag_35_0_pipe <= output_imag_35_0_pipe;
		output_real_36_0_pipe <= output_real_36_0_pipe;
                output_imag_36_0_pipe <= output_imag_36_0_pipe;
		output_real_37_0_pipe <= output_real_37_0_pipe;
                output_imag_37_0_pipe <= output_imag_37_0_pipe;
		output_real_38_0_pipe <= output_real_38_0_pipe;
                output_imag_38_0_pipe <= output_imag_38_0_pipe;
		output_real_39_0_pipe <= output_real_39_0_pipe;
                output_imag_39_0_pipe <= output_imag_39_0_pipe;
		output_real_40_0_pipe <= output_real_40_0_pipe;
                output_imag_40_0_pipe <= output_imag_40_0_pipe;
		output_real_41_0_pipe <= output_real_41_0_pipe;
                output_imag_41_0_pipe <= output_imag_41_0_pipe;
		output_real_42_0_pipe <= output_real_42_0_pipe;
                output_imag_42_0_pipe <= output_imag_42_0_pipe;
		output_real_43_0_pipe <= output_real_43_0_pipe;
                output_imag_43_0_pipe <= output_imag_43_0_pipe;
		output_real_44_0_pipe <= output_real_44_0_pipe;
                output_imag_44_0_pipe <= output_imag_44_0_pipe;
		output_real_45_0_pipe <= output_real_45_0_pipe;
                output_imag_45_0_pipe <= output_imag_45_0_pipe;
		output_real_46_0_pipe <= output_real_46_0_pipe;
                output_imag_46_0_pipe <= output_imag_46_0_pipe;
		output_real_47_0_pipe <= output_real_47_0_pipe;
                output_imag_47_0_pipe <= output_imag_47_0_pipe;
		output_real_48_0_pipe <= output_real_48_0_pipe;
                output_imag_48_0_pipe <= output_imag_48_0_pipe;
		output_real_49_0_pipe <= output_real_49_0_pipe;
                output_imag_49_0_pipe <= output_imag_49_0_pipe;
		output_real_50_0_pipe <= output_real_50_0_pipe;
                output_imag_50_0_pipe <= output_imag_50_0_pipe;
		output_real_51_0_pipe <= output_real_51_0_pipe;
                output_imag_51_0_pipe <= output_imag_51_0_pipe;
		output_real_52_0_pipe <= output_real_52_0_pipe;
                output_imag_52_0_pipe <= output_imag_52_0_pipe;
		output_real_53_0_pipe <= output_real_53_0_pipe;
                output_imag_53_0_pipe <= output_imag_53_0_pipe;
		output_real_54_0_pipe <= output_real_54_0_pipe;
                output_imag_54_0_pipe <= output_imag_54_0_pipe;
		output_real_55_0_pipe <= output_real_55_0_pipe;
                output_imag_55_0_pipe <= output_imag_55_0_pipe;
		output_real_56_0_pipe <= output_real_56_0_pipe;
                output_imag_56_0_pipe <= output_imag_56_0_pipe;
		output_real_57_0_pipe <= output_real_57_0_pipe;
                output_imag_57_0_pipe <= output_imag_57_0_pipe;
		output_real_58_0_pipe <= output_real_58_0_pipe;
                output_imag_58_0_pipe <= output_imag_58_0_pipe;
		output_real_59_0_pipe <= output_real_59_0_pipe;
                output_imag_59_0_pipe <= output_imag_59_0_pipe;
		output_real_60_0_pipe <= output_real_60_0_pipe;
                output_imag_60_0_pipe <= output_imag_60_0_pipe;
		output_real_61_0_pipe <= output_real_61_0_pipe;
                output_imag_61_0_pipe <= output_imag_61_0_pipe;
		output_real_62_0_pipe <= output_real_62_0_pipe;
                output_imag_62_0_pipe <= output_imag_62_0_pipe;
		output_real_63_0_pipe <= output_real_63_0_pipe;
                output_imag_63_0_pipe <= output_imag_63_0_pipe;
		output_real_0_1_pipe <= output_real_0_1_pipe;
                output_imag_0_1_pipe <= output_imag_0_1_pipe;
		output_real_1_1_pipe <= output_real_1_1_pipe;
                output_imag_1_1_pipe <= output_imag_1_1_pipe;
		output_real_2_1_pipe <= output_real_2_1_pipe;
                output_imag_2_1_pipe <= output_imag_2_1_pipe;
		output_real_3_1_pipe <= output_real_3_1_pipe;
                output_imag_3_1_pipe <= output_imag_3_1_pipe;
		output_real_4_1_pipe <= output_real_4_1_pipe;
                output_imag_4_1_pipe <= output_imag_4_1_pipe;
		output_real_5_1_pipe <= output_real_5_1_pipe;
                output_imag_5_1_pipe <= output_imag_5_1_pipe;
		output_real_6_1_pipe <= output_real_6_1_pipe;
                output_imag_6_1_pipe <= output_imag_6_1_pipe;
		output_real_7_1_pipe <= output_real_7_1_pipe;
                output_imag_7_1_pipe <= output_imag_7_1_pipe;
		output_real_8_1_pipe <= output_real_8_1_pipe;
                output_imag_8_1_pipe <= output_imag_8_1_pipe;
		output_real_9_1_pipe <= output_real_9_1_pipe;
                output_imag_9_1_pipe <= output_imag_9_1_pipe;
		output_real_10_1_pipe <= output_real_10_1_pipe;
                output_imag_10_1_pipe <= output_imag_10_1_pipe;
		output_real_11_1_pipe <= output_real_11_1_pipe;
                output_imag_11_1_pipe <= output_imag_11_1_pipe;
		output_real_12_1_pipe <= output_real_12_1_pipe;
                output_imag_12_1_pipe <= output_imag_12_1_pipe;
		output_real_13_1_pipe <= output_real_13_1_pipe;
                output_imag_13_1_pipe <= output_imag_13_1_pipe;
		output_real_14_1_pipe <= output_real_14_1_pipe;
                output_imag_14_1_pipe <= output_imag_14_1_pipe;
		output_real_15_1_pipe <= output_real_15_1_pipe;
                output_imag_15_1_pipe <= output_imag_15_1_pipe;
		output_real_16_1_pipe <= output_real_16_1_pipe;
                output_imag_16_1_pipe <= output_imag_16_1_pipe;
		output_real_17_1_pipe <= output_real_17_1_pipe;
                output_imag_17_1_pipe <= output_imag_17_1_pipe;
		output_real_18_1_pipe <= output_real_18_1_pipe;
                output_imag_18_1_pipe <= output_imag_18_1_pipe;
		output_real_19_1_pipe <= output_real_19_1_pipe;
                output_imag_19_1_pipe <= output_imag_19_1_pipe;
		output_real_20_1_pipe <= output_real_20_1_pipe;
                output_imag_20_1_pipe <= output_imag_20_1_pipe;
		output_real_21_1_pipe <= output_real_21_1_pipe;
                output_imag_21_1_pipe <= output_imag_21_1_pipe;
		output_real_22_1_pipe <= output_real_22_1_pipe;
                output_imag_22_1_pipe <= output_imag_22_1_pipe;
		output_real_23_1_pipe <= output_real_23_1_pipe;
                output_imag_23_1_pipe <= output_imag_23_1_pipe;
		output_real_24_1_pipe <= output_real_24_1_pipe;
                output_imag_24_1_pipe <= output_imag_24_1_pipe;
		output_real_25_1_pipe <= output_real_25_1_pipe;
                output_imag_25_1_pipe <= output_imag_25_1_pipe;
		output_real_26_1_pipe <= output_real_26_1_pipe;
                output_imag_26_1_pipe <= output_imag_26_1_pipe;
		output_real_27_1_pipe <= output_real_27_1_pipe;
                output_imag_27_1_pipe <= output_imag_27_1_pipe;
		output_real_28_1_pipe <= output_real_28_1_pipe;
                output_imag_28_1_pipe <= output_imag_28_1_pipe;
		output_real_29_1_pipe <= output_real_29_1_pipe;
                output_imag_29_1_pipe <= output_imag_29_1_pipe;
		output_real_30_1_pipe <= output_real_30_1_pipe;
                output_imag_30_1_pipe <= output_imag_30_1_pipe;
		output_real_31_1_pipe <= output_real_31_1_pipe;
                output_imag_31_1_pipe <= output_imag_31_1_pipe;
		output_real_32_1_pipe <= output_real_32_1_pipe;
                output_imag_32_1_pipe <= output_imag_32_1_pipe;
		output_real_33_1_pipe <= output_real_33_1_pipe;
                output_imag_33_1_pipe <= output_imag_33_1_pipe;
		output_real_34_1_pipe <= output_real_34_1_pipe;
                output_imag_34_1_pipe <= output_imag_34_1_pipe;
		output_real_35_1_pipe <= output_real_35_1_pipe;
                output_imag_35_1_pipe <= output_imag_35_1_pipe;
		output_real_36_1_pipe <= output_real_36_1_pipe;
                output_imag_36_1_pipe <= output_imag_36_1_pipe;
		output_real_37_1_pipe <= output_real_37_1_pipe;
                output_imag_37_1_pipe <= output_imag_37_1_pipe;
		output_real_38_1_pipe <= output_real_38_1_pipe;
                output_imag_38_1_pipe <= output_imag_38_1_pipe;
		output_real_39_1_pipe <= output_real_39_1_pipe;
                output_imag_39_1_pipe <= output_imag_39_1_pipe;
		output_real_40_1_pipe <= output_real_40_1_pipe;
                output_imag_40_1_pipe <= output_imag_40_1_pipe;
		output_real_41_1_pipe <= output_real_41_1_pipe;
                output_imag_41_1_pipe <= output_imag_41_1_pipe;
		output_real_42_1_pipe <= output_real_42_1_pipe;
                output_imag_42_1_pipe <= output_imag_42_1_pipe;
		output_real_43_1_pipe <= output_real_43_1_pipe;
                output_imag_43_1_pipe <= output_imag_43_1_pipe;
		output_real_44_1_pipe <= output_real_44_1_pipe;
                output_imag_44_1_pipe <= output_imag_44_1_pipe;
		output_real_45_1_pipe <= output_real_45_1_pipe;
                output_imag_45_1_pipe <= output_imag_45_1_pipe;
		output_real_46_1_pipe <= output_real_46_1_pipe;
                output_imag_46_1_pipe <= output_imag_46_1_pipe;
		output_real_47_1_pipe <= output_real_47_1_pipe;
                output_imag_47_1_pipe <= output_imag_47_1_pipe;
		output_real_48_1_pipe <= output_real_48_1_pipe;
                output_imag_48_1_pipe <= output_imag_48_1_pipe;
		output_real_49_1_pipe <= output_real_49_1_pipe;
                output_imag_49_1_pipe <= output_imag_49_1_pipe;
		output_real_50_1_pipe <= output_real_50_1_pipe;
                output_imag_50_1_pipe <= output_imag_50_1_pipe;
		output_real_51_1_pipe <= output_real_51_1_pipe;
                output_imag_51_1_pipe <= output_imag_51_1_pipe;
		output_real_52_1_pipe <= output_real_52_1_pipe;
                output_imag_52_1_pipe <= output_imag_52_1_pipe;
		output_real_53_1_pipe <= output_real_53_1_pipe;
                output_imag_53_1_pipe <= output_imag_53_1_pipe;
		output_real_54_1_pipe <= output_real_54_1_pipe;
                output_imag_54_1_pipe <= output_imag_54_1_pipe;
		output_real_55_1_pipe <= output_real_55_1_pipe;
                output_imag_55_1_pipe <= output_imag_55_1_pipe;
		output_real_56_1_pipe <= output_real_56_1_pipe;
                output_imag_56_1_pipe <= output_imag_56_1_pipe;
		output_real_57_1_pipe <= output_real_57_1_pipe;
                output_imag_57_1_pipe <= output_imag_57_1_pipe;
		output_real_58_1_pipe <= output_real_58_1_pipe;
                output_imag_58_1_pipe <= output_imag_58_1_pipe;
		output_real_59_1_pipe <= output_real_59_1_pipe;
                output_imag_59_1_pipe <= output_imag_59_1_pipe;
		output_real_60_1_pipe <= output_real_60_1_pipe;
                output_imag_60_1_pipe <= output_imag_60_1_pipe;
		output_real_61_1_pipe <= output_real_61_1_pipe;
                output_imag_61_1_pipe <= output_imag_61_1_pipe;
		output_real_62_1_pipe <= output_real_62_1_pipe;
                output_imag_62_1_pipe <= output_imag_62_1_pipe;
		output_real_63_1_pipe <= output_real_63_1_pipe;
                output_imag_63_1_pipe <= output_imag_63_1_pipe;
		output_real_0_2_pipe <= output_real_0_2_pipe;
                output_imag_0_2_pipe <= output_imag_0_2_pipe;
		output_real_1_2_pipe <= output_real_1_2_pipe;
                output_imag_1_2_pipe <= output_imag_1_2_pipe;
		output_real_2_2_pipe <= output_real_2_2_pipe;
                output_imag_2_2_pipe <= output_imag_2_2_pipe;
		output_real_3_2_pipe <= output_real_3_2_pipe;
                output_imag_3_2_pipe <= output_imag_3_2_pipe;
		output_real_4_2_pipe <= output_real_4_2_pipe;
                output_imag_4_2_pipe <= output_imag_4_2_pipe;
		output_real_5_2_pipe <= output_real_5_2_pipe;
                output_imag_5_2_pipe <= output_imag_5_2_pipe;
		output_real_6_2_pipe <= output_real_6_2_pipe;
                output_imag_6_2_pipe <= output_imag_6_2_pipe;
		output_real_7_2_pipe <= output_real_7_2_pipe;
                output_imag_7_2_pipe <= output_imag_7_2_pipe;
		output_real_8_2_pipe <= output_real_8_2_pipe;
                output_imag_8_2_pipe <= output_imag_8_2_pipe;
		output_real_9_2_pipe <= output_real_9_2_pipe;
                output_imag_9_2_pipe <= output_imag_9_2_pipe;
		output_real_10_2_pipe <= output_real_10_2_pipe;
                output_imag_10_2_pipe <= output_imag_10_2_pipe;
		output_real_11_2_pipe <= output_real_11_2_pipe;
                output_imag_11_2_pipe <= output_imag_11_2_pipe;
		output_real_12_2_pipe <= output_real_12_2_pipe;
                output_imag_12_2_pipe <= output_imag_12_2_pipe;
		output_real_13_2_pipe <= output_real_13_2_pipe;
                output_imag_13_2_pipe <= output_imag_13_2_pipe;
		output_real_14_2_pipe <= output_real_14_2_pipe;
                output_imag_14_2_pipe <= output_imag_14_2_pipe;
		output_real_15_2_pipe <= output_real_15_2_pipe;
                output_imag_15_2_pipe <= output_imag_15_2_pipe;
		output_real_16_2_pipe <= output_real_16_2_pipe;
                output_imag_16_2_pipe <= output_imag_16_2_pipe;
		output_real_17_2_pipe <= output_real_17_2_pipe;
                output_imag_17_2_pipe <= output_imag_17_2_pipe;
		output_real_18_2_pipe <= output_real_18_2_pipe;
                output_imag_18_2_pipe <= output_imag_18_2_pipe;
		output_real_19_2_pipe <= output_real_19_2_pipe;
                output_imag_19_2_pipe <= output_imag_19_2_pipe;
		output_real_20_2_pipe <= output_real_20_2_pipe;
                output_imag_20_2_pipe <= output_imag_20_2_pipe;
		output_real_21_2_pipe <= output_real_21_2_pipe;
                output_imag_21_2_pipe <= output_imag_21_2_pipe;
		output_real_22_2_pipe <= output_real_22_2_pipe;
                output_imag_22_2_pipe <= output_imag_22_2_pipe;
		output_real_23_2_pipe <= output_real_23_2_pipe;
                output_imag_23_2_pipe <= output_imag_23_2_pipe;
		output_real_24_2_pipe <= output_real_24_2_pipe;
                output_imag_24_2_pipe <= output_imag_24_2_pipe;
		output_real_25_2_pipe <= output_real_25_2_pipe;
                output_imag_25_2_pipe <= output_imag_25_2_pipe;
		output_real_26_2_pipe <= output_real_26_2_pipe;
                output_imag_26_2_pipe <= output_imag_26_2_pipe;
		output_real_27_2_pipe <= output_real_27_2_pipe;
                output_imag_27_2_pipe <= output_imag_27_2_pipe;
		output_real_28_2_pipe <= output_real_28_2_pipe;
                output_imag_28_2_pipe <= output_imag_28_2_pipe;
		output_real_29_2_pipe <= output_real_29_2_pipe;
                output_imag_29_2_pipe <= output_imag_29_2_pipe;
		output_real_30_2_pipe <= output_real_30_2_pipe;
                output_imag_30_2_pipe <= output_imag_30_2_pipe;
		output_real_31_2_pipe <= output_real_31_2_pipe;
                output_imag_31_2_pipe <= output_imag_31_2_pipe;
		output_real_32_2_pipe <= output_real_32_2_pipe;
                output_imag_32_2_pipe <= output_imag_32_2_pipe;
		output_real_33_2_pipe <= output_real_33_2_pipe;
                output_imag_33_2_pipe <= output_imag_33_2_pipe;
		output_real_34_2_pipe <= output_real_34_2_pipe;
                output_imag_34_2_pipe <= output_imag_34_2_pipe;
		output_real_35_2_pipe <= output_real_35_2_pipe;
                output_imag_35_2_pipe <= output_imag_35_2_pipe;
		output_real_36_2_pipe <= output_real_36_2_pipe;
                output_imag_36_2_pipe <= output_imag_36_2_pipe;
		output_real_37_2_pipe <= output_real_37_2_pipe;
                output_imag_37_2_pipe <= output_imag_37_2_pipe;
		output_real_38_2_pipe <= output_real_38_2_pipe;
                output_imag_38_2_pipe <= output_imag_38_2_pipe;
		output_real_39_2_pipe <= output_real_39_2_pipe;
                output_imag_39_2_pipe <= output_imag_39_2_pipe;
		output_real_40_2_pipe <= output_real_40_2_pipe;
                output_imag_40_2_pipe <= output_imag_40_2_pipe;
		output_real_41_2_pipe <= output_real_41_2_pipe;
                output_imag_41_2_pipe <= output_imag_41_2_pipe;
		output_real_42_2_pipe <= output_real_42_2_pipe;
                output_imag_42_2_pipe <= output_imag_42_2_pipe;
		output_real_43_2_pipe <= output_real_43_2_pipe;
                output_imag_43_2_pipe <= output_imag_43_2_pipe;
		output_real_44_2_pipe <= output_real_44_2_pipe;
                output_imag_44_2_pipe <= output_imag_44_2_pipe;
		output_real_45_2_pipe <= output_real_45_2_pipe;
                output_imag_45_2_pipe <= output_imag_45_2_pipe;
		output_real_46_2_pipe <= output_real_46_2_pipe;
                output_imag_46_2_pipe <= output_imag_46_2_pipe;
		output_real_47_2_pipe <= output_real_47_2_pipe;
                output_imag_47_2_pipe <= output_imag_47_2_pipe;
		output_real_48_2_pipe <= output_real_48_2_pipe;
                output_imag_48_2_pipe <= output_imag_48_2_pipe;
		output_real_49_2_pipe <= output_real_49_2_pipe;
                output_imag_49_2_pipe <= output_imag_49_2_pipe;
		output_real_50_2_pipe <= output_real_50_2_pipe;
                output_imag_50_2_pipe <= output_imag_50_2_pipe;
		output_real_51_2_pipe <= output_real_51_2_pipe;
                output_imag_51_2_pipe <= output_imag_51_2_pipe;
		output_real_52_2_pipe <= output_real_52_2_pipe;
                output_imag_52_2_pipe <= output_imag_52_2_pipe;
		output_real_53_2_pipe <= output_real_53_2_pipe;
                output_imag_53_2_pipe <= output_imag_53_2_pipe;
		output_real_54_2_pipe <= output_real_54_2_pipe;
                output_imag_54_2_pipe <= output_imag_54_2_pipe;
		output_real_55_2_pipe <= output_real_55_2_pipe;
                output_imag_55_2_pipe <= output_imag_55_2_pipe;
		output_real_56_2_pipe <= output_real_56_2_pipe;
                output_imag_56_2_pipe <= output_imag_56_2_pipe;
		output_real_57_2_pipe <= output_real_57_2_pipe;
                output_imag_57_2_pipe <= output_imag_57_2_pipe;
		output_real_58_2_pipe <= output_real_58_2_pipe;
                output_imag_58_2_pipe <= output_imag_58_2_pipe;
		output_real_59_2_pipe <= output_real_59_2_pipe;
                output_imag_59_2_pipe <= output_imag_59_2_pipe;
		output_real_60_2_pipe <= output_real_60_2_pipe;
                output_imag_60_2_pipe <= output_imag_60_2_pipe;
		output_real_61_2_pipe <= output_real_61_2_pipe;
                output_imag_61_2_pipe <= output_imag_61_2_pipe;
		output_real_62_2_pipe <= output_real_62_2_pipe;
                output_imag_62_2_pipe <= output_imag_62_2_pipe;
		output_real_63_2_pipe <= output_real_63_2_pipe;
                output_imag_63_2_pipe <= output_imag_63_2_pipe;
		output_real_0_3_pipe <= output_real_0_3_pipe;
                output_imag_0_3_pipe <= output_imag_0_3_pipe;
		output_real_1_3_pipe <= output_real_1_3_pipe;
                output_imag_1_3_pipe <= output_imag_1_3_pipe;
		output_real_2_3_pipe <= output_real_2_3_pipe;
                output_imag_2_3_pipe <= output_imag_2_3_pipe;
		output_real_3_3_pipe <= output_real_3_3_pipe;
                output_imag_3_3_pipe <= output_imag_3_3_pipe;
		output_real_4_3_pipe <= output_real_4_3_pipe;
                output_imag_4_3_pipe <= output_imag_4_3_pipe;
		output_real_5_3_pipe <= output_real_5_3_pipe;
                output_imag_5_3_pipe <= output_imag_5_3_pipe;
		output_real_6_3_pipe <= output_real_6_3_pipe;
                output_imag_6_3_pipe <= output_imag_6_3_pipe;
		output_real_7_3_pipe <= output_real_7_3_pipe;
                output_imag_7_3_pipe <= output_imag_7_3_pipe;
		output_real_8_3_pipe <= output_real_8_3_pipe;
                output_imag_8_3_pipe <= output_imag_8_3_pipe;
		output_real_9_3_pipe <= output_real_9_3_pipe;
                output_imag_9_3_pipe <= output_imag_9_3_pipe;
		output_real_10_3_pipe <= output_real_10_3_pipe;
                output_imag_10_3_pipe <= output_imag_10_3_pipe;
		output_real_11_3_pipe <= output_real_11_3_pipe;
                output_imag_11_3_pipe <= output_imag_11_3_pipe;
		output_real_12_3_pipe <= output_real_12_3_pipe;
                output_imag_12_3_pipe <= output_imag_12_3_pipe;
		output_real_13_3_pipe <= output_real_13_3_pipe;
                output_imag_13_3_pipe <= output_imag_13_3_pipe;
		output_real_14_3_pipe <= output_real_14_3_pipe;
                output_imag_14_3_pipe <= output_imag_14_3_pipe;
		output_real_15_3_pipe <= output_real_15_3_pipe;
                output_imag_15_3_pipe <= output_imag_15_3_pipe;
		output_real_16_3_pipe <= output_real_16_3_pipe;
                output_imag_16_3_pipe <= output_imag_16_3_pipe;
		output_real_17_3_pipe <= output_real_17_3_pipe;
                output_imag_17_3_pipe <= output_imag_17_3_pipe;
		output_real_18_3_pipe <= output_real_18_3_pipe;
                output_imag_18_3_pipe <= output_imag_18_3_pipe;
		output_real_19_3_pipe <= output_real_19_3_pipe;
                output_imag_19_3_pipe <= output_imag_19_3_pipe;
		output_real_20_3_pipe <= output_real_20_3_pipe;
                output_imag_20_3_pipe <= output_imag_20_3_pipe;
		output_real_21_3_pipe <= output_real_21_3_pipe;
                output_imag_21_3_pipe <= output_imag_21_3_pipe;
		output_real_22_3_pipe <= output_real_22_3_pipe;
                output_imag_22_3_pipe <= output_imag_22_3_pipe;
		output_real_23_3_pipe <= output_real_23_3_pipe;
                output_imag_23_3_pipe <= output_imag_23_3_pipe;
		output_real_24_3_pipe <= output_real_24_3_pipe;
                output_imag_24_3_pipe <= output_imag_24_3_pipe;
		output_real_25_3_pipe <= output_real_25_3_pipe;
                output_imag_25_3_pipe <= output_imag_25_3_pipe;
		output_real_26_3_pipe <= output_real_26_3_pipe;
                output_imag_26_3_pipe <= output_imag_26_3_pipe;
		output_real_27_3_pipe <= output_real_27_3_pipe;
                output_imag_27_3_pipe <= output_imag_27_3_pipe;
		output_real_28_3_pipe <= output_real_28_3_pipe;
                output_imag_28_3_pipe <= output_imag_28_3_pipe;
		output_real_29_3_pipe <= output_real_29_3_pipe;
                output_imag_29_3_pipe <= output_imag_29_3_pipe;
		output_real_30_3_pipe <= output_real_30_3_pipe;
                output_imag_30_3_pipe <= output_imag_30_3_pipe;
		output_real_31_3_pipe <= output_real_31_3_pipe;
                output_imag_31_3_pipe <= output_imag_31_3_pipe;
		output_real_32_3_pipe <= output_real_32_3_pipe;
                output_imag_32_3_pipe <= output_imag_32_3_pipe;
		output_real_33_3_pipe <= output_real_33_3_pipe;
                output_imag_33_3_pipe <= output_imag_33_3_pipe;
		output_real_34_3_pipe <= output_real_34_3_pipe;
                output_imag_34_3_pipe <= output_imag_34_3_pipe;
		output_real_35_3_pipe <= output_real_35_3_pipe;
                output_imag_35_3_pipe <= output_imag_35_3_pipe;
		output_real_36_3_pipe <= output_real_36_3_pipe;
                output_imag_36_3_pipe <= output_imag_36_3_pipe;
		output_real_37_3_pipe <= output_real_37_3_pipe;
                output_imag_37_3_pipe <= output_imag_37_3_pipe;
		output_real_38_3_pipe <= output_real_38_3_pipe;
                output_imag_38_3_pipe <= output_imag_38_3_pipe;
		output_real_39_3_pipe <= output_real_39_3_pipe;
                output_imag_39_3_pipe <= output_imag_39_3_pipe;
		output_real_40_3_pipe <= output_real_40_3_pipe;
                output_imag_40_3_pipe <= output_imag_40_3_pipe;
		output_real_41_3_pipe <= output_real_41_3_pipe;
                output_imag_41_3_pipe <= output_imag_41_3_pipe;
		output_real_42_3_pipe <= output_real_42_3_pipe;
                output_imag_42_3_pipe <= output_imag_42_3_pipe;
		output_real_43_3_pipe <= output_real_43_3_pipe;
                output_imag_43_3_pipe <= output_imag_43_3_pipe;
		output_real_44_3_pipe <= output_real_44_3_pipe;
                output_imag_44_3_pipe <= output_imag_44_3_pipe;
		output_real_45_3_pipe <= output_real_45_3_pipe;
                output_imag_45_3_pipe <= output_imag_45_3_pipe;
		output_real_46_3_pipe <= output_real_46_3_pipe;
                output_imag_46_3_pipe <= output_imag_46_3_pipe;
		output_real_47_3_pipe <= output_real_47_3_pipe;
                output_imag_47_3_pipe <= output_imag_47_3_pipe;
		output_real_48_3_pipe <= output_real_48_3_pipe;
                output_imag_48_3_pipe <= output_imag_48_3_pipe;
		output_real_49_3_pipe <= output_real_49_3_pipe;
                output_imag_49_3_pipe <= output_imag_49_3_pipe;
		output_real_50_3_pipe <= output_real_50_3_pipe;
                output_imag_50_3_pipe <= output_imag_50_3_pipe;
		output_real_51_3_pipe <= output_real_51_3_pipe;
                output_imag_51_3_pipe <= output_imag_51_3_pipe;
		output_real_52_3_pipe <= output_real_52_3_pipe;
                output_imag_52_3_pipe <= output_imag_52_3_pipe;
		output_real_53_3_pipe <= output_real_53_3_pipe;
                output_imag_53_3_pipe <= output_imag_53_3_pipe;
		output_real_54_3_pipe <= output_real_54_3_pipe;
                output_imag_54_3_pipe <= output_imag_54_3_pipe;
		output_real_55_3_pipe <= output_real_55_3_pipe;
                output_imag_55_3_pipe <= output_imag_55_3_pipe;
		output_real_56_3_pipe <= output_real_56_3_pipe;
                output_imag_56_3_pipe <= output_imag_56_3_pipe;
		output_real_57_3_pipe <= output_real_57_3_pipe;
                output_imag_57_3_pipe <= output_imag_57_3_pipe;
		output_real_58_3_pipe <= output_real_58_3_pipe;
                output_imag_58_3_pipe <= output_imag_58_3_pipe;
		output_real_59_3_pipe <= output_real_59_3_pipe;
                output_imag_59_3_pipe <= output_imag_59_3_pipe;
		output_real_60_3_pipe <= output_real_60_3_pipe;
                output_imag_60_3_pipe <= output_imag_60_3_pipe;
		output_real_61_3_pipe <= output_real_61_3_pipe;
                output_imag_61_3_pipe <= output_imag_61_3_pipe;
		output_real_62_3_pipe <= output_real_62_3_pipe;
                output_imag_62_3_pipe <= output_imag_62_3_pipe;
		output_real_63_3_pipe <= output_real_63_3_pipe;
                output_imag_63_3_pipe <= output_imag_63_3_pipe;
                end
        end
end




assign output_real_0_0 = output_real_0_0_pipe;
assign output_imag_0_0 = output_imag_0_0_pipe;
assign output_real_1_0 = output_real_1_0_pipe;
assign output_imag_1_0 = output_imag_1_0_pipe;
assign output_real_2_0 = output_real_2_0_pipe;
assign output_imag_2_0 = output_imag_2_0_pipe;
assign output_real_3_0 = output_real_3_0_pipe;
assign output_imag_3_0 = output_imag_3_0_pipe;
assign output_real_4_0 = output_real_4_0_pipe;
assign output_imag_4_0 = output_imag_4_0_pipe;
assign output_real_5_0 = output_real_5_0_pipe;
assign output_imag_5_0 = output_imag_5_0_pipe;
assign output_real_6_0 = output_real_6_0_pipe;
assign output_imag_6_0 = output_imag_6_0_pipe;
assign output_real_7_0 = output_real_7_0_pipe;
assign output_imag_7_0 = output_imag_7_0_pipe;
assign output_real_8_0 = output_real_8_0_pipe;
assign output_imag_8_0 = output_imag_8_0_pipe;
assign output_real_9_0 = output_real_9_0_pipe;
assign output_imag_9_0 = output_imag_9_0_pipe;
assign output_real_10_0 = output_real_10_0_pipe;
assign output_imag_10_0 = output_imag_10_0_pipe;
assign output_real_11_0 = output_real_11_0_pipe;
assign output_imag_11_0 = output_imag_11_0_pipe;
assign output_real_12_0 = output_real_12_0_pipe;
assign output_imag_12_0 = output_imag_12_0_pipe;
assign output_real_13_0 = output_real_13_0_pipe;
assign output_imag_13_0 = output_imag_13_0_pipe;
assign output_real_14_0 = output_real_14_0_pipe;
assign output_imag_14_0 = output_imag_14_0_pipe;
assign output_real_15_0 = output_real_15_0_pipe;
assign output_imag_15_0 = output_imag_15_0_pipe;
assign output_real_16_0 = output_real_16_0_pipe;
assign output_imag_16_0 = output_imag_16_0_pipe;
assign output_real_17_0 = output_real_17_0_pipe;
assign output_imag_17_0 = output_imag_17_0_pipe;
assign output_real_18_0 = output_real_18_0_pipe;
assign output_imag_18_0 = output_imag_18_0_pipe;
assign output_real_19_0 = output_real_19_0_pipe;
assign output_imag_19_0 = output_imag_19_0_pipe;
assign output_real_20_0 = output_real_20_0_pipe;
assign output_imag_20_0 = output_imag_20_0_pipe;
assign output_real_21_0 = output_real_21_0_pipe;
assign output_imag_21_0 = output_imag_21_0_pipe;
assign output_real_22_0 = output_real_22_0_pipe;
assign output_imag_22_0 = output_imag_22_0_pipe;
assign output_real_23_0 = output_real_23_0_pipe;
assign output_imag_23_0 = output_imag_23_0_pipe;
assign output_real_24_0 = output_real_24_0_pipe;
assign output_imag_24_0 = output_imag_24_0_pipe;
assign output_real_25_0 = output_real_25_0_pipe;
assign output_imag_25_0 = output_imag_25_0_pipe;
assign output_real_26_0 = output_real_26_0_pipe;
assign output_imag_26_0 = output_imag_26_0_pipe;
assign output_real_27_0 = output_real_27_0_pipe;
assign output_imag_27_0 = output_imag_27_0_pipe;
assign output_real_28_0 = output_real_28_0_pipe;
assign output_imag_28_0 = output_imag_28_0_pipe;
assign output_real_29_0 = output_real_29_0_pipe;
assign output_imag_29_0 = output_imag_29_0_pipe;
assign output_real_30_0 = output_real_30_0_pipe;
assign output_imag_30_0 = output_imag_30_0_pipe;
assign output_real_31_0 = output_real_31_0_pipe;
assign output_imag_31_0 = output_imag_31_0_pipe;
assign output_real_32_0 = output_real_32_0_pipe;
assign output_imag_32_0 = output_imag_32_0_pipe;
assign output_real_33_0 = output_real_33_0_pipe;
assign output_imag_33_0 = output_imag_33_0_pipe;
assign output_real_34_0 = output_real_34_0_pipe;
assign output_imag_34_0 = output_imag_34_0_pipe;
assign output_real_35_0 = output_real_35_0_pipe;
assign output_imag_35_0 = output_imag_35_0_pipe;
assign output_real_36_0 = output_real_36_0_pipe;
assign output_imag_36_0 = output_imag_36_0_pipe;
assign output_real_37_0 = output_real_37_0_pipe;
assign output_imag_37_0 = output_imag_37_0_pipe;
assign output_real_38_0 = output_real_38_0_pipe;
assign output_imag_38_0 = output_imag_38_0_pipe;
assign output_real_39_0 = output_real_39_0_pipe;
assign output_imag_39_0 = output_imag_39_0_pipe;
assign output_real_40_0 = output_real_40_0_pipe;
assign output_imag_40_0 = output_imag_40_0_pipe;
assign output_real_41_0 = output_real_41_0_pipe;
assign output_imag_41_0 = output_imag_41_0_pipe;
assign output_real_42_0 = output_real_42_0_pipe;
assign output_imag_42_0 = output_imag_42_0_pipe;
assign output_real_43_0 = output_real_43_0_pipe;
assign output_imag_43_0 = output_imag_43_0_pipe;
assign output_real_44_0 = output_real_44_0_pipe;
assign output_imag_44_0 = output_imag_44_0_pipe;
assign output_real_45_0 = output_real_45_0_pipe;
assign output_imag_45_0 = output_imag_45_0_pipe;
assign output_real_46_0 = output_real_46_0_pipe;
assign output_imag_46_0 = output_imag_46_0_pipe;
assign output_real_47_0 = output_real_47_0_pipe;
assign output_imag_47_0 = output_imag_47_0_pipe;
assign output_real_48_0 = output_real_48_0_pipe;
assign output_imag_48_0 = output_imag_48_0_pipe;
assign output_real_49_0 = output_real_49_0_pipe;
assign output_imag_49_0 = output_imag_49_0_pipe;
assign output_real_50_0 = output_real_50_0_pipe;
assign output_imag_50_0 = output_imag_50_0_pipe;
assign output_real_51_0 = output_real_51_0_pipe;
assign output_imag_51_0 = output_imag_51_0_pipe;
assign output_real_52_0 = output_real_52_0_pipe;
assign output_imag_52_0 = output_imag_52_0_pipe;
assign output_real_53_0 = output_real_53_0_pipe;
assign output_imag_53_0 = output_imag_53_0_pipe;
assign output_real_54_0 = output_real_54_0_pipe;
assign output_imag_54_0 = output_imag_54_0_pipe;
assign output_real_55_0 = output_real_55_0_pipe;
assign output_imag_55_0 = output_imag_55_0_pipe;
assign output_real_56_0 = output_real_56_0_pipe;
assign output_imag_56_0 = output_imag_56_0_pipe;
assign output_real_57_0 = output_real_57_0_pipe;
assign output_imag_57_0 = output_imag_57_0_pipe;
assign output_real_58_0 = output_real_58_0_pipe;
assign output_imag_58_0 = output_imag_58_0_pipe;
assign output_real_59_0 = output_real_59_0_pipe;
assign output_imag_59_0 = output_imag_59_0_pipe;
assign output_real_60_0 = output_real_60_0_pipe;
assign output_imag_60_0 = output_imag_60_0_pipe;
assign output_real_61_0 = output_real_61_0_pipe;
assign output_imag_61_0 = output_imag_61_0_pipe;
assign output_real_62_0 = output_real_62_0_pipe;
assign output_imag_62_0 = output_imag_62_0_pipe;
assign output_real_63_0 = output_real_63_0_pipe;
assign output_imag_63_0 = output_imag_63_0_pipe;
assign output_real_0_1 = output_real_0_1_pipe;
assign output_imag_0_1 = output_imag_0_1_pipe;
assign output_real_1_1 = output_real_1_1_pipe;
assign output_imag_1_1 = output_imag_1_1_pipe;
assign output_real_2_1 = output_real_2_1_pipe;
assign output_imag_2_1 = output_imag_2_1_pipe;
assign output_real_3_1 = output_real_3_1_pipe;
assign output_imag_3_1 = output_imag_3_1_pipe;
assign output_real_4_1 = output_real_4_1_pipe;
assign output_imag_4_1 = output_imag_4_1_pipe;
assign output_real_5_1 = output_real_5_1_pipe;
assign output_imag_5_1 = output_imag_5_1_pipe;
assign output_real_6_1 = output_real_6_1_pipe;
assign output_imag_6_1 = output_imag_6_1_pipe;
assign output_real_7_1 = output_real_7_1_pipe;
assign output_imag_7_1 = output_imag_7_1_pipe;
assign output_real_8_1 = output_real_8_1_pipe;
assign output_imag_8_1 = output_imag_8_1_pipe;
assign output_real_9_1 = output_real_9_1_pipe;
assign output_imag_9_1 = output_imag_9_1_pipe;
assign output_real_10_1 = output_real_10_1_pipe;
assign output_imag_10_1 = output_imag_10_1_pipe;
assign output_real_11_1 = output_real_11_1_pipe;
assign output_imag_11_1 = output_imag_11_1_pipe;
assign output_real_12_1 = output_real_12_1_pipe;
assign output_imag_12_1 = output_imag_12_1_pipe;
assign output_real_13_1 = output_real_13_1_pipe;
assign output_imag_13_1 = output_imag_13_1_pipe;
assign output_real_14_1 = output_real_14_1_pipe;
assign output_imag_14_1 = output_imag_14_1_pipe;
assign output_real_15_1 = output_real_15_1_pipe;
assign output_imag_15_1 = output_imag_15_1_pipe;
assign output_real_16_1 = output_real_16_1_pipe;
assign output_imag_16_1 = output_imag_16_1_pipe;
assign output_real_17_1 = output_real_17_1_pipe;
assign output_imag_17_1 = output_imag_17_1_pipe;
assign output_real_18_1 = output_real_18_1_pipe;
assign output_imag_18_1 = output_imag_18_1_pipe;
assign output_real_19_1 = output_real_19_1_pipe;
assign output_imag_19_1 = output_imag_19_1_pipe;
assign output_real_20_1 = output_real_20_1_pipe;
assign output_imag_20_1 = output_imag_20_1_pipe;
assign output_real_21_1 = output_real_21_1_pipe;
assign output_imag_21_1 = output_imag_21_1_pipe;
assign output_real_22_1 = output_real_22_1_pipe;
assign output_imag_22_1 = output_imag_22_1_pipe;
assign output_real_23_1 = output_real_23_1_pipe;
assign output_imag_23_1 = output_imag_23_1_pipe;
assign output_real_24_1 = output_real_24_1_pipe;
assign output_imag_24_1 = output_imag_24_1_pipe;
assign output_real_25_1 = output_real_25_1_pipe;
assign output_imag_25_1 = output_imag_25_1_pipe;
assign output_real_26_1 = output_real_26_1_pipe;
assign output_imag_26_1 = output_imag_26_1_pipe;
assign output_real_27_1 = output_real_27_1_pipe;
assign output_imag_27_1 = output_imag_27_1_pipe;
assign output_real_28_1 = output_real_28_1_pipe;
assign output_imag_28_1 = output_imag_28_1_pipe;
assign output_real_29_1 = output_real_29_1_pipe;
assign output_imag_29_1 = output_imag_29_1_pipe;
assign output_real_30_1 = output_real_30_1_pipe;
assign output_imag_30_1 = output_imag_30_1_pipe;
assign output_real_31_1 = output_real_31_1_pipe;
assign output_imag_31_1 = output_imag_31_1_pipe;
assign output_real_32_1 = output_real_32_1_pipe;
assign output_imag_32_1 = output_imag_32_1_pipe;
assign output_real_33_1 = output_real_33_1_pipe;
assign output_imag_33_1 = output_imag_33_1_pipe;
assign output_real_34_1 = output_real_34_1_pipe;
assign output_imag_34_1 = output_imag_34_1_pipe;
assign output_real_35_1 = output_real_35_1_pipe;
assign output_imag_35_1 = output_imag_35_1_pipe;
assign output_real_36_1 = output_real_36_1_pipe;
assign output_imag_36_1 = output_imag_36_1_pipe;
assign output_real_37_1 = output_real_37_1_pipe;
assign output_imag_37_1 = output_imag_37_1_pipe;
assign output_real_38_1 = output_real_38_1_pipe;
assign output_imag_38_1 = output_imag_38_1_pipe;
assign output_real_39_1 = output_real_39_1_pipe;
assign output_imag_39_1 = output_imag_39_1_pipe;
assign output_real_40_1 = output_real_40_1_pipe;
assign output_imag_40_1 = output_imag_40_1_pipe;
assign output_real_41_1 = output_real_41_1_pipe;
assign output_imag_41_1 = output_imag_41_1_pipe;
assign output_real_42_1 = output_real_42_1_pipe;
assign output_imag_42_1 = output_imag_42_1_pipe;
assign output_real_43_1 = output_real_43_1_pipe;
assign output_imag_43_1 = output_imag_43_1_pipe;
assign output_real_44_1 = output_real_44_1_pipe;
assign output_imag_44_1 = output_imag_44_1_pipe;
assign output_real_45_1 = output_real_45_1_pipe;
assign output_imag_45_1 = output_imag_45_1_pipe;
assign output_real_46_1 = output_real_46_1_pipe;
assign output_imag_46_1 = output_imag_46_1_pipe;
assign output_real_47_1 = output_real_47_1_pipe;
assign output_imag_47_1 = output_imag_47_1_pipe;
assign output_real_48_1 = output_real_48_1_pipe;
assign output_imag_48_1 = output_imag_48_1_pipe;
assign output_real_49_1 = output_real_49_1_pipe;
assign output_imag_49_1 = output_imag_49_1_pipe;
assign output_real_50_1 = output_real_50_1_pipe;
assign output_imag_50_1 = output_imag_50_1_pipe;
assign output_real_51_1 = output_real_51_1_pipe;
assign output_imag_51_1 = output_imag_51_1_pipe;
assign output_real_52_1 = output_real_52_1_pipe;
assign output_imag_52_1 = output_imag_52_1_pipe;
assign output_real_53_1 = output_real_53_1_pipe;
assign output_imag_53_1 = output_imag_53_1_pipe;
assign output_real_54_1 = output_real_54_1_pipe;
assign output_imag_54_1 = output_imag_54_1_pipe;
assign output_real_55_1 = output_real_55_1_pipe;
assign output_imag_55_1 = output_imag_55_1_pipe;
assign output_real_56_1 = output_real_56_1_pipe;
assign output_imag_56_1 = output_imag_56_1_pipe;
assign output_real_57_1 = output_real_57_1_pipe;
assign output_imag_57_1 = output_imag_57_1_pipe;
assign output_real_58_1 = output_real_58_1_pipe;
assign output_imag_58_1 = output_imag_58_1_pipe;
assign output_real_59_1 = output_real_59_1_pipe;
assign output_imag_59_1 = output_imag_59_1_pipe;
assign output_real_60_1 = output_real_60_1_pipe;
assign output_imag_60_1 = output_imag_60_1_pipe;
assign output_real_61_1 = output_real_61_1_pipe;
assign output_imag_61_1 = output_imag_61_1_pipe;
assign output_real_62_1 = output_real_62_1_pipe;
assign output_imag_62_1 = output_imag_62_1_pipe;
assign output_real_63_1 = output_real_63_1_pipe;
assign output_imag_63_1 = output_imag_63_1_pipe;
assign output_real_0_2 = output_real_0_2_pipe;
assign output_imag_0_2 = output_imag_0_2_pipe;
assign output_real_1_2 = output_real_1_2_pipe;
assign output_imag_1_2 = output_imag_1_2_pipe;
assign output_real_2_2 = output_real_2_2_pipe;
assign output_imag_2_2 = output_imag_2_2_pipe;
assign output_real_3_2 = output_real_3_2_pipe;
assign output_imag_3_2 = output_imag_3_2_pipe;
assign output_real_4_2 = output_real_4_2_pipe;
assign output_imag_4_2 = output_imag_4_2_pipe;
assign output_real_5_2 = output_real_5_2_pipe;
assign output_imag_5_2 = output_imag_5_2_pipe;
assign output_real_6_2 = output_real_6_2_pipe;
assign output_imag_6_2 = output_imag_6_2_pipe;
assign output_real_7_2 = output_real_7_2_pipe;
assign output_imag_7_2 = output_imag_7_2_pipe;
assign output_real_8_2 = output_real_8_2_pipe;
assign output_imag_8_2 = output_imag_8_2_pipe;
assign output_real_9_2 = output_real_9_2_pipe;
assign output_imag_9_2 = output_imag_9_2_pipe;
assign output_real_10_2 = output_real_10_2_pipe;
assign output_imag_10_2 = output_imag_10_2_pipe;
assign output_real_11_2 = output_real_11_2_pipe;
assign output_imag_11_2 = output_imag_11_2_pipe;
assign output_real_12_2 = output_real_12_2_pipe;
assign output_imag_12_2 = output_imag_12_2_pipe;
assign output_real_13_2 = output_real_13_2_pipe;
assign output_imag_13_2 = output_imag_13_2_pipe;
assign output_real_14_2 = output_real_14_2_pipe;
assign output_imag_14_2 = output_imag_14_2_pipe;
assign output_real_15_2 = output_real_15_2_pipe;
assign output_imag_15_2 = output_imag_15_2_pipe;
assign output_real_16_2 = output_real_16_2_pipe;
assign output_imag_16_2 = output_imag_16_2_pipe;
assign output_real_17_2 = output_real_17_2_pipe;
assign output_imag_17_2 = output_imag_17_2_pipe;
assign output_real_18_2 = output_real_18_2_pipe;
assign output_imag_18_2 = output_imag_18_2_pipe;
assign output_real_19_2 = output_real_19_2_pipe;
assign output_imag_19_2 = output_imag_19_2_pipe;
assign output_real_20_2 = output_real_20_2_pipe;
assign output_imag_20_2 = output_imag_20_2_pipe;
assign output_real_21_2 = output_real_21_2_pipe;
assign output_imag_21_2 = output_imag_21_2_pipe;
assign output_real_22_2 = output_real_22_2_pipe;
assign output_imag_22_2 = output_imag_22_2_pipe;
assign output_real_23_2 = output_real_23_2_pipe;
assign output_imag_23_2 = output_imag_23_2_pipe;
assign output_real_24_2 = output_real_24_2_pipe;
assign output_imag_24_2 = output_imag_24_2_pipe;
assign output_real_25_2 = output_real_25_2_pipe;
assign output_imag_25_2 = output_imag_25_2_pipe;
assign output_real_26_2 = output_real_26_2_pipe;
assign output_imag_26_2 = output_imag_26_2_pipe;
assign output_real_27_2 = output_real_27_2_pipe;
assign output_imag_27_2 = output_imag_27_2_pipe;
assign output_real_28_2 = output_real_28_2_pipe;
assign output_imag_28_2 = output_imag_28_2_pipe;
assign output_real_29_2 = output_real_29_2_pipe;
assign output_imag_29_2 = output_imag_29_2_pipe;
assign output_real_30_2 = output_real_30_2_pipe;
assign output_imag_30_2 = output_imag_30_2_pipe;
assign output_real_31_2 = output_real_31_2_pipe;
assign output_imag_31_2 = output_imag_31_2_pipe;
assign output_real_32_2 = output_real_32_2_pipe;
assign output_imag_32_2 = output_imag_32_2_pipe;
assign output_real_33_2 = output_real_33_2_pipe;
assign output_imag_33_2 = output_imag_33_2_pipe;
assign output_real_34_2 = output_real_34_2_pipe;
assign output_imag_34_2 = output_imag_34_2_pipe;
assign output_real_35_2 = output_real_35_2_pipe;
assign output_imag_35_2 = output_imag_35_2_pipe;
assign output_real_36_2 = output_real_36_2_pipe;
assign output_imag_36_2 = output_imag_36_2_pipe;
assign output_real_37_2 = output_real_37_2_pipe;
assign output_imag_37_2 = output_imag_37_2_pipe;
assign output_real_38_2 = output_real_38_2_pipe;
assign output_imag_38_2 = output_imag_38_2_pipe;
assign output_real_39_2 = output_real_39_2_pipe;
assign output_imag_39_2 = output_imag_39_2_pipe;
assign output_real_40_2 = output_real_40_2_pipe;
assign output_imag_40_2 = output_imag_40_2_pipe;
assign output_real_41_2 = output_real_41_2_pipe;
assign output_imag_41_2 = output_imag_41_2_pipe;
assign output_real_42_2 = output_real_42_2_pipe;
assign output_imag_42_2 = output_imag_42_2_pipe;
assign output_real_43_2 = output_real_43_2_pipe;
assign output_imag_43_2 = output_imag_43_2_pipe;
assign output_real_44_2 = output_real_44_2_pipe;
assign output_imag_44_2 = output_imag_44_2_pipe;
assign output_real_45_2 = output_real_45_2_pipe;
assign output_imag_45_2 = output_imag_45_2_pipe;
assign output_real_46_2 = output_real_46_2_pipe;
assign output_imag_46_2 = output_imag_46_2_pipe;
assign output_real_47_2 = output_real_47_2_pipe;
assign output_imag_47_2 = output_imag_47_2_pipe;
assign output_real_48_2 = output_real_48_2_pipe;
assign output_imag_48_2 = output_imag_48_2_pipe;
assign output_real_49_2 = output_real_49_2_pipe;
assign output_imag_49_2 = output_imag_49_2_pipe;
assign output_real_50_2 = output_real_50_2_pipe;
assign output_imag_50_2 = output_imag_50_2_pipe;
assign output_real_51_2 = output_real_51_2_pipe;
assign output_imag_51_2 = output_imag_51_2_pipe;
assign output_real_52_2 = output_real_52_2_pipe;
assign output_imag_52_2 = output_imag_52_2_pipe;
assign output_real_53_2 = output_real_53_2_pipe;
assign output_imag_53_2 = output_imag_53_2_pipe;
assign output_real_54_2 = output_real_54_2_pipe;
assign output_imag_54_2 = output_imag_54_2_pipe;
assign output_real_55_2 = output_real_55_2_pipe;
assign output_imag_55_2 = output_imag_55_2_pipe;
assign output_real_56_2 = output_real_56_2_pipe;
assign output_imag_56_2 = output_imag_56_2_pipe;
assign output_real_57_2 = output_real_57_2_pipe;
assign output_imag_57_2 = output_imag_57_2_pipe;
assign output_real_58_2 = output_real_58_2_pipe;
assign output_imag_58_2 = output_imag_58_2_pipe;
assign output_real_59_2 = output_real_59_2_pipe;
assign output_imag_59_2 = output_imag_59_2_pipe;
assign output_real_60_2 = output_real_60_2_pipe;
assign output_imag_60_2 = output_imag_60_2_pipe;
assign output_real_61_2 = output_real_61_2_pipe;
assign output_imag_61_2 = output_imag_61_2_pipe;
assign output_real_62_2 = output_real_62_2_pipe;
assign output_imag_62_2 = output_imag_62_2_pipe;
assign output_real_63_2 = output_real_63_2_pipe;
assign output_imag_63_2 = output_imag_63_2_pipe;
assign output_real_0_3 = output_real_0_3_pipe;
assign output_imag_0_3 = output_imag_0_3_pipe;
assign output_real_1_3 = output_real_1_3_pipe;
assign output_imag_1_3 = output_imag_1_3_pipe;
assign output_real_2_3 = output_real_2_3_pipe;
assign output_imag_2_3 = output_imag_2_3_pipe;
assign output_real_3_3 = output_real_3_3_pipe;
assign output_imag_3_3 = output_imag_3_3_pipe;
assign output_real_4_3 = output_real_4_3_pipe;
assign output_imag_4_3 = output_imag_4_3_pipe;
assign output_real_5_3 = output_real_5_3_pipe;
assign output_imag_5_3 = output_imag_5_3_pipe;
assign output_real_6_3 = output_real_6_3_pipe;
assign output_imag_6_3 = output_imag_6_3_pipe;
assign output_real_7_3 = output_real_7_3_pipe;
assign output_imag_7_3 = output_imag_7_3_pipe;
assign output_real_8_3 = output_real_8_3_pipe;
assign output_imag_8_3 = output_imag_8_3_pipe;
assign output_real_9_3 = output_real_9_3_pipe;
assign output_imag_9_3 = output_imag_9_3_pipe;
assign output_real_10_3 = output_real_10_3_pipe;
assign output_imag_10_3 = output_imag_10_3_pipe;
assign output_real_11_3 = output_real_11_3_pipe;
assign output_imag_11_3 = output_imag_11_3_pipe;
assign output_real_12_3 = output_real_12_3_pipe;
assign output_imag_12_3 = output_imag_12_3_pipe;
assign output_real_13_3 = output_real_13_3_pipe;
assign output_imag_13_3 = output_imag_13_3_pipe;
assign output_real_14_3 = output_real_14_3_pipe;
assign output_imag_14_3 = output_imag_14_3_pipe;
assign output_real_15_3 = output_real_15_3_pipe;
assign output_imag_15_3 = output_imag_15_3_pipe;
assign output_real_16_3 = output_real_16_3_pipe;
assign output_imag_16_3 = output_imag_16_3_pipe;
assign output_real_17_3 = output_real_17_3_pipe;
assign output_imag_17_3 = output_imag_17_3_pipe;
assign output_real_18_3 = output_real_18_3_pipe;
assign output_imag_18_3 = output_imag_18_3_pipe;
assign output_real_19_3 = output_real_19_3_pipe;
assign output_imag_19_3 = output_imag_19_3_pipe;
assign output_real_20_3 = output_real_20_3_pipe;
assign output_imag_20_3 = output_imag_20_3_pipe;
assign output_real_21_3 = output_real_21_3_pipe;
assign output_imag_21_3 = output_imag_21_3_pipe;
assign output_real_22_3 = output_real_22_3_pipe;
assign output_imag_22_3 = output_imag_22_3_pipe;
assign output_real_23_3 = output_real_23_3_pipe;
assign output_imag_23_3 = output_imag_23_3_pipe;
assign output_real_24_3 = output_real_24_3_pipe;
assign output_imag_24_3 = output_imag_24_3_pipe;
assign output_real_25_3 = output_real_25_3_pipe;
assign output_imag_25_3 = output_imag_25_3_pipe;
assign output_real_26_3 = output_real_26_3_pipe;
assign output_imag_26_3 = output_imag_26_3_pipe;
assign output_real_27_3 = output_real_27_3_pipe;
assign output_imag_27_3 = output_imag_27_3_pipe;
assign output_real_28_3 = output_real_28_3_pipe;
assign output_imag_28_3 = output_imag_28_3_pipe;
assign output_real_29_3 = output_real_29_3_pipe;
assign output_imag_29_3 = output_imag_29_3_pipe;
assign output_real_30_3 = output_real_30_3_pipe;
assign output_imag_30_3 = output_imag_30_3_pipe;
assign output_real_31_3 = output_real_31_3_pipe;
assign output_imag_31_3 = output_imag_31_3_pipe;
assign output_real_32_3 = output_real_32_3_pipe;
assign output_imag_32_3 = output_imag_32_3_pipe;
assign output_real_33_3 = output_real_33_3_pipe;
assign output_imag_33_3 = output_imag_33_3_pipe;
assign output_real_34_3 = output_real_34_3_pipe;
assign output_imag_34_3 = output_imag_34_3_pipe;
assign output_real_35_3 = output_real_35_3_pipe;
assign output_imag_35_3 = output_imag_35_3_pipe;
assign output_real_36_3 = output_real_36_3_pipe;
assign output_imag_36_3 = output_imag_36_3_pipe;
assign output_real_37_3 = output_real_37_3_pipe;
assign output_imag_37_3 = output_imag_37_3_pipe;
assign output_real_38_3 = output_real_38_3_pipe;
assign output_imag_38_3 = output_imag_38_3_pipe;
assign output_real_39_3 = output_real_39_3_pipe;
assign output_imag_39_3 = output_imag_39_3_pipe;
assign output_real_40_3 = output_real_40_3_pipe;
assign output_imag_40_3 = output_imag_40_3_pipe;
assign output_real_41_3 = output_real_41_3_pipe;
assign output_imag_41_3 = output_imag_41_3_pipe;
assign output_real_42_3 = output_real_42_3_pipe;
assign output_imag_42_3 = output_imag_42_3_pipe;
assign output_real_43_3 = output_real_43_3_pipe;
assign output_imag_43_3 = output_imag_43_3_pipe;
assign output_real_44_3 = output_real_44_3_pipe;
assign output_imag_44_3 = output_imag_44_3_pipe;
assign output_real_45_3 = output_real_45_3_pipe;
assign output_imag_45_3 = output_imag_45_3_pipe;
assign output_real_46_3 = output_real_46_3_pipe;
assign output_imag_46_3 = output_imag_46_3_pipe;
assign output_real_47_3 = output_real_47_3_pipe;
assign output_imag_47_3 = output_imag_47_3_pipe;
assign output_real_48_3 = output_real_48_3_pipe;
assign output_imag_48_3 = output_imag_48_3_pipe;
assign output_real_49_3 = output_real_49_3_pipe;
assign output_imag_49_3 = output_imag_49_3_pipe;
assign output_real_50_3 = output_real_50_3_pipe;
assign output_imag_50_3 = output_imag_50_3_pipe;
assign output_real_51_3 = output_real_51_3_pipe;
assign output_imag_51_3 = output_imag_51_3_pipe;
assign output_real_52_3 = output_real_52_3_pipe;
assign output_imag_52_3 = output_imag_52_3_pipe;
assign output_real_53_3 = output_real_53_3_pipe;
assign output_imag_53_3 = output_imag_53_3_pipe;
assign output_real_54_3 = output_real_54_3_pipe;
assign output_imag_54_3 = output_imag_54_3_pipe;
assign output_real_55_3 = output_real_55_3_pipe;
assign output_imag_55_3 = output_imag_55_3_pipe;
assign output_real_56_3 = output_real_56_3_pipe;
assign output_imag_56_3 = output_imag_56_3_pipe;
assign output_real_57_3 = output_real_57_3_pipe;
assign output_imag_57_3 = output_imag_57_3_pipe;
assign output_real_58_3 = output_real_58_3_pipe;
assign output_imag_58_3 = output_imag_58_3_pipe;
assign output_real_59_3 = output_real_59_3_pipe;
assign output_imag_59_3 = output_imag_59_3_pipe;
assign output_real_60_3 = output_real_60_3_pipe;
assign output_imag_60_3 = output_imag_60_3_pipe;
assign output_real_61_3 = output_real_61_3_pipe;
assign output_imag_61_3 = output_imag_61_3_pipe;
assign output_real_62_3 = output_real_62_3_pipe;
assign output_imag_62_3 = output_imag_62_3_pipe;
assign output_real_63_3 = output_real_63_3_pipe;
assign output_imag_63_3 = output_imag_63_3_pipe;


endmodule
