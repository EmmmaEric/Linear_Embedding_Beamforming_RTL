
module memory_rom_33(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbccabc25;
    11'b00000000001: data <= 32'hb9a3b852;
    11'b00000000010: data <= 32'h397b392a;
    11'b00000000011: data <= 32'h39953ef5;
    11'b00000000100: data <= 32'hbc183d91;
    11'b00000000101: data <= 32'hc0b620ba;
    11'b00000000110: data <= 32'hbf18b7b7;
    11'b00000000111: data <= 32'hb3e337e5;
    11'b00000001000: data <= 32'h390d3cca;
    11'b00000001001: data <= 32'h3b103522;
    11'b00000001010: data <= 32'h3d49ba6a;
    11'b00000001011: data <= 32'h3e91b166;
    11'b00000001100: data <= 32'h3bc13ea0;
    11'b00000001101: data <= 32'hb284404c;
    11'b00000001110: data <= 32'hb66b36f0;
    11'b00000001111: data <= 32'h3761be42;
    11'b00000010000: data <= 32'h3a35bfe0;
    11'b00000010001: data <= 32'hb0aabd25;
    11'b00000010010: data <= 32'hba24bba2;
    11'b00000010011: data <= 32'h33f1bbb1;
    11'b00000010100: data <= 32'h3e67b640;
    11'b00000010101: data <= 32'h3c03382d;
    11'b00000010110: data <= 32'hbd6838fb;
    11'b00000010111: data <= 32'hc1b3ad0b;
    11'b00000011000: data <= 32'hc01bb470;
    11'b00000011001: data <= 32'hb6fb3624;
    11'b00000011010: data <= 32'h2e8238b5;
    11'b00000011011: data <= 32'hb14cb578;
    11'b00000011100: data <= 32'h2fdcbb37;
    11'b00000011101: data <= 32'h3b4e370a;
    11'b00000011110: data <= 32'h3bfe4110;
    11'b00000011111: data <= 32'h3431418d;
    11'b00000100000: data <= 32'haf7c3a35;
    11'b00000100001: data <= 32'h343ebc67;
    11'b00000100010: data <= 32'h36a7bc67;
    11'b00000100011: data <= 32'hac8fb470;
    11'b00000100100: data <= 32'h9f09b690;
    11'b00000100101: data <= 32'h3d55bce6;
    11'b00000100110: data <= 32'h40d9bcbb;
    11'b00000100111: data <= 32'h3d76b107;
    11'b00000101000: data <= 32'hbc733727;
    11'b00000101001: data <= 32'hc0b128c2;
    11'b00000101010: data <= 32'hbd89b6f3;
    11'b00000101011: data <= 32'hb0d8b5e4;
    11'b00000101100: data <= 32'hb68ab7ec;
    11'b00000101101: data <= 32'hbd0abcae;
    11'b00000101110: data <= 32'hbb17bca0;
    11'b00000101111: data <= 32'h37af3828;
    11'b00000110000: data <= 32'h3c1140fc;
    11'b00000110001: data <= 32'h31964111;
    11'b00000110010: data <= 32'hb9943a19;
    11'b00000110011: data <= 32'hb911b6d7;
    11'b00000110100: data <= 32'hb3dd312f;
    11'b00000110101: data <= 32'haf703b65;
    11'b00000110110: data <= 32'h3698305b;
    11'b00000110111: data <= 32'h3efcbd3d;
    11'b00000111000: data <= 32'h4130bd5a;
    11'b00000111001: data <= 32'h3e4b2eaa;
    11'b00000111010: data <= 32'hb6953c2f;
    11'b00000111011: data <= 32'hbc773728;
    11'b00000111100: data <= 32'hb1f5b912;
    11'b00000111101: data <= 32'h35c2bc54;
    11'b00000111110: data <= 32'hb979bd00;
    11'b00000111111: data <= 32'hbf1fbe86;
    11'b00001000000: data <= 32'hbc31bde0;
    11'b00001000001: data <= 32'h39e3ac0a;
    11'b00001000010: data <= 32'h3cca3dfc;
    11'b00001000011: data <= 32'hb26f3e2e;
    11'b00001000100: data <= 32'hbe6336c1;
    11'b00001000101: data <= 32'hbe4d2dcf;
    11'b00001000110: data <= 32'hba893c46;
    11'b00001000111: data <= 32'hb5eb3e19;
    11'b00001001000: data <= 32'h2d6e327d;
    11'b00001001001: data <= 32'h3c7dbd6f;
    11'b00001001010: data <= 32'h3fd5bb90;
    11'b00001001011: data <= 32'h3dfa3c0e;
    11'b00001001100: data <= 32'h356a4003;
    11'b00001001101: data <= 32'h2d8f3bb4;
    11'b00001001110: data <= 32'h3a08b8ba;
    11'b00001001111: data <= 32'h3945bc7b;
    11'b00001010000: data <= 32'hb9cfbc3d;
    11'b00001010001: data <= 32'hbe3cbd82;
    11'b00001010010: data <= 32'hb558be9a;
    11'b00001010011: data <= 32'h3e36bbca;
    11'b00001010100: data <= 32'h3e3630ce;
    11'b00001010101: data <= 32'hb70b3737;
    11'b00001010110: data <= 32'hc01629f5;
    11'b00001010111: data <= 32'hbf3f340f;
    11'b00001011000: data <= 32'hbb0b3ca8;
    11'b00001011001: data <= 32'hb9a63cb6;
    11'b00001011010: data <= 32'hbad1b56b;
    11'b00001011011: data <= 32'hb230be11;
    11'b00001011100: data <= 32'h3b4ab763;
    11'b00001011101: data <= 32'h3ce13f3c;
    11'b00001011110: data <= 32'h39e4412f;
    11'b00001011111: data <= 32'h38943ce5;
    11'b00001100000: data <= 32'h3ac2b449;
    11'b00001100001: data <= 32'h3731b577;
    11'b00001100010: data <= 32'hb9a72ad7;
    11'b00001100011: data <= 32'hbb9cb844;
    11'b00001100100: data <= 32'h3921be6c;
    11'b00001100101: data <= 32'h40aebeb6;
    11'b00001100110: data <= 32'h3f83b9ca;
    11'b00001100111: data <= 32'hb49ea8ab;
    11'b00001101000: data <= 32'hbe69a62a;
    11'b00001101001: data <= 32'hbc323076;
    11'b00001101010: data <= 32'hb52b38b2;
    11'b00001101011: data <= 32'hbb59337d;
    11'b00001101100: data <= 32'hbf63bc84;
    11'b00001101101: data <= 32'hbd8fbf16;
    11'b00001101110: data <= 32'h30b4b587;
    11'b00001101111: data <= 32'h3c0d3f3a;
    11'b00001110000: data <= 32'h395d408c;
    11'b00001110001: data <= 32'h31d53bcb;
    11'b00001110010: data <= 32'h2f9a3032;
    11'b00001110011: data <= 32'hb1433a91;
    11'b00001110100: data <= 32'hba423dbd;
    11'b00001110101: data <= 32'hb85a35b5;
    11'b00001110110: data <= 32'h3c44bdbc;
    11'b00001110111: data <= 32'h40e7bf52;
    11'b00001111000: data <= 32'h3f92b94e;
    11'b00001111001: data <= 32'h317a35b0;
    11'b00001111010: data <= 32'hb77e3514;
    11'b00001111011: data <= 32'h351da161;
    11'b00001111100: data <= 32'h384aac9c;
    11'b00001111101: data <= 32'hbb4db814;
    11'b00001111110: data <= 32'hc0afbe35;
    11'b00001111111: data <= 32'hbf09bfc3;
    11'b00010000000: data <= 32'h3122b9d1;
    11'b00010000001: data <= 32'h3c613b2e;
    11'b00010000010: data <= 32'h359b3c81;
    11'b00010000011: data <= 32'hb90134a9;
    11'b00010000100: data <= 32'hba4735ab;
    11'b00010000101: data <= 32'hb9b43ebe;
    11'b00010000110: data <= 32'hbb89407f;
    11'b00010000111: data <= 32'hb9b8399a;
    11'b00010001000: data <= 32'h3828bd64;
    11'b00010001001: data <= 32'h3eb2bdf3;
    11'b00010001010: data <= 32'h3df3300b;
    11'b00010001011: data <= 32'h38fc3cfe;
    11'b00010001100: data <= 32'h39763a8b;
    11'b00010001101: data <= 32'h3deca40a;
    11'b00010001110: data <= 32'h3c94b304;
    11'b00010001111: data <= 32'hba43b629;
    11'b00010010000: data <= 32'hc052bcbb;
    11'b00010010001: data <= 32'hbcc2bf4e;
    11'b00010010010: data <= 32'h3b03bd65;
    11'b00010010011: data <= 32'h3dbab63c;
    11'b00010010100: data <= 32'h2e56b22d;
    11'b00010010101: data <= 32'hbc8cb6c1;
    11'b00010010110: data <= 32'hbc4a34f4;
    11'b00010010111: data <= 32'hb9843f3d;
    11'b00010011000: data <= 32'hbc194023;
    11'b00010011001: data <= 32'hbd8834ba;
    11'b00010011010: data <= 32'hb9dbbde5;
    11'b00010011011: data <= 32'h367dbc11;
    11'b00010011100: data <= 32'h3ad63b8e;
    11'b00010011101: data <= 32'h3a403f7b;
    11'b00010011110: data <= 32'h3cbc3c14;
    11'b00010011111: data <= 32'h3f0e2e77;
    11'b00010100000: data <= 32'h3c733521;
    11'b00010100001: data <= 32'hb9ae394e;
    11'b00010100010: data <= 32'hbe54b017;
    11'b00010100011: data <= 32'hb33cbdaa;
    11'b00010100100: data <= 32'h3ebbbf28;
    11'b00010100101: data <= 32'h3ee2bd12;
    11'b00010100110: data <= 32'h2de6bb2a;
    11'b00010100111: data <= 32'hbb32b9bb;
    11'b00010101000: data <= 32'hb6032f2e;
    11'b00010101001: data <= 32'h2b893d15;
    11'b00010101010: data <= 32'hbb0b3cb0;
    11'b00010101011: data <= 32'hc034b7e9;
    11'b00010101100: data <= 32'hbfb0bed8;
    11'b00010101101: data <= 32'hb8bfba4c;
    11'b00010101110: data <= 32'h360e3c72;
    11'b00010101111: data <= 32'h38c53e76;
    11'b00010110000: data <= 32'h3ab038d4;
    11'b00010110001: data <= 32'h3c793149;
    11'b00010110010: data <= 32'h38373cd3;
    11'b00010110011: data <= 32'hba384010;
    11'b00010110100: data <= 32'hbc673c0b;
    11'b00010110101: data <= 32'h355ebb79;
    11'b00010110110: data <= 32'h3f72bf22;
    11'b00010110111: data <= 32'h3e66bcfe;
    11'b00010111000: data <= 32'h33f2b8f9;
    11'b00010111001: data <= 32'ha817b70d;
    11'b00010111010: data <= 32'h3bcdaa1a;
    11'b00010111011: data <= 32'h3cb13891;
    11'b00010111100: data <= 32'hb8483535;
    11'b00010111101: data <= 32'hc0d0bbdf;
    11'b00010111110: data <= 32'hc0a8bf1d;
    11'b00010111111: data <= 32'hb9dfbb38;
    11'b00011000000: data <= 32'h35943744;
    11'b00011000001: data <= 32'h340637df;
    11'b00011000010: data <= 32'h22d5b54f;
    11'b00011000011: data <= 32'h30b42817;
    11'b00011000100: data <= 32'had673f6d;
    11'b00011000101: data <= 32'hbaf641c3;
    11'b00011000110: data <= 32'hbc303e2b;
    11'b00011000111: data <= 32'h25cdb97f;
    11'b00011001000: data <= 32'h3c77bd92;
    11'b00011001001: data <= 32'h3ba2b765;
    11'b00011001010: data <= 32'h356834d6;
    11'b00011001011: data <= 32'h3b1a2f0d;
    11'b00011001100: data <= 32'h4057addd;
    11'b00011001101: data <= 32'h400133c1;
    11'b00011001110: data <= 32'hb240338e;
    11'b00011001111: data <= 32'hc04bb94a;
    11'b00011010000: data <= 32'hbf1bbdc9;
    11'b00011010001: data <= 32'ha64fbcac;
    11'b00011010010: data <= 32'h39b5b8bc;
    11'b00011010011: data <= 32'ha56ebae7;
    11'b00011010100: data <= 32'hb91cbd2e;
    11'b00011010101: data <= 32'hb551b44e;
    11'b00011010110: data <= 32'hafc73f7e;
    11'b00011010111: data <= 32'hba254175;
    11'b00011011000: data <= 32'hbd833cbd;
    11'b00011011001: data <= 32'hbbdfba79;
    11'b00011011010: data <= 32'hb1e2bb3f;
    11'b00011011011: data <= 32'h2a843767;
    11'b00011011100: data <= 32'h32633c5d;
    11'b00011011101: data <= 32'h3d043624;
    11'b00011011110: data <= 32'h40fdafd0;
    11'b00011011111: data <= 32'h401f3794;
    11'b00011100000: data <= 32'had093c29;
    11'b00011100001: data <= 32'hbe3136a5;
    11'b00011100010: data <= 32'hb9deba0f;
    11'b00011100011: data <= 32'h3b5fbd1f;
    11'b00011100100: data <= 32'h3c51bd3f;
    11'b00011100101: data <= 32'hb079be79;
    11'b00011100110: data <= 32'hb969beea;
    11'b00011100111: data <= 32'h300ab875;
    11'b00011101000: data <= 32'h39113d35;
    11'b00011101001: data <= 32'hb59d3f1b;
    11'b00011101010: data <= 32'hbf01348d;
    11'b00011101011: data <= 32'hbffabc7d;
    11'b00011101100: data <= 32'hbcfdb8c0;
    11'b00011101101: data <= 32'hb8e63af9;
    11'b00011101110: data <= 32'hb01b3c44;
    11'b00011101111: data <= 32'h3adda536;
    11'b00011110000: data <= 32'h3f48b503;
    11'b00011110001: data <= 32'h3d9b3c0b;
    11'b00011110010: data <= 32'hb2cf406d;
    11'b00011110011: data <= 32'hbc073e7f;
    11'b00011110100: data <= 32'h2903aa12;
    11'b00011110101: data <= 32'h3d4abc52;
    11'b00011110110: data <= 32'h3beebce3;
    11'b00011110111: data <= 32'hb2d3bd5d;
    11'b00011111000: data <= 32'hb0d0bdb1;
    11'b00011111001: data <= 32'h3d18b960;
    11'b00011111010: data <= 32'h3f46387a;
    11'b00011111011: data <= 32'h340d39fd;
    11'b00011111100: data <= 32'hbf44b6b4;
    11'b00011111101: data <= 32'hc09fbcf9;
    11'b00011111110: data <= 32'hbda3b815;
    11'b00011111111: data <= 32'hb9503856;
    11'b00100000000: data <= 32'hb76330e3;
    11'b00100000001: data <= 32'h0c1abc16;
    11'b00100000010: data <= 32'h3994b9cb;
    11'b00100000011: data <= 32'h38b73d8a;
    11'b00100000100: data <= 32'hb60d41e8;
    11'b00100000101: data <= 32'hba4e4067;
    11'b00100000110: data <= 32'h28cf346c;
    11'b00100000111: data <= 32'h3a5cb942;
    11'b00100001000: data <= 32'h34a8b666;
    11'b00100001001: data <= 32'hb688b4bd;
    11'b00100001010: data <= 32'h3782b98e;
    11'b00100001011: data <= 32'h40b1b90d;
    11'b00100001100: data <= 32'h416e2e46;
    11'b00100001101: data <= 32'h39c935e2;
    11'b00100001110: data <= 32'hbde7b529;
    11'b00100001111: data <= 32'hbedabb05;
    11'b00100010000: data <= 32'hb8e0b7ee;
    11'b00100010001: data <= 32'hb0f1b203;
    11'b00100010010: data <= 32'hb935bc44;
    11'b00100010011: data <= 32'hba0fc025;
    11'b00100010100: data <= 32'haa93bcd1;
    11'b00100010101: data <= 32'h35163d18;
    11'b00100010110: data <= 32'hb44f417f;
    11'b00100010111: data <= 32'hbad53f24;
    11'b00100011000: data <= 32'hb9282a8a;
    11'b00100011001: data <= 32'hb5b7b3ab;
    11'b00100011010: data <= 32'hb9b338e3;
    11'b00100011011: data <= 32'hba2739e7;
    11'b00100011100: data <= 32'h3952b1da;
    11'b00100011101: data <= 32'h4137b91e;
    11'b00100011110: data <= 32'h41812dbc;
    11'b00100011111: data <= 32'h3a483ac4;
    11'b00100100000: data <= 32'hbb5e38b9;
    11'b00100100001: data <= 32'hb8c5ad7d;
    11'b00100100010: data <= 32'h3876b5a5;
    11'b00100100011: data <= 32'h3723b996;
    11'b00100100100: data <= 32'hb9c7bf05;
    11'b00100100101: data <= 32'hbc06c10a;
    11'b00100100110: data <= 32'h2d6dbdf9;
    11'b00100100111: data <= 32'h3b2139ba;
    11'b00100101000: data <= 32'h33b83eeb;
    11'b00100101001: data <= 32'hbb9e3984;
    11'b00100101010: data <= 32'hbda8b7c5;
    11'b00100101011: data <= 32'hbd622006;
    11'b00100101100: data <= 32'hbdb63cd1;
    11'b00100101101: data <= 32'hbc9f3c1e;
    11'b00100101110: data <= 32'h33d2b632;
    11'b00100101111: data <= 32'h3f7dbb3c;
    11'b00100110000: data <= 32'h3fb5358b;
    11'b00100110001: data <= 32'h372d3f03;
    11'b00100110010: data <= 32'hb73f3edc;
    11'b00100110011: data <= 32'h356b39aa;
    11'b00100110100: data <= 32'h3d11a8a0;
    11'b00100110101: data <= 32'h389ab85b;
    11'b00100110110: data <= 32'hbac0bdaf;
    11'b00100110111: data <= 32'hba09c02d;
    11'b00100111000: data <= 32'h3b99bdbf;
    11'b00100111001: data <= 32'h3fec29bc;
    11'b00100111010: data <= 32'h3b9b3874;
    11'b00100111011: data <= 32'hbacdb501;
    11'b00100111100: data <= 32'hbe7fbab9;
    11'b00100111101: data <= 32'hbdd42f33;
    11'b00100111110: data <= 32'hbd983c8d;
    11'b00100111111: data <= 32'hbd74368f;
    11'b00101000000: data <= 32'hb86dbd1c;
    11'b00101000001: data <= 32'h38fabdb9;
    11'b00101000010: data <= 32'h3aa2381c;
    11'b00101000011: data <= 32'h28b740b4;
    11'b00101000100: data <= 32'hb3ab407d;
    11'b00101000101: data <= 32'h38af3bfd;
    11'b00101000110: data <= 32'h3c2e3510;
    11'b00101000111: data <= 32'h1d6933ab;
    11'b00101001000: data <= 32'hbc9fb43f;
    11'b00101001001: data <= 32'hb5eabc62;
    11'b00101001010: data <= 32'h3f66bc97;
    11'b00101001011: data <= 32'h41aab632;
    11'b00101001100: data <= 32'h3dbaab44;
    11'b00101001101: data <= 32'hb82eb844;
    11'b00101001110: data <= 32'hbc25b909;
    11'b00101001111: data <= 32'hb87d3380;
    11'b00101010000: data <= 32'hb93f3948;
    11'b00101010001: data <= 32'hbd41b8e4;
    11'b00101010010: data <= 32'hbd0fc091;
    11'b00101010011: data <= 32'hb57abfdb;
    11'b00101010100: data <= 32'h336735c0;
    11'b00101010101: data <= 32'ha8f34040;
    11'b00101010110: data <= 32'hb2f63efc;
    11'b00101010111: data <= 32'h315538a0;
    11'b00101011000: data <= 32'h2f4e3828;
    11'b00101011001: data <= 32'hbb9d3ccb;
    11'b00101011010: data <= 32'hbe693bbe;
    11'b00101011011: data <= 32'hb449b413;
    11'b00101011100: data <= 32'h401fbb8a;
    11'b00101011101: data <= 32'h419ab755;
    11'b00101011110: data <= 32'h3d6030f0;
    11'b00101011111: data <= 32'hb0aa3042;
    11'b00101100000: data <= 32'h28252ea9;
    11'b00101100001: data <= 32'h3a5337ce;
    11'b00101100010: data <= 32'h345834a1;
    11'b00101100011: data <= 32'hbc9abce5;
    11'b00101100100: data <= 32'hbe32c15e;
    11'b00101100101: data <= 32'hb787c04d;
    11'b00101100110: data <= 32'h3845ac1d;
    11'b00101100111: data <= 32'h36473c91;
    11'b00101101000: data <= 32'hb23037b3;
    11'b00101101001: data <= 32'hb6cfb461;
    11'b00101101010: data <= 32'hba2f382b;
    11'b00101101011: data <= 32'hbe8b3f38;
    11'b00101101100: data <= 32'hbfc43e13;
    11'b00101101101: data <= 32'hb8d4b142;
    11'b00101101110: data <= 32'h3d64bc65;
    11'b00101101111: data <= 32'h3f4db525;
    11'b00101110000: data <= 32'h39b33ad9;
    11'b00101110001: data <= 32'h2cd63c84;
    11'b00101110010: data <= 32'h3bb83b07;
    11'b00101110011: data <= 32'h3f033a77;
    11'b00101110100: data <= 32'h39ba3691;
    11'b00101110101: data <= 32'hbc87bb2e;
    11'b00101110110: data <= 32'hbda0c03f;
    11'b00101110111: data <= 32'h315cbf54;
    11'b00101111000: data <= 32'h3ddeb7fe;
    11'b00101111001: data <= 32'h3c58a4c6;
    11'b00101111010: data <= 32'ha997ba2a;
    11'b00101111011: data <= 32'hb8efbbb3;
    11'b00101111100: data <= 32'hbaff3743;
    11'b00101111101: data <= 32'hbe073f52;
    11'b00101111110: data <= 32'hbfb73c8f;
    11'b00101111111: data <= 32'hbcc0baf8;
    11'b00110000000: data <= 32'h2f4ebe6a;
    11'b00110000001: data <= 32'h37c3b37b;
    11'b00110000010: data <= 32'ha9e43d8d;
    11'b00110000011: data <= 32'h2db13e87;
    11'b00110000100: data <= 32'h3d263c65;
    11'b00110000101: data <= 32'h3f243bf0;
    11'b00110000110: data <= 32'h35c43c0e;
    11'b00110000111: data <= 32'hbd9f33b7;
    11'b00110001000: data <= 32'hbc7bbb38;
    11'b00110001001: data <= 32'h3bb5bcc5;
    11'b00110001010: data <= 32'h408bb9ac;
    11'b00110001011: data <= 32'h3e18b989;
    11'b00110001100: data <= 32'h3177bd08;
    11'b00110001101: data <= 32'hb164bbfe;
    11'b00110001110: data <= 32'h1ec23820;
    11'b00110001111: data <= 32'hb8713dd9;
    11'b00110010000: data <= 32'hbe293417;
    11'b00110010001: data <= 32'hbea8bf40;
    11'b00110010010: data <= 32'hbb2ac03a;
    11'b00110010011: data <= 32'hb640b53b;
    11'b00110010100: data <= 32'hb67b3d07;
    11'b00110010101: data <= 32'h25603c92;
    11'b00110010110: data <= 32'h3bd837f6;
    11'b00110010111: data <= 32'h3c153b0d;
    11'b00110011000: data <= 32'hb8153ef3;
    11'b00110011001: data <= 32'hbf623e08;
    11'b00110011010: data <= 32'hbc033328;
    11'b00110011011: data <= 32'h3ce9b95e;
    11'b00110011100: data <= 32'h407eb93f;
    11'b00110011101: data <= 32'h3d25b8b8;
    11'b00110011110: data <= 32'h3451ba4b;
    11'b00110011111: data <= 32'h396fb614;
    11'b00110100000: data <= 32'h3d893a24;
    11'b00110100001: data <= 32'h393f3c76;
    11'b00110100010: data <= 32'hbc23b5ef;
    11'b00110100011: data <= 32'hbf2ac06d;
    11'b00110100100: data <= 32'hbc80c060;
    11'b00110100101: data <= 32'hb4fcb823;
    11'b00110100110: data <= 32'haff63792;
    11'b00110100111: data <= 32'h28e3b09a;
    11'b00110101000: data <= 32'h371db90e;
    11'b00110101001: data <= 32'h31023838;
    11'b00110101010: data <= 32'hbcc44052;
    11'b00110101011: data <= 32'hc036404d;
    11'b00110101100: data <= 32'hbc9e3881;
    11'b00110101101: data <= 32'h3980b915;
    11'b00110101110: data <= 32'h3d03b7e9;
    11'b00110101111: data <= 32'h3641283b;
    11'b00110110000: data <= 32'h305430d0;
    11'b00110110001: data <= 32'h3da63621;
    11'b00110110010: data <= 32'h40dd3c2d;
    11'b00110110011: data <= 32'h3d7e3c69;
    11'b00110110100: data <= 32'hba3fb20f;
    11'b00110110101: data <= 32'hbe62be93;
    11'b00110110110: data <= 32'hb8a0be82;
    11'b00110110111: data <= 32'h3835b8dd;
    11'b00110111000: data <= 32'h3853b7b2;
    11'b00110111001: data <= 32'h3170bde9;
    11'b00110111010: data <= 32'h3164be73;
    11'b00110111011: data <= 32'hab9f31f3;
    11'b00110111100: data <= 32'hbc404036;
    11'b00110111101: data <= 32'hbf8c3f7c;
    11'b00110111110: data <= 32'hbdaba249;
    11'b00110111111: data <= 32'hb573bc57;
    11'b00111000000: data <= 32'hb14ab670;
    11'b00111000001: data <= 32'hb96738da;
    11'b00111000010: data <= 32'hb12239e1;
    11'b00111000011: data <= 32'h3e8138e8;
    11'b00111000100: data <= 32'h41233c3f;
    11'b00111000101: data <= 32'h3cbd3dad;
    11'b00111000110: data <= 32'hbbbc3a01;
    11'b00111000111: data <= 32'hbd3bb59d;
    11'b00111001000: data <= 32'h3324b962;
    11'b00111001001: data <= 32'h3d87b7b5;
    11'b00111001010: data <= 32'h3bf5bc16;
    11'b00111001011: data <= 32'h342ac026;
    11'b00111001100: data <= 32'h35f7bf6b;
    11'b00111001101: data <= 32'h39162fb0;
    11'b00111001110: data <= 32'haac13ee8;
    11'b00111001111: data <= 32'hbcc23c08;
    11'b00111010000: data <= 32'hbe2bbbc8;
    11'b00111010001: data <= 32'hbccbbe72;
    11'b00111010010: data <= 32'hbca2b68e;
    11'b00111010011: data <= 32'hbd1d3964;
    11'b00111010100: data <= 32'hb66736a5;
    11'b00111010101: data <= 32'h3d2da7ef;
    11'b00111010110: data <= 32'h3f65394d;
    11'b00111010111: data <= 32'h35413f29;
    11'b00111011000: data <= 32'hbdaa3f68;
    11'b00111011001: data <= 32'hbc8b3b2c;
    11'b00111011010: data <= 32'h39273025;
    11'b00111011011: data <= 32'h3e06b2b7;
    11'b00111011100: data <= 32'h39d9bb02;
    11'b00111011101: data <= 32'h2e7ebeaf;
    11'b00111011110: data <= 32'h3b0dbd27;
    11'b00111011111: data <= 32'h3f5d35df;
    11'b00111100000: data <= 32'h3d1e3d64;
    11'b00111100001: data <= 32'hb6003437;
    11'b00111100010: data <= 32'hbda0be05;
    11'b00111100011: data <= 32'hbd72beb6;
    11'b00111100100: data <= 32'hbcacb60e;
    11'b00111100101: data <= 32'hbc623296;
    11'b00111100110: data <= 32'hb6a1b996;
    11'b00111100111: data <= 32'h39ebbd1b;
    11'b00111101000: data <= 32'h3b38a424;
    11'b00111101001: data <= 32'hb7783fab;
    11'b00111101010: data <= 32'hbec040d0;
    11'b00111101011: data <= 32'hbc6b3d60;
    11'b00111101100: data <= 32'h364134fe;
    11'b00111101101: data <= 32'h3977253a;
    11'b00111101110: data <= 32'hb456b3a8;
    11'b00111101111: data <= 32'hb5cab97c;
    11'b00111110000: data <= 32'h3d2eb6f2;
    11'b00111110001: data <= 32'h41923958;
    11'b00111110010: data <= 32'h403e3cc5;
    11'b00111110011: data <= 32'h2cbf320d;
    11'b00111110100: data <= 32'hbc64bc6a;
    11'b00111110101: data <= 32'hba60bc1b;
    11'b00111110110: data <= 32'hb508b0bd;
    11'b00111110111: data <= 32'hb5edb6b2;
    11'b00111111000: data <= 32'hb409bfab;
    11'b00111111001: data <= 32'h35bcc0cb;
    11'b00111111010: data <= 32'h3768b8ca;
    11'b00111111011: data <= 32'hb80b3ece;
    11'b00111111100: data <= 32'hbd9a4032;
    11'b00111111101: data <= 32'hbc423a44;
    11'b00111111110: data <= 32'hb4e7b118;
    11'b00111111111: data <= 32'hb8e72db8;
    11'b01000000000: data <= 32'hbdf5368f;
    11'b01000000001: data <= 32'hbb802da7;
    11'b01000000010: data <= 32'h3d3aa90c;
    11'b01000000011: data <= 32'h41c3392d;
    11'b01000000100: data <= 32'h3fea3cf2;
    11'b01000000101: data <= 32'had9f3a70;
    11'b01000000110: data <= 32'hba812b7b;
    11'b01000000111: data <= 32'h2bc12d6f;
    11'b01000001000: data <= 32'h3994349f;
    11'b01000001001: data <= 32'h33afb9c5;
    11'b01000001010: data <= 32'hb18bc0ef;
    11'b01000001011: data <= 32'h353ac16f;
    11'b01000001100: data <= 32'h3ac9b9e8;
    11'b01000001101: data <= 32'h35d63d30;
    11'b01000001110: data <= 32'hb8693cc3;
    11'b01000001111: data <= 32'hbae2b4d2;
    11'b01000010000: data <= 32'hbb2bbaa0;
    11'b01000010001: data <= 32'hbe332c9b;
    11'b01000010010: data <= 32'hc0683966;
    11'b01000010011: data <= 32'hbd382ba0;
    11'b01000010100: data <= 32'h3b51b845;
    11'b01000010101: data <= 32'h403f2f35;
    11'b01000010110: data <= 32'h3c1f3d19;
    11'b01000010111: data <= 32'hb9443e77;
    11'b01000011000: data <= 32'hb94f3cf8;
    11'b01000011001: data <= 32'h392a3c1e;
    11'b01000011010: data <= 32'h3c5d39f2;
    11'b01000011011: data <= 32'h3059b79d;
    11'b01000011100: data <= 32'hb714c00e;
    11'b01000011101: data <= 32'h3818c030;
    11'b01000011110: data <= 32'h3f01b669;
    11'b01000011111: data <= 32'h3e803b8c;
    11'b01000100000: data <= 32'h36d934f5;
    11'b01000100001: data <= 32'hb7ddbc54;
    11'b01000100010: data <= 32'hbb5dbc3e;
    11'b01000100011: data <= 32'hbe1d31ea;
    11'b01000100100: data <= 32'hc0033815;
    11'b01000100101: data <= 32'hbd13b9fe;
    11'b01000100110: data <= 32'h3610beca;
    11'b01000100111: data <= 32'h3c40b9f3;
    11'b01000101000: data <= 32'h204f3c81;
    11'b01000101001: data <= 32'hbc693ffb;
    11'b01000101010: data <= 32'hb8a43ea5;
    11'b01000101011: data <= 32'h395d3cf7;
    11'b01000101100: data <= 32'h38923bca;
    11'b01000101101: data <= 32'hba2c3118;
    11'b01000101110: data <= 32'hbc56bb98;
    11'b01000101111: data <= 32'h38febc27;
    11'b01000110000: data <= 32'h40f92ccb;
    11'b01000110001: data <= 32'h40e13a1a;
    11'b01000110010: data <= 32'h3b9ea422;
    11'b01000110011: data <= 32'hb009bbd9;
    11'b01000110100: data <= 32'hb549b828;
    11'b01000110101: data <= 32'hb8cc38b0;
    11'b01000110110: data <= 32'hbc713274;
    11'b01000110111: data <= 32'hbb87bef2;
    11'b01000111000: data <= 32'h9e21c195;
    11'b01000111001: data <= 32'h3660bdc4;
    11'b01000111010: data <= 32'hb53c3a5e;
    11'b01000111011: data <= 32'hbb8e3e84;
    11'b01000111100: data <= 32'hb6313c29;
    11'b01000111101: data <= 32'h34b03920;
    11'b01000111110: data <= 32'hb79e3b31;
    11'b01000111111: data <= 32'hbfdb3a63;
    11'b01001000000: data <= 32'hbf3d25fe;
    11'b01001000001: data <= 32'h377fb5a6;
    11'b01001000010: data <= 32'h40fd328c;
    11'b01001000011: data <= 32'h4080396f;
    11'b01001000100: data <= 32'h39a43489;
    11'b01001000101: data <= 32'h2a84ad34;
    11'b01001000110: data <= 32'h3820387c;
    11'b01001000111: data <= 32'h38b13cca;
    11'b01001001000: data <= 32'hb3112f26;
    11'b01001001001: data <= 32'hb988c056;
    11'b01001001010: data <= 32'hb04dc228;
    11'b01001001011: data <= 32'h37a9be2e;
    11'b01001001100: data <= 32'h34453748;
    11'b01001001101: data <= 32'hb07339c8;
    11'b01001001110: data <= 32'h200eb24e;
    11'b01001001111: data <= 32'ha9f8b4a2;
    11'b01001010000: data <= 32'hbd14399a;
    11'b01001010001: data <= 32'hc1523c86;
    11'b01001010010: data <= 32'hc0623487;
    11'b01001010011: data <= 32'h2dbab878;
    11'b01001010100: data <= 32'h3ee3b43e;
    11'b01001010101: data <= 32'h3cad3833;
    11'b01001010110: data <= 32'hae873a89;
    11'b01001010111: data <= 32'h24d63b7e;
    11'b01001011000: data <= 32'h3c943e03;
    11'b01001011001: data <= 32'h3d003ee0;
    11'b01001011010: data <= 32'ha6de365a;
    11'b01001011011: data <= 32'hbaf5beca;
    11'b01001011100: data <= 32'hb026c0b0;
    11'b01001011101: data <= 32'h3c59bc03;
    11'b01001011110: data <= 32'h3d5b3458;
    11'b01001011111: data <= 32'h3ac7b1f8;
    11'b01001100000: data <= 32'h37dcbced;
    11'b01001100001: data <= 32'h25beba9e;
    11'b01001100010: data <= 32'hbccc3990;
    11'b01001100011: data <= 32'hc0c13c81;
    11'b01001100100: data <= 32'hbff9b329;
    11'b01001100101: data <= 32'hb4c4be0d;
    11'b01001100110: data <= 32'h3920bc83;
    11'b01001100111: data <= 32'hadd93337;
    11'b01001101000: data <= 32'hbad63c35;
    11'b01001101001: data <= 32'ha91b3d26;
    11'b01001101010: data <= 32'h3d393ea4;
    11'b01001101011: data <= 32'h3c223f5b;
    11'b01001101100: data <= 32'hb9a33b56;
    11'b01001101101: data <= 32'hbe09b8cd;
    11'b01001101110: data <= 32'hb22abc46;
    11'b01001101111: data <= 32'h3e8db31b;
    11'b01001110000: data <= 32'h4021340e;
    11'b01001110001: data <= 32'h3d60b904;
    11'b01001110010: data <= 32'h3a6ebdbb;
    11'b01001110011: data <= 32'h3851b84a;
    11'b01001110100: data <= 32'hb3fe3c4e;
    11'b01001110101: data <= 32'hbd253c03;
    11'b01001110110: data <= 32'hbd7ebbf3;
    11'b01001110111: data <= 32'hb80fc100;
    11'b01001111000: data <= 32'haf8abf4a;
    11'b01001111001: data <= 32'hb9d3aeff;
    11'b01001111010: data <= 32'hbbc239b0;
    11'b01001111011: data <= 32'h2f05391c;
    11'b01001111100: data <= 32'h3c763b1f;
    11'b01001111101: data <= 32'h334a3dfe;
    11'b01001111110: data <= 32'hbf163d84;
    11'b01001111111: data <= 32'hc07f372e;
    11'b01010000000: data <= 32'hb679ad6e;
    11'b01010000001: data <= 32'h3e7b3289;
    11'b01010000010: data <= 32'h3f5c33bf;
    11'b01010000011: data <= 32'h3bb0b810;
    11'b01010000100: data <= 32'h3a07ba5b;
    11'b01010000101: data <= 32'h3ce23664;
    11'b01010000110: data <= 32'h3bff3edc;
    11'b01010000111: data <= 32'haebd3c0d;
    11'b01010001000: data <= 32'hba77bd6d;
    11'b01010001001: data <= 32'hb842c17d;
    11'b01010001010: data <= 32'hb298bf4d;
    11'b01010001011: data <= 32'hb69fb457;
    11'b01010001100: data <= 32'hb555aaef;
    11'b01010001101: data <= 32'h3842b93b;
    11'b01010001110: data <= 32'h3b49b515;
    11'b01010001111: data <= 32'hb7593bcd;
    11'b01010010000: data <= 32'hc0d73e52;
    11'b01010010001: data <= 32'hc1223ae4;
    11'b01010010010: data <= 32'hb9431cef;
    11'b01010010011: data <= 32'h3ba8ac35;
    11'b01010010100: data <= 32'h39a82c81;
    11'b01010010101: data <= 32'haeb4b046;
    11'b01010010110: data <= 32'h36682d31;
    11'b01010010111: data <= 32'h3ecc3d25;
    11'b01010011000: data <= 32'h3f34406b;
    11'b01010011001: data <= 32'h36583ce9;
    11'b01010011010: data <= 32'hba06bbaf;
    11'b01010011011: data <= 32'hb830bfd9;
    11'b01010011100: data <= 32'h3356bc32;
    11'b01010011101: data <= 32'h37bbb0c4;
    11'b01010011110: data <= 32'h38b0ba74;
    11'b01010011111: data <= 32'h3c15bf41;
    11'b01010100000: data <= 32'h3bb6bcb0;
    11'b01010100001: data <= 32'hb6d339a1;
    11'b01010100010: data <= 32'hc0303e2c;
    11'b01010100011: data <= 32'hc0563840;
    11'b01010100100: data <= 32'hba21b9f3;
    11'b01010100101: data <= 32'h27cababe;
    11'b01010100110: data <= 32'hb95ab418;
    11'b01010100111: data <= 32'hbcb82c44;
    11'b01010101000: data <= 32'h2a1d36f0;
    11'b01010101001: data <= 32'h3f343da2;
    11'b01010101010: data <= 32'h3f0a4056;
    11'b01010101011: data <= 32'haa343e07;
    11'b01010101100: data <= 32'hbd1f9f71;
    11'b01010101101: data <= 32'hb8fab89e;
    11'b01010101110: data <= 32'h39a02af1;
    11'b01010101111: data <= 32'h3cb430bb;
    11'b01010110000: data <= 32'h3c38bca5;
    11'b01010110001: data <= 32'h3ce1c060;
    11'b01010110010: data <= 32'h3d26bc90;
    11'b01010110011: data <= 32'h36543b8a;
    11'b01010110100: data <= 32'hbb3e3dd0;
    11'b01010110101: data <= 32'hbcefb02c;
    11'b01010110110: data <= 32'hb931bea7;
    11'b01010110111: data <= 32'hb8fabe0c;
    11'b01010111000: data <= 32'hbde9b82d;
    11'b01010111001: data <= 32'hbe53b04b;
    11'b01010111010: data <= 32'h24f0af04;
    11'b01010111011: data <= 32'h3e863870;
    11'b01010111100: data <= 32'h3c563e24;
    11'b01010111101: data <= 32'hbc103e92;
    11'b01010111110: data <= 32'hbff73b5f;
    11'b01010111111: data <= 32'hba6e389c;
    11'b01011000000: data <= 32'h3a2f3a5a;
    11'b01011000001: data <= 32'h3c1d35a5;
    11'b01011000010: data <= 32'h38d5bc2e;
    11'b01011000011: data <= 32'h3b46bec9;
    11'b01011000100: data <= 32'h3ea2b562;
    11'b01011000101: data <= 32'h3e123e2a;
    11'b01011000110: data <= 32'h370f3dd9;
    11'b01011000111: data <= 32'hb557b844;
    11'b01011001000: data <= 32'hb6b5bfd7;
    11'b01011001001: data <= 32'hb989bdda;
    11'b01011001010: data <= 32'hbd4db771;
    11'b01011001011: data <= 32'hbc72b8f3;
    11'b01011001100: data <= 32'h362abd1b;
    11'b01011001101: data <= 32'h3dc7ba7c;
    11'b01011001110: data <= 32'h365d3951;
    11'b01011001111: data <= 32'hbec53e3a;
    11'b01011010000: data <= 32'hc08d3d2c;
    11'b01011010001: data <= 32'hbb103abc;
    11'b01011010010: data <= 32'h35a639d6;
    11'b01011010011: data <= 32'h23733441;
    11'b01011010100: data <= 32'hb8deb99a;
    11'b01011010101: data <= 32'h32b0badd;
    11'b01011010110: data <= 32'h3f513871;
    11'b01011010111: data <= 32'h40844008;
    11'b01011011000: data <= 32'h3c843e31;
    11'b01011011001: data <= 32'ha804b56c;
    11'b01011011010: data <= 32'hb49ebd24;
    11'b01011011011: data <= 32'hb493b870;
    11'b01011011100: data <= 32'hb7fca006;
    11'b01011011101: data <= 32'hb2debc38;
    11'b01011011110: data <= 32'h3aebc0b8;
    11'b01011011111: data <= 32'h3da7bf70;
    11'b01011100000: data <= 32'h34542ee6;
    11'b01011100001: data <= 32'hbddd3d6d;
    11'b01011100010: data <= 32'hbf0e3bde;
    11'b01011100011: data <= 32'hb96f3229;
    11'b01011100100: data <= 32'hb4322081;
    11'b01011100101: data <= 32'hbd1daabb;
    11'b01011100110: data <= 32'hbf89b744;
    11'b01011100111: data <= 32'hb762b635;
    11'b01011101000: data <= 32'h3ee73a21;
    11'b01011101001: data <= 32'h40713f90;
    11'b01011101010: data <= 32'h3a7a3e31;
    11'b01011101011: data <= 32'hb7693512;
    11'b01011101100: data <= 32'hb5e12274;
    11'b01011101101: data <= 32'h328c3a03;
    11'b01011101110: data <= 32'h3453390d;
    11'b01011101111: data <= 32'h354cbcaf;
    11'b01011110000: data <= 32'h3c06c174;
    11'b01011110001: data <= 32'h3e00bfe9;
    11'b01011110010: data <= 32'h3a8a329c;
    11'b01011110011: data <= 32'hb5d63ce4;
    11'b01011110100: data <= 32'hb90b3528;
    11'b01011110101: data <= 32'hb28dba20;
    11'b01011110110: data <= 32'hb932b9c4;
    11'b01011110111: data <= 32'hc023b499;
    11'b01011111000: data <= 32'hc0ebb770;
    11'b01011111001: data <= 32'hb967b979;
    11'b01011111010: data <= 32'h3ded1d5b;
    11'b01011111011: data <= 32'h3e393c49;
    11'b01011111100: data <= 32'hb12b3d4c;
    11'b01011111101: data <= 32'hbcda3bb2;
    11'b01011111110: data <= 32'hb84a3c90;
    11'b01011111111: data <= 32'h36b63ec3;
    11'b01100000000: data <= 32'h35683c47;
    11'b01100000001: data <= 32'ha615bb91;
    11'b01100000010: data <= 32'h3849c07f;
    11'b01100000011: data <= 32'h3e19bccf;
    11'b01100000100: data <= 32'h3e963a8b;
    11'b01100000101: data <= 32'h3b973ce8;
    11'b01100000110: data <= 32'h37d6b1f9;
    11'b01100000111: data <= 32'h34dbbcf9;
    11'b01100001000: data <= 32'hb895ba28;
    11'b01100001001: data <= 32'hbfbaae6f;
    11'b01100001010: data <= 32'hc01cb908;
    11'b01100001011: data <= 32'hb550be3e;
    11'b01100001100: data <= 32'h3d28bd47;
    11'b01100001101: data <= 32'h3a5ba7f0;
    11'b01100001110: data <= 32'hbbe83b5e;
    11'b01100001111: data <= 32'hbe603c99;
    11'b01100010000: data <= 32'hb8233dae;
    11'b01100010001: data <= 32'h34903eeb;
    11'b01100010010: data <= 32'hb65a3c31;
    11'b01100010011: data <= 32'hbcc0b8ab;
    11'b01100010100: data <= 32'hb65ebd70;
    11'b01100010101: data <= 32'h3d67b222;
    11'b01100010110: data <= 32'h40583d8d;
    11'b01100010111: data <= 32'h3e993cfb;
    11'b01100011000: data <= 32'h3b7cb3b4;
    11'b01100011001: data <= 32'h3868baa9;
    11'b01100011010: data <= 32'hb01f2d34;
    11'b01100011011: data <= 32'hbc4c38a6;
    11'b01100011100: data <= 32'hbc49b9ae;
    11'b01100011101: data <= 32'h3382c0d0;
    11'b01100011110: data <= 32'h3cdfc0c2;
    11'b01100011111: data <= 32'h374cba26;
    11'b01100100000: data <= 32'hbc083864;
    11'b01100100001: data <= 32'hbc9a3a30;
    11'b01100100010: data <= 32'haed93a10;
    11'b01100100011: data <= 32'h25f63bb0;
    11'b01100100100: data <= 32'hbdc23947;
    11'b01100100101: data <= 32'hc0f2b513;
    11'b01100100110: data <= 32'hbd1fb9b7;
    11'b01100100111: data <= 32'h3c193400;
    11'b01100101000: data <= 32'h40133d61;
    11'b01100101001: data <= 32'h3d513c42;
    11'b01100101010: data <= 32'h37fa2cb1;
    11'b01100101011: data <= 32'h36ec32b1;
    11'b01100101100: data <= 32'h35f53d95;
    11'b01100101101: data <= 32'hb1413dd3;
    11'b01100101110: data <= 32'hb506b879;
    11'b01100101111: data <= 32'h3798c149;
    11'b01100110000: data <= 32'h3ca0c104;
    11'b01100110001: data <= 32'h3972b9ae;
    11'b01100110010: data <= 32'hb156369f;
    11'b01100110011: data <= 32'ha4192e56;
    11'b01100110100: data <= 32'h38f2b4ff;
    11'b01100110101: data <= 32'habf9298e;
    11'b01100110110: data <= 32'hc025350e;
    11'b01100110111: data <= 32'hc224b2e7;
    11'b01100111000: data <= 32'hbe54b9b8;
    11'b01100111001: data <= 32'h39d8b401;
    11'b01100111010: data <= 32'h3d60384c;
    11'b01100111011: data <= 32'h345638b4;
    11'b01100111100: data <= 32'hb6903647;
    11'b01100111101: data <= 32'h30e83ca3;
    11'b01100111110: data <= 32'h395740bc;
    11'b01100111111: data <= 32'h3169400f;
    11'b01101000000: data <= 32'hb68cb372;
    11'b01101000001: data <= 32'h2881c03d;
    11'b01101000010: data <= 32'h3b80beac;
    11'b01101000011: data <= 32'h3caf269e;
    11'b01101000100: data <= 32'h3b9e3827;
    11'b01101000101: data <= 32'h3c98b776;
    11'b01101000110: data <= 32'h3d3bbc1a;
    11'b01101000111: data <= 32'h3159b42c;
    11'b01101001000: data <= 32'hbf7c372c;
    11'b01101001001: data <= 32'hc13fb118;
    11'b01101001010: data <= 32'hbc9ebd00;
    11'b01101001011: data <= 32'h38f5bd76;
    11'b01101001100: data <= 32'h3852b8ea;
    11'b01101001101: data <= 32'hba1da87f;
    11'b01101001110: data <= 32'hbc28360e;
    11'b01101001111: data <= 32'h2e193d6b;
    11'b01101010000: data <= 32'h39cb40c9;
    11'b01101010001: data <= 32'hb3773fe3;
    11'b01101010010: data <= 32'hbd672d02;
    11'b01101010011: data <= 32'hbb8bbcc7;
    11'b01101010100: data <= 32'h3827b791;
    11'b01101010101: data <= 32'h3dce3aaa;
    11'b01101010110: data <= 32'h3e323911;
    11'b01101010111: data <= 32'h3e6db972;
    11'b01101011000: data <= 32'h3e4bbb77;
    11'b01101011001: data <= 32'h38cc35b8;
    11'b01101011010: data <= 32'hbbd53ca5;
    11'b01101011011: data <= 32'hbded2443;
    11'b01101011100: data <= 32'hb5dbbf46;
    11'b01101011101: data <= 32'h3940c09b;
    11'b01101011110: data <= 32'h2c76bd8d;
    11'b01101011111: data <= 32'hbc59b7bb;
    11'b01101100000: data <= 32'hbab6a861;
    11'b01101100001: data <= 32'h38253938;
    11'b01101100010: data <= 32'h39bf3dfa;
    11'b01101100011: data <= 32'hbbd33d8d;
    11'b01101100100: data <= 32'hc0fe336f;
    11'b01101100101: data <= 32'hbf86b710;
    11'b01101100110: data <= 32'h2c00341c;
    11'b01101100111: data <= 32'h3cea3c2d;
    11'b01101101000: data <= 32'h3cb7376b;
    11'b01101101001: data <= 32'h3c4bb8e6;
    11'b01101101010: data <= 32'h3d30b272;
    11'b01101101011: data <= 32'h3bf83e13;
    11'b01101101100: data <= 32'h24df4036;
    11'b01101101101: data <= 32'hb740357d;
    11'b01101101110: data <= 32'h3069bfae;
    11'b01101101111: data <= 32'h3912c0be;
    11'b01101110000: data <= 32'h2c3dbd14;
    11'b01101110001: data <= 32'hb880b812;
    11'b01101110010: data <= 32'h301eb900;
    11'b01101110011: data <= 32'h3d46b7db;
    11'b01101110100: data <= 32'h3abf3537;
    11'b01101110101: data <= 32'hbdbf3a34;
    11'b01101110110: data <= 32'hc20d3445;
    11'b01101110111: data <= 32'hc051b38f;
    11'b01101111000: data <= 32'hb1ac2cf2;
    11'b01101111001: data <= 32'h38b236c4;
    11'b01101111010: data <= 32'h2b1dad65;
    11'b01101111011: data <= 32'habd9b83b;
    11'b01101111100: data <= 32'h3a0b3853;
    11'b01101111101: data <= 32'h3ccf40d5;
    11'b01101111110: data <= 32'h38444161;
    11'b01101111111: data <= 32'hb3423961;
    11'b01110000000: data <= 32'hade4bda3;
    11'b01110000001: data <= 32'h35c0bde0;
    11'b01110000010: data <= 32'h34e9b560;
    11'b01110000011: data <= 32'h3519b117;
    11'b01110000100: data <= 32'h3cd7bc5c;
    11'b01110000101: data <= 32'h401bbd73;
    11'b01110000110: data <= 32'h3c87b4c0;
    11'b01110000111: data <= 32'hbcd43964;
    11'b01110001000: data <= 32'hc10935ab;
    11'b01110001001: data <= 32'hbe44b828;
    11'b01110001010: data <= 32'haca7ba36;
    11'b01110001011: data <= 32'haf7cb912;
    11'b01110001100: data <= 32'hbc7bba3c;
    11'b01110001101: data <= 32'hbc03b93e;
    11'b01110001110: data <= 32'h3716395c;
    11'b01110001111: data <= 32'h3d0a40c5;
    11'b01110010000: data <= 32'h35ff4104;
    11'b01110010001: data <= 32'hbb1a3a75;
    11'b01110010010: data <= 32'hbba9b897;
    11'b01110010011: data <= 32'hb0b5b0b0;
    11'b01110010100: data <= 32'h36da3a33;
    11'b01110010101: data <= 32'h3a80332b;
    11'b01110010110: data <= 32'h3e7abd1d;
    11'b01110010111: data <= 32'h407abe01;
    11'b01110011000: data <= 32'h3dbf2669;
    11'b01110011001: data <= 32'hb62c3d02;
    11'b01110011010: data <= 32'hbd0c38f6;
    11'b01110011011: data <= 32'hb7cfbb29;
    11'b01110011100: data <= 32'h33acbe4d;
    11'b01110011101: data <= 32'hb84ebd73;
    11'b01110011110: data <= 32'hbea5bcc9;
    11'b01110011111: data <= 32'hbc73bbf8;
    11'b01110100000: data <= 32'h39a2230a;
    11'b01110100001: data <= 32'h3d573d8a;
    11'b01110100010: data <= 32'hb0f13ea0;
    11'b01110100011: data <= 32'hbf763981;
    11'b01110100100: data <= 32'hbf672f44;
    11'b01110100101: data <= 32'hb8ef3a53;
    11'b01110100110: data <= 32'h33093d3c;
    11'b01110100111: data <= 32'h375e33da;
    11'b01110101000: data <= 32'h3bffbd18;
    11'b01110101001: data <= 32'h3eebbbfb;
    11'b01110101010: data <= 32'h3e4e3bed;
    11'b01110101011: data <= 32'h384c404a;
    11'b01110101100: data <= 32'ha8b63bf5;
    11'b01110101101: data <= 32'h359cbba4;
    11'b01110101110: data <= 32'h3706be85;
    11'b01110101111: data <= 32'hb8adbcb1;
    11'b01110110000: data <= 32'hbd7dbc21;
    11'b01110110001: data <= 32'hb5dbbd71;
    11'b01110110010: data <= 32'h3dc4bc37;
    11'b01110110011: data <= 32'h3e22282c;
    11'b01110110100: data <= 32'hb83339a1;
    11'b01110110101: data <= 32'hc0b33793;
    11'b01110110110: data <= 32'hc0253566;
    11'b01110110111: data <= 32'hb9b93ace;
    11'b01110111000: data <= 32'hb39c3b7d;
    11'b01110111001: data <= 32'hb8c4b31b;
    11'b01110111010: data <= 32'hb4e0bd1c;
    11'b01110111011: data <= 32'h3ad1b61c;
    11'b01110111100: data <= 32'h3e0d3f46;
    11'b01110111101: data <= 32'h3c2f4161;
    11'b01110111110: data <= 32'h36e63cee;
    11'b01110111111: data <= 32'h3660b8a5;
    11'b01111000000: data <= 32'h345bba3f;
    11'b01111000001: data <= 32'hb6f7ad94;
    11'b01111000010: data <= 32'hb931b5cf;
    11'b01111000011: data <= 32'h38f8be33;
    11'b01111000100: data <= 32'h404cbf9a;
    11'b01111000101: data <= 32'h3f1ebaa5;
    11'b01111000110: data <= 32'hb61c34bb;
    11'b01111000111: data <= 32'hbf8436b0;
    11'b01111001000: data <= 32'hbd633071;
    11'b01111001001: data <= 32'hb51831cf;
    11'b01111001010: data <= 32'hb96214d0;
    11'b01111001011: data <= 32'hbef1bb2d;
    11'b01111001100: data <= 32'hbdefbda0;
    11'b01111001101: data <= 32'h32b0b2de;
    11'b01111001110: data <= 32'h3d913f3b;
    11'b01111001111: data <= 32'h3ba940cb;
    11'b01111010000: data <= 32'ha6203c72;
    11'b01111010001: data <= 32'hb5031d83;
    11'b01111010010: data <= 32'hb2c33803;
    11'b01111010011: data <= 32'hb5a33d07;
    11'b01111010100: data <= 32'hb13c35e3;
    11'b01111010101: data <= 32'h3c24be1a;
    11'b01111010110: data <= 32'h4082c02e;
    11'b01111010111: data <= 32'h3f7eb9d9;
    11'b01111011000: data <= 32'h32f5397a;
    11'b01111011001: data <= 32'hb94b392a;
    11'b01111011010: data <= 32'ha989b18a;
    11'b01111011011: data <= 32'h359bb888;
    11'b01111011100: data <= 32'hbadcb9bb;
    11'b01111011101: data <= 32'hc0a0bd0b;
    11'b01111011110: data <= 32'hbf51be59;
    11'b01111011111: data <= 32'h33cdb977;
    11'b01111100000: data <= 32'h3d9d3ac3;
    11'b01111100001: data <= 32'h38093d56;
    11'b01111100010: data <= 32'hbb4d391b;
    11'b01111100011: data <= 32'hbcb3370b;
    11'b01111100100: data <= 32'hb9363dd9;
    11'b01111100101: data <= 32'hb7474015;
    11'b01111100110: data <= 32'hb5e43939;
    11'b01111100111: data <= 32'h373cbdb5;
    11'b01111101000: data <= 32'h3e38beaa;
    11'b01111101001: data <= 32'h3eb12f52;
    11'b01111101010: data <= 32'h3b0e3e16;
    11'b01111101011: data <= 32'h389e3c06;
    11'b01111101100: data <= 32'h3c3cb4a5;
    11'b01111101101: data <= 32'h3accb9cf;
    11'b01111101110: data <= 32'hba35b87c;
    11'b01111101111: data <= 32'hc033bb83;
    11'b01111110000: data <= 32'hbceebe91;
    11'b01111110001: data <= 32'h3b2dbdfd;
    11'b01111110010: data <= 32'h3e5eb81b;
    11'b01111110011: data <= 32'h2f712efc;
    11'b01111110100: data <= 32'hbdd92dd4;
    11'b01111110101: data <= 32'hbdb43806;
    11'b01111110110: data <= 32'hb9043e61;
    11'b01111110111: data <= 32'hb9253f63;
    11'b01111111000: data <= 32'hbcbf34df;
    11'b01111111001: data <= 32'hbad0bdaa;
    11'b01111111010: data <= 32'h3680bc41;
    11'b01111111011: data <= 32'h3d043bc2;
    11'b01111111100: data <= 32'h3ccc402d;
    11'b01111111101: data <= 32'h3c743c9f;
    11'b01111111110: data <= 32'h3d45b069;
    11'b01111111111: data <= 32'h3abfadc5;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    