
module memory_rom_56(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h38e4bdd1;
    11'b00000000001: data <= 32'h34c2bb29;
    11'b00000000010: data <= 32'hb5ac3a6e;
    11'b00000000011: data <= 32'hbd903d00;
    11'b00000000100: data <= 32'hbea6b709;
    11'b00000000101: data <= 32'hba72c064;
    11'b00000000110: data <= 32'haf98bf8a;
    11'b00000000111: data <= 32'hb82ab05e;
    11'b00000001000: data <= 32'hbb7f3bc1;
    11'b00000001001: data <= 32'hac8b3b92;
    11'b00000001010: data <= 32'h3ca63bd5;
    11'b00000001011: data <= 32'h39f33def;
    11'b00000001100: data <= 32'hbcc03de3;
    11'b00000001101: data <= 32'hc03a3851;
    11'b00000001110: data <= 32'hb900b35c;
    11'b00000001111: data <= 32'h3e4aad42;
    11'b00000010000: data <= 32'h40432ef5;
    11'b00000010001: data <= 32'h3cd5b82b;
    11'b00000010010: data <= 32'h393dbc28;
    11'b00000010011: data <= 32'h3bd0b039;
    11'b00000010100: data <= 32'h3b463d6c;
    11'b00000010101: data <= 32'hb0113caf;
    11'b00000010110: data <= 32'hbc0cbbeb;
    11'b00000010111: data <= 32'hbae6c167;
    11'b00000011000: data <= 32'hb681c02f;
    11'b00000011001: data <= 32'hb7e8b578;
    11'b00000011010: data <= 32'hb84d34b2;
    11'b00000011011: data <= 32'h3377b3ee;
    11'b00000011100: data <= 32'h3b28b275;
    11'b00000011101: data <= 32'hab2c3bac;
    11'b00000011110: data <= 32'hc0083f09;
    11'b00000011111: data <= 32'hc1243cb9;
    11'b00000100000: data <= 32'hbadb314a;
    11'b00000100001: data <= 32'h3c58aee1;
    11'b00000100010: data <= 32'h3cd228ea;
    11'b00000100011: data <= 32'h3439b0af;
    11'b00000100100: data <= 32'h35a6b0fc;
    11'b00000100101: data <= 32'h3e323a8d;
    11'b00000100110: data <= 32'h3fb03f97;
    11'b00000100111: data <= 32'h39343d36;
    11'b00000101000: data <= 32'hba05baa4;
    11'b00000101001: data <= 32'hba80c066;
    11'b00000101010: data <= 32'hab90be01;
    11'b00000101011: data <= 32'h34c3b48e;
    11'b00000101100: data <= 32'h354cb814;
    11'b00000101101: data <= 32'h397cbe2f;
    11'b00000101110: data <= 32'h3a99bd0a;
    11'b00000101111: data <= 32'hb466386b;
    11'b00000110000: data <= 32'hbfef3f08;
    11'b00000110001: data <= 32'hc0bc3c22;
    11'b00000110010: data <= 32'hbc07b608;
    11'b00000110011: data <= 32'h31f7b9fb;
    11'b00000110100: data <= 32'hb256b277;
    11'b00000110101: data <= 32'hbb4831cc;
    11'b00000110110: data <= 32'hab7b36ad;
    11'b00000110111: data <= 32'h3f013cc6;
    11'b00000111000: data <= 32'h40444006;
    11'b00000111001: data <= 32'h37bd3e46;
    11'b00000111010: data <= 32'hbc631b98;
    11'b00000111011: data <= 32'hba99bb46;
    11'b00000111100: data <= 32'h37f5b690;
    11'b00000111101: data <= 32'h3c8c19e1;
    11'b00000111110: data <= 32'h3bc4bbf6;
    11'b00000111111: data <= 32'h3bb5c064;
    11'b00001000000: data <= 32'h3c3ebe1f;
    11'b00001000001: data <= 32'h357838d4;
    11'b00001000010: data <= 32'hbbe93e7f;
    11'b00001000011: data <= 32'hbe22360e;
    11'b00001000100: data <= 32'hbb88bd58;
    11'b00001000101: data <= 32'hb8aebdf4;
    11'b00001000110: data <= 32'hbcfab775;
    11'b00001000111: data <= 32'hbe523056;
    11'b00001001000: data <= 32'hb3a1308f;
    11'b00001001001: data <= 32'h3e6c38c0;
    11'b00001001010: data <= 32'h3e4c3e15;
    11'b00001001011: data <= 32'hb6673f06;
    11'b00001001100: data <= 32'hbf213bff;
    11'b00001001101: data <= 32'hbb913660;
    11'b00001001110: data <= 32'h3a0a3822;
    11'b00001001111: data <= 32'h3d2034af;
    11'b00001010000: data <= 32'h3a4abbce;
    11'b00001010001: data <= 32'h3a45bfac;
    11'b00001010010: data <= 32'h3dbebb59;
    11'b00001010011: data <= 32'h3dc83c65;
    11'b00001010100: data <= 32'h36733e34;
    11'b00001010101: data <= 32'hb866b21d;
    11'b00001010110: data <= 32'hb9a3bf91;
    11'b00001010111: data <= 32'hba7abeb1;
    11'b00001011000: data <= 32'hbd77b7db;
    11'b00001011001: data <= 32'hbd7ab45b;
    11'b00001011010: data <= 32'ha48dbb31;
    11'b00001011011: data <= 32'h3d69b9a7;
    11'b00001011100: data <= 32'h3a553946;
    11'b00001011101: data <= 32'hbcff3ee4;
    11'b00001011110: data <= 32'hc0743e38;
    11'b00001011111: data <= 32'hbc2a3b9d;
    11'b00001100000: data <= 32'h37e939c0;
    11'b00001100001: data <= 32'h37ec3579;
    11'b00001100010: data <= 32'hb43bb8ed;
    11'b00001100011: data <= 32'h30e5bc56;
    11'b00001100100: data <= 32'h3eb326a7;
    11'b00001100101: data <= 32'h40b43e8c;
    11'b00001100110: data <= 32'h3d613e5b;
    11'b00001100111: data <= 32'ha5e6b2d2;
    11'b00001101000: data <= 32'hb7dfbe0d;
    11'b00001101001: data <= 32'hb77cbbea;
    11'b00001101010: data <= 32'hb939affc;
    11'b00001101011: data <= 32'hb84fb9f5;
    11'b00001101100: data <= 32'h36e5c029;
    11'b00001101101: data <= 32'h3ce8bfbb;
    11'b00001101110: data <= 32'h36efaa53;
    11'b00001101111: data <= 32'hbd513e0f;
    11'b00001110000: data <= 32'hbfce3d96;
    11'b00001110001: data <= 32'hbb4b3819;
    11'b00001110010: data <= 32'had8c30ff;
    11'b00001110011: data <= 32'hba4b2f66;
    11'b00001110100: data <= 32'hbe70b430;
    11'b00001110101: data <= 32'hb8b1b69c;
    11'b00001110110: data <= 32'h3e8637fb;
    11'b00001110111: data <= 32'h41123ed2;
    11'b00001111000: data <= 32'h3d373e73;
    11'b00001111001: data <= 32'hb3e4352c;
    11'b00001111010: data <= 32'hb779b587;
    11'b00001111011: data <= 32'h2e293452;
    11'b00001111100: data <= 32'h33da3810;
    11'b00001111101: data <= 32'h31d4bba0;
    11'b00001111110: data <= 32'h397fc15e;
    11'b00001111111: data <= 32'h3d0fc0b3;
    11'b00010000000: data <= 32'h3a3eb148;
    11'b00010000001: data <= 32'hb7523d3f;
    11'b00010000010: data <= 32'hbbac39ee;
    11'b00010000011: data <= 32'hb7eab783;
    11'b00010000100: data <= 32'hb87ab925;
    11'b00010000101: data <= 32'hbf1bb0a4;
    11'b00010000110: data <= 32'hc0e4b0f4;
    11'b00010000111: data <= 32'hbbd7b737;
    11'b00010001000: data <= 32'h3d8225db;
    11'b00010001001: data <= 32'h3fe73c4b;
    11'b00010001010: data <= 32'h36e03dd2;
    11'b00010001011: data <= 32'hbbb23c09;
    11'b00010001100: data <= 32'hb8bf3b2e;
    11'b00010001101: data <= 32'h37743d89;
    11'b00010001110: data <= 32'h38bb3c3a;
    11'b00010001111: data <= 32'h2fc1ba49;
    11'b00010010000: data <= 32'h364fc0cf;
    11'b00010010001: data <= 32'h3d44bf1e;
    11'b00010010010: data <= 32'h3e4a3538;
    11'b00010010011: data <= 32'h3ae53cf7;
    11'b00010010100: data <= 32'h333e2de1;
    11'b00010010101: data <= 32'h296ebcc4;
    11'b00010010110: data <= 32'hb8c8bb97;
    11'b00010010111: data <= 32'hbf92ad96;
    11'b00010011000: data <= 32'hc09fb45e;
    11'b00010011001: data <= 32'hba6fbcc2;
    11'b00010011010: data <= 32'h3c77bcc8;
    11'b00010011011: data <= 32'h3c8c1db0;
    11'b00010011100: data <= 32'hb8713c5c;
    11'b00010011101: data <= 32'hbe163d5e;
    11'b00010011110: data <= 32'hb9143dc2;
    11'b00010011111: data <= 32'h37503ecd;
    11'b00010100000: data <= 32'h2de13ccd;
    11'b00010100001: data <= 32'hbab8b655;
    11'b00010100010: data <= 32'hb6fabe21;
    11'b00010100011: data <= 32'h3cd5b9d9;
    11'b00010100100: data <= 32'h40743bc4;
    11'b00010100101: data <= 32'h3f273d00;
    11'b00010100110: data <= 32'h3b39b09d;
    11'b00010100111: data <= 32'h3675bc53;
    11'b00010101000: data <= 32'hb242b5cf;
    11'b00010101001: data <= 32'hbc9d3767;
    11'b00010101010: data <= 32'hbda6b651;
    11'b00010101011: data <= 32'hb440c034;
    11'b00010101100: data <= 32'h3bd7c0cd;
    11'b00010101101: data <= 32'h38cdbb13;
    11'b00010101110: data <= 32'hbb123971;
    11'b00010101111: data <= 32'hbd6c3c59;
    11'b00010110000: data <= 32'hb5853be3;
    11'b00010110001: data <= 32'h32ef3c6e;
    11'b00010110010: data <= 32'hbb4d3b4a;
    11'b00010110011: data <= 32'hc051a96e;
    11'b00010110100: data <= 32'hbd86b9ba;
    11'b00010110101: data <= 32'h3b4ca787;
    11'b00010110110: data <= 32'h408e3ca3;
    11'b00010110111: data <= 32'h3ef43c91;
    11'b00010111000: data <= 32'h398d2c78;
    11'b00010111001: data <= 32'h367eb232;
    11'b00010111010: data <= 32'h35e73aec;
    11'b00010111011: data <= 32'hb0793d44;
    11'b00010111100: data <= 32'hb7c4b505;
    11'b00010111101: data <= 32'h2fbfc114;
    11'b00010111110: data <= 32'h3b5cc1a2;
    11'b00010111111: data <= 32'h3932bc3d;
    11'b00011000000: data <= 32'hb4aa3737;
    11'b00011000001: data <= 32'hb67636af;
    11'b00011000010: data <= 32'h34caad97;
    11'b00011000011: data <= 32'h2bb9302d;
    11'b00011000100: data <= 32'hbed93822;
    11'b00011000101: data <= 32'hc201302c;
    11'b00011000110: data <= 32'hbf85b7c2;
    11'b00011000111: data <= 32'h38a3b344;
    11'b00011001000: data <= 32'h3ebb38af;
    11'b00011001001: data <= 32'h3a583a1e;
    11'b00011001010: data <= 32'hb14f36c1;
    11'b00011001011: data <= 32'h30e83ab6;
    11'b00011001100: data <= 32'h3a3b3ff8;
    11'b00011001101: data <= 32'h371a4007;
    11'b00011001110: data <= 32'hb45ca314;
    11'b00011001111: data <= 32'hade6c066;
    11'b00011010000: data <= 32'h3a29c063;
    11'b00011010001: data <= 32'h3c69b766;
    11'b00011010010: data <= 32'h3a6737c9;
    11'b00011010011: data <= 32'h3a65b41b;
    11'b00011010100: data <= 32'h3c19bc13;
    11'b00011010101: data <= 32'h3299b70c;
    11'b00011010110: data <= 32'hbef83791;
    11'b00011010111: data <= 32'hc1ab31f8;
    11'b00011011000: data <= 32'hbe91bb1f;
    11'b00011011001: data <= 32'h3651bcd1;
    11'b00011011010: data <= 32'h3a97b7f6;
    11'b00011011011: data <= 32'hb60031d2;
    11'b00011011100: data <= 32'hbbd63832;
    11'b00011011101: data <= 32'ha0253d16;
    11'b00011011110: data <= 32'h3b4e4098;
    11'b00011011111: data <= 32'h3438404b;
    11'b00011100000: data <= 32'hbbda356d;
    11'b00011100001: data <= 32'hbb69bd38;
    11'b00011100010: data <= 32'h36d6bbe0;
    11'b00011100011: data <= 32'h3df636b9;
    11'b00011100100: data <= 32'h3e613906;
    11'b00011100101: data <= 32'h3df3b8da;
    11'b00011100110: data <= 32'h3db8bcd7;
    11'b00011100111: data <= 32'h38f3af70;
    11'b00011101000: data <= 32'hbbca3c08;
    11'b00011101001: data <= 32'hbf3234cc;
    11'b00011101010: data <= 32'hbb1abe09;
    11'b00011101011: data <= 32'h3654c084;
    11'b00011101100: data <= 32'h3258bdab;
    11'b00011101101: data <= 32'hbbe9b53f;
    11'b00011101110: data <= 32'hbc5432a0;
    11'b00011101111: data <= 32'h33d43a37;
    11'b00011110000: data <= 32'h3b2f3e65;
    11'b00011110001: data <= 32'hb6ed3eb3;
    11'b00011110010: data <= 32'hc043387e;
    11'b00011110011: data <= 32'hbfa6b6b5;
    11'b00011110100: data <= 32'ha407a346;
    11'b00011110101: data <= 32'h3db33b19;
    11'b00011110110: data <= 32'h3df538a9;
    11'b00011110111: data <= 32'h3cd0b8ce;
    11'b00011111000: data <= 32'h3d2eb918;
    11'b00011111001: data <= 32'h3c483b69;
    11'b00011111010: data <= 32'h2e1c3fa2;
    11'b00011111011: data <= 32'hb8fa3886;
    11'b00011111100: data <= 32'hb2f7bf25;
    11'b00011111101: data <= 32'h36cdc134;
    11'b00011111110: data <= 32'h2bc1be33;
    11'b00011111111: data <= 32'hb9b7b794;
    11'b00100000000: data <= 32'hb559b61b;
    11'b00100000001: data <= 32'h3b75b582;
    11'b00100000010: data <= 32'h3b9f364d;
    11'b00100000011: data <= 32'hbc213c00;
    11'b00100000100: data <= 32'hc1c738f7;
    11'b00100000101: data <= 32'hc0cca69d;
    11'b00100000110: data <= 32'hb5262ecd;
    11'b00100000111: data <= 32'h3af5384b;
    11'b00100001000: data <= 32'h37f53197;
    11'b00100001001: data <= 32'h308bb79a;
    11'b00100001010: data <= 32'h3a36314c;
    11'b00100001011: data <= 32'h3d693fd5;
    11'b00100001100: data <= 32'h3a8a4140;
    11'b00100001101: data <= 32'hadff3b2b;
    11'b00100001110: data <= 32'hb1dfbdc4;
    11'b00100001111: data <= 32'h3446bfb8;
    11'b00100010000: data <= 32'h3483ba3f;
    11'b00100010001: data <= 32'h2fd5b25b;
    11'b00100010010: data <= 32'h3a17bb68;
    11'b00100010011: data <= 32'h3ecebd93;
    11'b00100010100: data <= 32'h3cbbb7c9;
    11'b00100010101: data <= 32'hbc11397f;
    11'b00100010110: data <= 32'hc157393e;
    11'b00100010111: data <= 32'hc00db291;
    11'b00100011000: data <= 32'hb4dfb8c2;
    11'b00100011001: data <= 32'h3030b6bc;
    11'b00100011010: data <= 32'hba34b785;
    11'b00100011011: data <= 32'hbbc6b809;
    11'b00100011100: data <= 32'h35453817;
    11'b00100011101: data <= 32'h3dbd406d;
    11'b00100011110: data <= 32'h3acc4152;
    11'b00100011111: data <= 32'hb8133c5f;
    11'b00100100000: data <= 32'hbaf4b92c;
    11'b00100100001: data <= 32'hb08db900;
    11'b00100100010: data <= 32'h3800363b;
    11'b00100100011: data <= 32'h3a553391;
    11'b00100100100: data <= 32'h3d98bccb;
    11'b00100100101: data <= 32'h401cbf21;
    11'b00100100110: data <= 32'h3df8b77e;
    11'b00100100111: data <= 32'hb5283c2f;
    11'b00100101000: data <= 32'hbe323a9f;
    11'b00100101001: data <= 32'hbc02b907;
    11'b00100101010: data <= 32'ha1d4bdf3;
    11'b00100101011: data <= 32'hb665bd26;
    11'b00100101100: data <= 32'hbe4abbc2;
    11'b00100101101: data <= 32'hbd91ba38;
    11'b00100101110: data <= 32'h36092ba1;
    11'b00100101111: data <= 32'h3dd83dc0;
    11'b00100110000: data <= 32'h35cd3fca;
    11'b00100110001: data <= 32'hbddf3c23;
    11'b00100110010: data <= 32'hbf2e3046;
    11'b00100110011: data <= 32'hb8e33822;
    11'b00100110100: data <= 32'h36be3cbc;
    11'b00100110101: data <= 32'h398f36d0;
    11'b00100110110: data <= 32'h3c34bcd8;
    11'b00100110111: data <= 32'h3edebdb2;
    11'b00100111000: data <= 32'h3ec335ba;
    11'b00100111001: data <= 32'h391e3f7e;
    11'b00100111010: data <= 32'hb2bf3c94;
    11'b00100111011: data <= 32'h19e8babc;
    11'b00100111100: data <= 32'h347fbf39;
    11'b00100111101: data <= 32'hb83fbd79;
    11'b00100111110: data <= 32'hbe10bbab;
    11'b00100111111: data <= 32'hbb16bc9b;
    11'b00101000000: data <= 32'h3bc7bbb1;
    11'b00101000001: data <= 32'h3e532d6a;
    11'b00101000010: data <= 32'hb03a3b82;
    11'b00101000011: data <= 32'hc0573a78;
    11'b00101000100: data <= 32'hc07b37ed;
    11'b00101000101: data <= 32'hba783ad8;
    11'b00101000110: data <= 32'h281c3c69;
    11'b00101000111: data <= 32'hb2cd305b;
    11'b00101001000: data <= 32'hb09dbc9e;
    11'b00101001001: data <= 32'h3b02ba13;
    11'b00101001010: data <= 32'h3eb33d37;
    11'b00101001011: data <= 32'h3d3b411c;
    11'b00101001100: data <= 32'h38463da6;
    11'b00101001101: data <= 32'h355cb8e3;
    11'b00101001110: data <= 32'h3465bcca;
    11'b00101001111: data <= 32'hb5f8b7b2;
    11'b00101010000: data <= 32'hbabdb629;
    11'b00101010001: data <= 32'h2e24bd9b;
    11'b00101010010: data <= 32'h3edabfc5;
    11'b00101010011: data <= 32'h3f2bbc09;
    11'b00101010100: data <= 32'hb1bc34d3;
    11'b00101010101: data <= 32'hbff9393b;
    11'b00101010110: data <= 32'hbf1035d7;
    11'b00101010111: data <= 32'hb836356f;
    11'b00101011000: data <= 32'hb6dc34a3;
    11'b00101011001: data <= 32'hbda4b7a5;
    11'b00101011010: data <= 32'hbdddbcce;
    11'b00101011011: data <= 32'h2d82b65d;
    11'b00101011100: data <= 32'h3e203e53;
    11'b00101011101: data <= 32'h3d7a4106;
    11'b00101011110: data <= 32'h351f3d8a;
    11'b00101011111: data <= 32'hb177ac4a;
    11'b00101100000: data <= 32'hadc42835;
    11'b00101100001: data <= 32'hb25f3b1f;
    11'b00101100010: data <= 32'hb2753673;
    11'b00101100011: data <= 32'h39e6bdad;
    11'b00101100100: data <= 32'h4006c0ad;
    11'b00101100101: data <= 32'h3fb3bcd1;
    11'b00101100110: data <= 32'h34c8371a;
    11'b00101100111: data <= 32'hbb863a0d;
    11'b00101101000: data <= 32'hb86a10b7;
    11'b00101101001: data <= 32'h2fbdb7c4;
    11'b00101101010: data <= 32'hb97cb877;
    11'b00101101011: data <= 32'hc066bb91;
    11'b00101101100: data <= 32'hc038bd66;
    11'b00101101101: data <= 32'hafbab963;
    11'b00101101110: data <= 32'h3dd23af6;
    11'b00101101111: data <= 32'h3b8c3e82;
    11'b00101110000: data <= 32'hb84c3be0;
    11'b00101110001: data <= 32'hbc3536e7;
    11'b00101110010: data <= 32'hb8573c9f;
    11'b00101110011: data <= 32'hb27a3fae;
    11'b00101110100: data <= 32'hb14e3b11;
    11'b00101110101: data <= 32'h372abd2c;
    11'b00101110110: data <= 32'h3e1ac013;
    11'b00101110111: data <= 32'h3f37b811;
    11'b00101111000: data <= 32'h3bd93cc8;
    11'b00101111001: data <= 32'h35eb3c3e;
    11'b00101111010: data <= 32'h3995b3e0;
    11'b00101111011: data <= 32'h39e6bb24;
    11'b00101111100: data <= 32'hb925b984;
    11'b00101111101: data <= 32'hc061ba8b;
    11'b00101111110: data <= 32'hbf0bbdc3;
    11'b00101111111: data <= 32'h35d7bdb6;
    11'b00110000000: data <= 32'h3e3ab731;
    11'b00110000001: data <= 32'h372535ed;
    11'b00110000010: data <= 32'hbd263686;
    11'b00110000011: data <= 32'hbe2738b1;
    11'b00110000100: data <= 32'hb93d3e23;
    11'b00110000101: data <= 32'hb5ab400c;
    11'b00110000110: data <= 32'hbaa239f0;
    11'b00110000111: data <= 32'hb9acbcd0;
    11'b00110001000: data <= 32'h371fbd91;
    11'b00110001001: data <= 32'h3db13733;
    11'b00110001010: data <= 32'h3da93fa2;
    11'b00110001011: data <= 32'h3c973d18;
    11'b00110001100: data <= 32'h3cf8b28d;
    11'b00110001101: data <= 32'h3b65b7fa;
    11'b00110001110: data <= 32'hb6d930f4;
    11'b00110001111: data <= 32'hbe36a558;
    11'b00110010000: data <= 32'hba68bd4d;
    11'b00110010001: data <= 32'h3c7bc050;
    11'b00110010010: data <= 32'h3ef1be46;
    11'b00110010011: data <= 32'h3418b80b;
    11'b00110010100: data <= 32'hbd2c21b5;
    11'b00110010101: data <= 32'hbc7035e2;
    11'b00110010110: data <= 32'hb1913c41;
    11'b00110010111: data <= 32'hb7723d12;
    11'b00110011000: data <= 32'hbf143056;
    11'b00110011001: data <= 32'hc019bcf0;
    11'b00110011010: data <= 32'hb8d4bb6d;
    11'b00110011011: data <= 32'h3bf23b0b;
    11'b00110011100: data <= 32'h3d693faa;
    11'b00110011101: data <= 32'h3be13c4f;
    11'b00110011110: data <= 32'h3aab23fa;
    11'b00110011111: data <= 32'h38ca37a7;
    11'b00110100000: data <= 32'hb3da3e28;
    11'b00110100001: data <= 32'hbac63c27;
    11'b00110100010: data <= 32'ha8a2bc16;
    11'b00110100011: data <= 32'h3de8c0ca;
    11'b00110100100: data <= 32'h3ef1bf44;
    11'b00110100101: data <= 32'h3719b7fe;
    11'b00110100110: data <= 32'hb7c02825;
    11'b00110100111: data <= 32'h2f1ba1b5;
    11'b00110101000: data <= 32'h39fa3290;
    11'b00110101001: data <= 32'hb6073540;
    11'b00110101010: data <= 32'hc0bfb64a;
    11'b00110101011: data <= 32'hc17fbd25;
    11'b00110101100: data <= 32'hbbe3bb9d;
    11'b00110101101: data <= 32'h3a4c3667;
    11'b00110101110: data <= 32'h3b293c21;
    11'b00110101111: data <= 32'h2f86368d;
    11'b00110110000: data <= 32'haeb43101;
    11'b00110110001: data <= 32'h2dcf3d98;
    11'b00110110010: data <= 32'hb1ee4141;
    11'b00110110011: data <= 32'hb8cc3eec;
    11'b00110110100: data <= 32'haf04b9bb;
    11'b00110110101: data <= 32'h3c07c013;
    11'b00110110110: data <= 32'h3d75bc85;
    11'b00110110111: data <= 32'h3a243456;
    11'b00110111000: data <= 32'h38e63609;
    11'b00110111001: data <= 32'h3db0b4be;
    11'b00110111010: data <= 32'h3e71b5f5;
    11'b00110111011: data <= 32'haeda98bb;
    11'b00110111100: data <= 32'hc091b4cd;
    11'b00110111101: data <= 32'hc0d9bca1;
    11'b00110111110: data <= 32'hb82dbd6f;
    11'b00110111111: data <= 32'h3b39b996;
    11'b00111000000: data <= 32'h35f6b494;
    11'b00111000001: data <= 32'hba22b711;
    11'b00111000010: data <= 32'hba29294e;
    11'b00111000011: data <= 32'hacbc3eb0;
    11'b00111000100: data <= 32'hb0f1418b;
    11'b00111000101: data <= 32'hbb823ea0;
    11'b00111000110: data <= 32'hbc2ab8d8;
    11'b00111000111: data <= 32'hb01cbd7b;
    11'b00111001000: data <= 32'h398bac54;
    11'b00111001001: data <= 32'h3b2c3c8f;
    11'b00111001010: data <= 32'h3d0d393b;
    11'b00111001011: data <= 32'h400eb668;
    11'b00111001100: data <= 32'h3fa7b462;
    11'b00111001101: data <= 32'h317a38f1;
    11'b00111001110: data <= 32'hbe78384e;
    11'b00111001111: data <= 32'hbd8db9ff;
    11'b00111010000: data <= 32'h35d2bf08;
    11'b00111010001: data <= 32'h3c9abeae;
    11'b00111010010: data <= 32'h2c7dbcf5;
    11'b00111010011: data <= 32'hbc26bc05;
    11'b00111010100: data <= 32'hb881b4a0;
    11'b00111010101: data <= 32'h36df3ca7;
    11'b00111010110: data <= 32'h23cd3fe0;
    11'b00111010111: data <= 32'hbe263b9c;
    11'b00111011000: data <= 32'hc06fb9a1;
    11'b00111011001: data <= 32'hbd11ba92;
    11'b00111011010: data <= 32'h2a3a38c8;
    11'b00111011011: data <= 32'h395f3d76;
    11'b00111011100: data <= 32'h3c2f3754;
    11'b00111011101: data <= 32'h3e65b705;
    11'b00111011110: data <= 32'h3e1f35ce;
    11'b00111011111: data <= 32'h34d03f4f;
    11'b00111100000: data <= 32'hbac83ec5;
    11'b00111100001: data <= 32'hb6a4b22d;
    11'b00111100010: data <= 32'h3b78bf26;
    11'b00111100011: data <= 32'h3cb2bf65;
    11'b00111100100: data <= 32'h26f2bcfb;
    11'b00111100101: data <= 32'hb87abbd0;
    11'b00111100110: data <= 32'h3799b921;
    11'b00111100111: data <= 32'h3dc8340f;
    11'b00111101000: data <= 32'h361e3acb;
    11'b00111101001: data <= 32'hbf9332ed;
    11'b00111101010: data <= 32'hc1aaba69;
    11'b00111101011: data <= 32'hbec3b92a;
    11'b00111101100: data <= 32'hb29336fe;
    11'b00111101101: data <= 32'h327e3964;
    11'b00111101110: data <= 32'h3051b4c0;
    11'b00111101111: data <= 32'h381ab8b8;
    11'b00111110000: data <= 32'h3aa73c06;
    11'b00111110001: data <= 32'h34be41a3;
    11'b00111110010: data <= 32'hb6ef40e8;
    11'b00111110011: data <= 32'hb1e332ea;
    11'b00111110100: data <= 32'h3959bd7f;
    11'b00111110101: data <= 32'h39dfbc77;
    11'b00111110110: data <= 32'h2b4eb5bf;
    11'b00111110111: data <= 32'h33afb77c;
    11'b00111111000: data <= 32'h3eb7bad6;
    11'b00111111001: data <= 32'h40cdb760;
    11'b00111111010: data <= 32'h3a783369;
    11'b00111111011: data <= 32'hbed02dec;
    11'b00111111100: data <= 32'hc0ebb908;
    11'b00111111101: data <= 32'hbc95ba23;
    11'b00111111110: data <= 32'h28c0b5a0;
    11'b00111111111: data <= 32'hb40eb838;
    11'b01000000000: data <= 32'hbae7bd0b;
    11'b01000000001: data <= 32'hb6b6bb46;
    11'b01000000010: data <= 32'h370a3c8d;
    11'b01000000011: data <= 32'h357441d2;
    11'b01000000100: data <= 32'hb80c40ac;
    11'b01000000101: data <= 32'hba6333dd;
    11'b01000000110: data <= 32'hb560ba09;
    11'b01000000111: data <= 32'habce2979;
    11'b01000001000: data <= 32'hab553a09;
    11'b01000001001: data <= 32'h39b028fa;
    11'b01000001010: data <= 32'h4076bb8c;
    11'b01000001011: data <= 32'h4167b8d4;
    11'b01000001100: data <= 32'h3c3b3841;
    11'b01000001101: data <= 32'hbc3d3a3f;
    11'b01000001110: data <= 32'hbd58ae6a;
    11'b01000001111: data <= 32'ha8fbbb2b;
    11'b01000010000: data <= 32'h3814bc70;
    11'b01000010001: data <= 32'hb827bdb3;
    11'b01000010010: data <= 32'hbd65bf75;
    11'b01000010011: data <= 32'hb83dbd12;
    11'b01000010100: data <= 32'h3a2f38f5;
    11'b01000010101: data <= 32'h38ee400f;
    11'b01000010110: data <= 32'hba923dc2;
    11'b01000010111: data <= 32'hbef0ac00;
    11'b01000011000: data <= 32'hbda8b419;
    11'b01000011001: data <= 32'hba453b36;
    11'b01000011010: data <= 32'hb5ec3d2d;
    11'b01000011011: data <= 32'h3736285f;
    11'b01000011100: data <= 32'h3ef2bc42;
    11'b01000011101: data <= 32'h4054b406;
    11'b01000011110: data <= 32'h3c033dec;
    11'b01000011111: data <= 32'hb5823f78;
    11'b01000100000: data <= 32'hb2113884;
    11'b01000100001: data <= 32'h3ab8ba42;
    11'b01000100010: data <= 32'h39f4bcd5;
    11'b01000100011: data <= 32'hb8f3bd81;
    11'b01000100100: data <= 32'hbc98bee8;
    11'b01000100101: data <= 32'h3366bde4;
    11'b01000100110: data <= 32'h3ed5b3a7;
    11'b01000100111: data <= 32'h3c703a09;
    11'b01000101000: data <= 32'hbbeb3673;
    11'b01000101001: data <= 32'hc077b637;
    11'b01000101010: data <= 32'hbf2caa6d;
    11'b01000101011: data <= 32'hbbd43c08;
    11'b01000101100: data <= 32'hb9ed3b26;
    11'b01000101101: data <= 32'hb6c9b8fb;
    11'b01000101110: data <= 32'h3818bd65;
    11'b01000101111: data <= 32'h3cb83178;
    11'b01000110000: data <= 32'h3a1440a6;
    11'b01000110001: data <= 32'h2cca412f;
    11'b01000110010: data <= 32'h34c33bb7;
    11'b01000110011: data <= 32'h3b0cb696;
    11'b01000110100: data <= 32'h36ceb7db;
    11'b01000110101: data <= 32'hb9c0b5eb;
    11'b01000110110: data <= 32'hb8bfbbab;
    11'b01000110111: data <= 32'h3d0fbdcd;
    11'b01000111000: data <= 32'h4144bb82;
    11'b01000111001: data <= 32'h3e4aaeca;
    11'b01000111010: data <= 32'hba47a942;
    11'b01000111011: data <= 32'hbf65b5db;
    11'b01000111100: data <= 32'hbc96ab11;
    11'b01000111101: data <= 32'hb81a37ac;
    11'b01000111110: data <= 32'hbbd2af41;
    11'b01000111111: data <= 32'hbd94be3d;
    11'b01001000000: data <= 32'hb931befa;
    11'b01001000001: data <= 32'h3755338e;
    11'b01001000010: data <= 32'h38fd40c3;
    11'b01001000011: data <= 32'h2e4840c8;
    11'b01001000100: data <= 32'haa013a84;
    11'b01001000101: data <= 32'h2e2024bb;
    11'b01001000110: data <= 32'hb565391d;
    11'b01001000111: data <= 32'hbb863ba8;
    11'b01001001000: data <= 32'hb38baf97;
    11'b01001001001: data <= 32'h3f08bd53;
    11'b01001001010: data <= 32'h41bfbc9b;
    11'b01001001011: data <= 32'h3ec4ad11;
    11'b01001001100: data <= 32'hb4ad366a;
    11'b01001001101: data <= 32'hb9fe2f4c;
    11'b01001001110: data <= 32'h3110ab3a;
    11'b01001001111: data <= 32'h3498affb;
    11'b01001010000: data <= 32'hbc12bb74;
    11'b01001010001: data <= 32'hbfb6c040;
    11'b01001010010: data <= 32'hbc21c00d;
    11'b01001010011: data <= 32'h3824b19f;
    11'b01001010100: data <= 32'h3a993e10;
    11'b01001010101: data <= 32'had543d42;
    11'b01001010110: data <= 32'hba5c3234;
    11'b01001010111: data <= 32'hbb0b348d;
    11'b01001011000: data <= 32'hbc2b3e1c;
    11'b01001011001: data <= 32'hbcec3f13;
    11'b01001011010: data <= 32'hb701319f;
    11'b01001011011: data <= 32'h3d12bd63;
    11'b01001011100: data <= 32'h405cbb6d;
    11'b01001011101: data <= 32'h3d66393e;
    11'b01001011110: data <= 32'h323c3d6f;
    11'b01001011111: data <= 32'h36a93a2f;
    11'b01001100000: data <= 32'h3d3b2d61;
    11'b01001100001: data <= 32'h3abfb36e;
    11'b01001100010: data <= 32'hbbd8bb03;
    11'b01001100011: data <= 32'hbf61bf72;
    11'b01001100100: data <= 32'hb80abfee;
    11'b01001100101: data <= 32'h3d30ba92;
    11'b01001100110: data <= 32'h3d40334c;
    11'b01001100111: data <= 32'hb1ef219d;
    11'b01001101000: data <= 32'hbd06b78d;
    11'b01001101001: data <= 32'hbcf6352e;
    11'b01001101010: data <= 32'hbc943ef3;
    11'b01001101011: data <= 32'hbd9c3e79;
    11'b01001101100: data <= 32'hbc80b4ba;
    11'b01001101101: data <= 32'h288cbe77;
    11'b01001101110: data <= 32'h3b81b8cb;
    11'b01001101111: data <= 32'h3a0e3daf;
    11'b01001110000: data <= 32'h36c0401a;
    11'b01001110001: data <= 32'h3bf33c73;
    11'b01001110010: data <= 32'h3e7634f7;
    11'b01001110011: data <= 32'h39f23555;
    11'b01001110100: data <= 32'hbc313050;
    11'b01001110101: data <= 32'hbd98bad4;
    11'b01001110110: data <= 32'h36a2be73;
    11'b01001110111: data <= 32'h405abd3e;
    11'b01001111000: data <= 32'h3ef9b9af;
    11'b01001111001: data <= 32'hac88b9bc;
    11'b01001111010: data <= 32'hbbdeb9a5;
    11'b01001111011: data <= 32'hb8b7342d;
    11'b01001111100: data <= 32'hb7763d4f;
    11'b01001111101: data <= 32'hbd3c3a0c;
    11'b01001111110: data <= 32'hbf84bcac;
    11'b01001111111: data <= 32'hbcc4c000;
    11'b01010000000: data <= 32'had22b7e4;
    11'b01010000001: data <= 32'h353b3e34;
    11'b01010000010: data <= 32'h35b43f63;
    11'b01010000011: data <= 32'h3a2b3a42;
    11'b01010000100: data <= 32'h3c063712;
    11'b01010000101: data <= 32'h2c643d03;
    11'b01010000110: data <= 32'hbd163e14;
    11'b01010000111: data <= 32'hbc2c349c;
    11'b01010001000: data <= 32'h3b8dbcac;
    11'b01010001001: data <= 32'h40d3bd9c;
    11'b01010001010: data <= 32'h3ee0ba6e;
    11'b01010001011: data <= 32'h313db7b9;
    11'b01010001100: data <= 32'had07b586;
    11'b01010001101: data <= 32'h3a22343d;
    11'b01010001110: data <= 32'h39123a18;
    11'b01010001111: data <= 32'hbc04ac17;
    11'b01010010000: data <= 32'hc086beed;
    11'b01010010001: data <= 32'hbec4c05b;
    11'b01010010010: data <= 32'hb429b98a;
    11'b01010010011: data <= 32'h35e73adb;
    11'b01010010100: data <= 32'h317339cb;
    11'b01010010101: data <= 32'h2dbfb018;
    11'b01010010110: data <= 32'h2c1035ae;
    11'b01010010111: data <= 32'hb9103fe3;
    11'b01010011000: data <= 32'hbdfc40e2;
    11'b01010011001: data <= 32'hbc543acc;
    11'b01010011010: data <= 32'h38d4bbdb;
    11'b01010011011: data <= 32'h3ebbbc9d;
    11'b01010011100: data <= 32'h3c6db103;
    11'b01010011101: data <= 32'h34d8367e;
    11'b01010011110: data <= 32'h3b4134cc;
    11'b01010011111: data <= 32'h400d35f4;
    11'b01010100000: data <= 32'h3dee3852;
    11'b01010100001: data <= 32'hb9c6b043;
    11'b01010100010: data <= 32'hc041bdc8;
    11'b01010100011: data <= 32'hbd0ebf94;
    11'b01010100100: data <= 32'h369abc07;
    11'b01010100101: data <= 32'h3a96b3ea;
    11'b01010100110: data <= 32'h2b4bb97f;
    11'b01010100111: data <= 32'hb708bc6d;
    11'b01010101000: data <= 32'hb6502f21;
    11'b01010101001: data <= 32'hb9d34035;
    11'b01010101010: data <= 32'hbdde40ce;
    11'b01010101011: data <= 32'hbddd382f;
    11'b01010101100: data <= 32'hb72abcc1;
    11'b01010101101: data <= 32'h3565ba95;
    11'b01010101110: data <= 32'h31ff391c;
    11'b01010101111: data <= 32'h32e73cac;
    11'b01010110000: data <= 32'h3d8a3929;
    11'b01010110001: data <= 32'h40e93711;
    11'b01010110010: data <= 32'h3e443ab7;
    11'b01010110011: data <= 32'hb98639a1;
    11'b01010110100: data <= 32'hbeb8b588;
    11'b01010110101: data <= 32'hb58cbcc9;
    11'b01010110110: data <= 32'h3d54bca4;
    11'b01010110111: data <= 32'h3d11bc44;
    11'b01010111000: data <= 32'h2b49be31;
    11'b01010111001: data <= 32'hb640be45;
    11'b01010111010: data <= 32'h2e00add4;
    11'b01010111011: data <= 32'h269e3ebd;
    11'b01010111100: data <= 32'hbc3d3e48;
    11'b01010111101: data <= 32'hbf80b5bb;
    11'b01010111110: data <= 32'hbe2abe58;
    11'b01010111111: data <= 32'hba96b91b;
    11'b01011000000: data <= 32'hb8153b9a;
    11'b01011000001: data <= 32'ha86e3c73;
    11'b01011000010: data <= 32'h3c8d3426;
    11'b01011000011: data <= 32'h3f9b3490;
    11'b01011000100: data <= 32'h3b593dae;
    11'b01011000101: data <= 32'hbb5b3fc7;
    11'b01011000110: data <= 32'hbd183b8c;
    11'b01011000111: data <= 32'h3539b732;
    11'b01011001000: data <= 32'h3ed1bc17;
    11'b01011001001: data <= 32'h3cd4bc7b;
    11'b01011001010: data <= 32'h28dbbd95;
    11'b01011001011: data <= 32'h3229bd1b;
    11'b01011001100: data <= 32'h3d35ae7b;
    11'b01011001101: data <= 32'h3d163c5a;
    11'b01011001110: data <= 32'hb6d73922;
    11'b01011001111: data <= 32'hbff5bc2e;
    11'b01011010000: data <= 32'hbfeebf01;
    11'b01011010001: data <= 32'hbc71b8fa;
    11'b01011010010: data <= 32'hb8b3386f;
    11'b01011010011: data <= 32'hb43f3070;
    11'b01011010100: data <= 32'h3703ba50;
    11'b01011010101: data <= 32'h3b13b072;
    11'b01011010110: data <= 32'h2f273f5f;
    11'b01011010111: data <= 32'hbc9b4197;
    11'b01011011000: data <= 32'hbc8b3e8a;
    11'b01011011001: data <= 32'h341cadec;
    11'b01011011010: data <= 32'h3c7eb983;
    11'b01011011011: data <= 32'h3789b750;
    11'b01011011100: data <= 32'hb114b77c;
    11'b01011011101: data <= 32'h3aeeb868;
    11'b01011011110: data <= 32'h40f426d7;
    11'b01011011111: data <= 32'h408a39d5;
    11'b01011100000: data <= 32'h2cc73547;
    11'b01011100001: data <= 32'hbee8bb49;
    11'b01011100010: data <= 32'hbe24bd75;
    11'b01011100011: data <= 32'hb6edb8e8;
    11'b01011100100: data <= 32'had92b36f;
    11'b01011100101: data <= 32'hb5b3bcba;
    11'b01011100110: data <= 32'hb233bfbe;
    11'b01011100111: data <= 32'h32d8b92b;
    11'b01011101000: data <= 32'hb0743f39;
    11'b01011101001: data <= 32'hbc304175;
    11'b01011101010: data <= 32'hbce23d59;
    11'b01011101011: data <= 32'hb7a5b4d8;
    11'b01011101100: data <= 32'hafddb5e6;
    11'b01011101101: data <= 32'hb90336a4;
    11'b01011101110: data <= 32'hb85c379b;
    11'b01011101111: data <= 32'h3c8caa82;
    11'b01011110000: data <= 32'h41c02acb;
    11'b01011110001: data <= 32'h40d73a18;
    11'b01011110010: data <= 32'h30d53adc;
    11'b01011110011: data <= 32'hbd102d23;
    11'b01011110100: data <= 32'hb878b7cb;
    11'b01011110101: data <= 32'h3916b712;
    11'b01011110110: data <= 32'h3805ba82;
    11'b01011110111: data <= 32'hb5f5c004;
    11'b01011111000: data <= 32'hb5ffc0ff;
    11'b01011111001: data <= 32'h3681bb93;
    11'b01011111010: data <= 32'h37e53d5f;
    11'b01011111011: data <= 32'hb7903f63;
    11'b01011111100: data <= 32'hbd2b356c;
    11'b01011111101: data <= 32'hbd3cbaa5;
    11'b01011111110: data <= 32'hbcfcb1f9;
    11'b01011111111: data <= 32'hbdda3b5f;
    11'b01100000000: data <= 32'hbb983996;
    11'b01100000001: data <= 32'h3a84b4d4;
    11'b01100000010: data <= 32'h4090b3f7;
    11'b01100000011: data <= 32'h3ec23c07;
    11'b01100000100: data <= 32'hb1e73f47;
    11'b01100000101: data <= 32'hbafa3d4f;
    11'b01100000110: data <= 32'h347a36df;
    11'b01100000111: data <= 32'h3d14ae2d;
    11'b01100001000: data <= 32'h38bbba0b;
    11'b01100001001: data <= 32'hb812bf4e;
    11'b01100001010: data <= 32'haf2fc055;
    11'b01100001011: data <= 32'h3d4ebb13;
    11'b01100001100: data <= 32'h3ec13a11;
    11'b01100001101: data <= 32'h35963a3a;
    11'b01100001110: data <= 32'hbc9db8b9;
    11'b01100001111: data <= 32'hbe69bc9d;
    11'b01100010000: data <= 32'hbe0dad53;
    11'b01100010001: data <= 32'hbe303a9a;
    11'b01100010010: data <= 32'hbc9c2410;
    11'b01100010011: data <= 32'h2f80bd27;
    11'b01100010100: data <= 32'h3c96baf7;
    11'b01100010101: data <= 32'h39483c91;
    11'b01100010110: data <= 32'hb8a640fb;
    11'b01100010111: data <= 32'hb9694002;
    11'b01100011000: data <= 32'h37c93abd;
    11'b01100011001: data <= 32'h3bd83439;
    11'b01100011010: data <= 32'hac62ace1;
    11'b01100011011: data <= 32'hbb34ba69;
    11'b01100011100: data <= 32'h340abcfc;
    11'b01100011101: data <= 32'h4098b8be;
    11'b01100011110: data <= 32'h415b35de;
    11'b01100011111: data <= 32'h3ba032da;
    11'b01100100000: data <= 32'hba73b9ff;
    11'b01100100001: data <= 32'hbc74bae9;
    11'b01100100010: data <= 32'hba112eea;
    11'b01100100011: data <= 32'hbb1d35b8;
    11'b01100100100: data <= 32'hbc60bc54;
    11'b01100100101: data <= 32'hb83bc0dc;
    11'b01100100110: data <= 32'h33f5be14;
    11'b01100100111: data <= 32'h2f7d3bb9;
    11'b01100101000: data <= 32'hb8c840b5;
    11'b01100101001: data <= 32'hb8cc3e99;
    11'b01100101010: data <= 32'h2ca83827;
    11'b01100101011: data <= 32'ha7643765;
    11'b01100101100: data <= 32'hbca53a69;
    11'b01100101101: data <= 32'hbdd83585;
    11'b01100101110: data <= 32'h3561b75a;
    11'b01100101111: data <= 32'h4133b6c1;
    11'b01100110000: data <= 32'h41943442;
    11'b01100110001: data <= 32'h3bba36d2;
    11'b01100110010: data <= 32'hb6daa1c9;
    11'b01100110011: data <= 32'hb0201563;
    11'b01100110100: data <= 32'h37db379f;
    11'b01100110101: data <= 32'ha62c1a66;
    11'b01100110110: data <= 32'hbb96bf2a;
    11'b01100110111: data <= 32'hba81c1f3;
    11'b01100111000: data <= 32'h305dbf3d;
    11'b01100111001: data <= 32'h37b13851;
    11'b01100111010: data <= 32'haab43dd2;
    11'b01100111011: data <= 32'hb77037e0;
    11'b01100111100: data <= 32'hb7fab437;
    11'b01100111101: data <= 32'hbc0f379a;
    11'b01100111110: data <= 32'hc0003d8a;
    11'b01100111111: data <= 32'hbfa23adf;
    11'b01101000000: data <= 32'h13f7b6d4;
    11'b01101000001: data <= 32'h3fe9b95c;
    11'b01101000010: data <= 32'h3fb234f3;
    11'b01101000011: data <= 32'h36763c6b;
    11'b01101000100: data <= 32'hb25c3c4f;
    11'b01101000101: data <= 32'h3a243b7e;
    11'b01101000110: data <= 32'h3d9a3b56;
    11'b01101000111: data <= 32'h35c13006;
    11'b01101001000: data <= 32'hbc01be44;
    11'b01101001001: data <= 32'hb9e8c112;
    11'b01101001010: data <= 32'h3a15be3c;
    11'b01101001011: data <= 32'h3dfc2eb2;
    11'b01101001100: data <= 32'h3a5d356f;
    11'b01101001101: data <= 32'hb1f8b99a;
    11'b01101001110: data <= 32'hb96ebb1f;
    11'b01101001111: data <= 32'hbce5377f;
    11'b01101010000: data <= 32'hc0053dd3;
    11'b01101010001: data <= 32'hbfe337aa;
    11'b01101010010: data <= 32'hb895bcd9;
    11'b01101010011: data <= 32'h3a6bbd42;
    11'b01101010100: data <= 32'h392e345e;
    11'b01101010101: data <= 32'hb4c93e79;
    11'b01101010110: data <= 32'hb05e3ebd;
    11'b01101010111: data <= 32'h3c7c3d3d;
    11'b01101011000: data <= 32'h3dac3cc6;
    11'b01101011001: data <= 32'hace739bc;
    11'b01101011010: data <= 32'hbd9db809;
    11'b01101011011: data <= 32'hb880bd8e;
    11'b01101011100: data <= 32'h3e27bbbb;
    11'b01101011101: data <= 32'h40cdb059;
    11'b01101011110: data <= 32'h3d8fb5a1;
    11'b01101011111: data <= 32'h305fbcac;
    11'b01101100000: data <= 32'hb386bac8;
    11'b01101100001: data <= 32'hb6ed3932;
    11'b01101100010: data <= 32'hbc9d3cbd;
    11'b01101100011: data <= 32'hbe86b65d;
    11'b01101100100: data <= 32'hbc3dc082;
    11'b01101100101: data <= 32'hb298bfea;
    11'b01101100110: data <= 32'hb2a22c2b;
    11'b01101100111: data <= 32'hb8b83ded;
    11'b01101101000: data <= 32'hae253d28;
    11'b01101101001: data <= 32'h3b393a93;
    11'b01101101010: data <= 32'h393a3c92;
    11'b01101101011: data <= 32'hbc363dc1;
    11'b01101101100: data <= 32'hbffd39e5;
    11'b01101101101: data <= 32'hb877b4af;
    11'b01101101110: data <= 32'h3f30b7f5;
    11'b01101101111: data <= 32'h40f0b172;
    11'b01101110000: data <= 32'h3d1ab545;
    11'b01101110001: data <= 32'h34f5b992;
    11'b01101110010: data <= 32'h38e3afc5;
    11'b01101110011: data <= 32'h3b343c3d;
    11'b01101110100: data <= 32'h21f53b97;
    11'b01101110101: data <= 32'hbcaebc1a;
    11'b01101110110: data <= 32'hbcfdc182;
    11'b01101110111: data <= 32'hb7f5c05d;
    11'b01101111000: data <= 32'hb02db2a0;
    11'b01101111001: data <= 32'hb2c63990;
    11'b01101111010: data <= 32'h2d002b20;
    11'b01101111011: data <= 32'h37b3b3dd;
    11'b01101111100: data <= 32'hb2ee3ab1;
    11'b01101111101: data <= 32'hbf633f9d;
    11'b01101111110: data <= 32'hc0cb3dab;
    11'b01101111111: data <= 32'hba5929bb;
    11'b01110000000: data <= 32'h3d06b859;
    11'b01110000001: data <= 32'h3e23b0dc;
    11'b01110000010: data <= 32'h373c31b8;
    11'b01110000011: data <= 32'h335233c8;
    11'b01110000100: data <= 32'h3d813a1d;
    11'b01110000101: data <= 32'h3fdc3df8;
    11'b01110000110: data <= 32'h39b83c1b;
    11'b01110000111: data <= 32'hbbe5bad0;
    11'b01110001000: data <= 32'hbcb2c082;
    11'b01110001001: data <= 32'hab1dbecc;
    11'b01110001010: data <= 32'h39a1b5a2;
    11'b01110001011: data <= 32'h3897b495;
    11'b01110001100: data <= 32'h360dbd21;
    11'b01110001101: data <= 32'h34eebccf;
    11'b01110001110: data <= 32'hb724387e;
    11'b01110001111: data <= 32'hbf3c3fcb;
    11'b01110010000: data <= 32'hc08a3ce4;
    11'b01110010001: data <= 32'hbc6fb83b;
    11'b01110010010: data <= 32'h32b5bc6b;
    11'b01110010011: data <= 32'h2f98b348;
    11'b01110010100: data <= 32'hb8b0391a;
    11'b01110010101: data <= 32'h9a483ab5;
    11'b01110010110: data <= 32'h3eb73c69;
    11'b01110010111: data <= 32'h40573e80;
    11'b01110011000: data <= 32'h38293d9a;
    11'b01110011001: data <= 32'hbd1b2de4;
    11'b01110011010: data <= 32'hbc2bbbd6;
    11'b01110011011: data <= 32'h390eba32;
    11'b01110011100: data <= 32'h3e42b47f;
    11'b01110011101: data <= 32'h3c92bb40;
    11'b01110011110: data <= 32'h38d8bfc3;
    11'b01110011111: data <= 32'h38adbdba;
    11'b01110100000: data <= 32'h33c638c7;
    11'b01110100001: data <= 32'hbab53edc;
    11'b01110100010: data <= 32'hbe72376d;
    11'b01110100011: data <= 32'hbd1cbdfb;
    11'b01110100100: data <= 32'hb9b0befd;
    11'b01110100101: data <= 32'hbb6eb623;
    11'b01110100110: data <= 32'hbcb738f0;
    11'b01110100111: data <= 32'hb0a53835;
    11'b01110101000: data <= 32'h3df23828;
    11'b01110101001: data <= 32'h3e2e3d23;
    11'b01110101010: data <= 32'hb59c3f40;
    11'b01110101011: data <= 32'hbf613cf1;
    11'b01110101100: data <= 32'hbc1534f3;
    11'b01110101101: data <= 32'h3baa2638;
    11'b01110101110: data <= 32'h3ec6ae03;
    11'b01110101111: data <= 32'h3ba4bb25;
    11'b01110110000: data <= 32'h3839be83;
    11'b01110110001: data <= 32'h3c91bac1;
    11'b01110110010: data <= 32'h3de63bc2;
    11'b01110110011: data <= 32'h381e3df5;
    11'b01110110100: data <= 32'hba68b204;
    11'b01110110101: data <= 32'hbcd5c012;
    11'b01110110110: data <= 32'hbbf1bf96;
    11'b01110110111: data <= 32'hbc1eb732;
    11'b01110111000: data <= 32'hbbd72d9a;
    11'b01110111001: data <= 32'ha7b3b8de;
    11'b01110111010: data <= 32'h3c5eb9cf;
    11'b01110111011: data <= 32'h398038f8;
    11'b01110111100: data <= 32'hbcaa3ff8;
    11'b01110111101: data <= 32'hc06d3f8d;
    11'b01110111110: data <= 32'hbc633abb;
    11'b01110111111: data <= 32'h3917326a;
    11'b01111000000: data <= 32'h3ad023cb;
    11'b01111000001: data <= 32'ha847b6b7;
    11'b01111000010: data <= 32'h2e28b9e5;
    11'b01111000011: data <= 32'h3e6f2914;
    11'b01111000100: data <= 32'h40fe3d8c;
    11'b01111000101: data <= 32'h3db43dd0;
    11'b01111000110: data <= 32'hb5a4b23c;
    11'b01111000111: data <= 32'hbc04be7f;
    11'b01111001000: data <= 32'hb8acbd14;
    11'b01111001001: data <= 32'hb46eb430;
    11'b01111001010: data <= 32'hb335b8c1;
    11'b01111001011: data <= 32'h3437bf95;
    11'b01111001100: data <= 32'h3ac7bf9a;
    11'b01111001101: data <= 32'h35102989;
    11'b01111001110: data <= 32'hbcd73f78;
    11'b01111001111: data <= 32'hbfdd3ee0;
    11'b01111010000: data <= 32'hbc6e3614;
    11'b01111010001: data <= 32'haf97b4af;
    11'b01111010010: data <= 32'hb80faa80;
    11'b01111010011: data <= 32'hbd302cd5;
    11'b01111010100: data <= 32'hb77fa905;
    11'b01111010101: data <= 32'h3ed13748;
    11'b01111010110: data <= 32'h416e3dba;
    11'b01111010111: data <= 32'h3d7d3e3e;
    11'b01111011000: data <= 32'hb8403792;
    11'b01111011001: data <= 32'hbac7b68d;
    11'b01111011010: data <= 32'h2f51afa3;
    11'b01111011011: data <= 32'h39303139;
    11'b01111011100: data <= 32'h3697bbd4;
    11'b01111011101: data <= 32'h36f6c11f;
    11'b01111011110: data <= 32'h3b36c099;
    11'b01111011111: data <= 32'h3a04acfb;
    11'b01111100000: data <= 32'hb4e53e54;
    11'b01111100001: data <= 32'hbc5d3bb5;
    11'b01111100010: data <= 32'hbb4eb8ec;
    11'b01111100011: data <= 32'hba42bbe6;
    11'b01111100100: data <= 32'hbe3bb1a6;
    11'b01111100101: data <= 32'hc02d3366;
    11'b01111100110: data <= 32'hba86b004;
    11'b01111100111: data <= 32'h3db8aaea;
    11'b01111101000: data <= 32'h40353b2c;
    11'b01111101001: data <= 32'h38103e74;
    11'b01111101010: data <= 32'hbc843d62;
    11'b01111101011: data <= 32'hba7f3b06;
    11'b01111101100: data <= 32'h389a3b3f;
    11'b01111101101: data <= 32'h3bcc38d4;
    11'b01111101110: data <= 32'h34dfbacc;
    11'b01111101111: data <= 32'h3227c089;
    11'b01111110000: data <= 32'h3c7abf06;
    11'b01111110001: data <= 32'h3ed634b8;
    11'b01111110010: data <= 32'h3c283d64;
    11'b01111110011: data <= 32'ha88c32c1;
    11'b01111110100: data <= 32'hb860bd4c;
    11'b01111110101: data <= 32'hbb4fbce4;
    11'b01111110110: data <= 32'hbebcaf19;
    11'b01111110111: data <= 32'hbfe42192;
    11'b01111111000: data <= 32'hb9e9bbec;
    11'b01111111001: data <= 32'h3c17bd22;
    11'b01111111010: data <= 32'h3cb3a529;
    11'b01111111011: data <= 32'hb72b3ddb;
    11'b01111111100: data <= 32'hbe583f44;
    11'b01111111101: data <= 32'hba503dc2;
    11'b01111111110: data <= 32'h38393cd6;
    11'b01111111111: data <= 32'h36433a63;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    