
module memory_rom_38(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbde138b1;
    11'b00000000001: data <= 32'hba81362b;
    11'b00000000010: data <= 32'h3afdb4fc;
    11'b00000000011: data <= 32'h3f76314c;
    11'b00000000100: data <= 32'h3a463e26;
    11'b00000000101: data <= 32'hbc3c4033;
    11'b00000000110: data <= 32'hbcfd3d75;
    11'b00000000111: data <= 32'h35003734;
    11'b00000001000: data <= 32'h3d69a15d;
    11'b00000001001: data <= 32'h3995b90d;
    11'b00000001010: data <= 32'haee2be25;
    11'b00000001011: data <= 32'h38b8be2c;
    11'b00000001100: data <= 32'h3fa4af8b;
    11'b00000001101: data <= 32'h3f4f3ca4;
    11'b00000001110: data <= 32'h32ee3889;
    11'b00000001111: data <= 32'hbcb2bc75;
    11'b00000010000: data <= 32'hbd97be61;
    11'b00000010001: data <= 32'hbcd8b782;
    11'b00000010010: data <= 32'hbccd33eb;
    11'b00000010011: data <= 32'hb9fdb932;
    11'b00000010100: data <= 32'h3604be67;
    11'b00000010101: data <= 32'h3b66b958;
    11'b00000010110: data <= 32'haaaf3de2;
    11'b00000010111: data <= 32'hbd7840ff;
    11'b00000011000: data <= 32'hbcc73ed7;
    11'b00000011001: data <= 32'h303b388f;
    11'b00000011010: data <= 32'h389631c0;
    11'b00000011011: data <= 32'hb5f19e57;
    11'b00000011100: data <= 32'hba01b824;
    11'b00000011101: data <= 32'h3a55b8ea;
    11'b00000011110: data <= 32'h4166342a;
    11'b00000011111: data <= 32'h41323c24;
    11'b00000100000: data <= 32'h393a377e;
    11'b00000100001: data <= 32'hbad1b9dc;
    11'b00000100010: data <= 32'hba59bb06;
    11'b00000100011: data <= 32'hb480ac67;
    11'b00000100100: data <= 32'hb5d9b18d;
    11'b00000100101: data <= 32'hb7b3beee;
    11'b00000100110: data <= 32'h2a8ec165;
    11'b00000100111: data <= 32'h37c3bd38;
    11'b00000101000: data <= 32'hae9d3cb5;
    11'b00000101001: data <= 32'hbc244035;
    11'b00000101010: data <= 32'hbc183c2c;
    11'b00000101011: data <= 32'hb665a7b7;
    11'b00000101100: data <= 32'hb8f7303c;
    11'b00000101101: data <= 32'hbe7138ac;
    11'b00000101110: data <= 32'hbdc73438;
    11'b00000101111: data <= 32'h394bb208;
    11'b00000110000: data <= 32'h41583357;
    11'b00000110001: data <= 32'h40b03bff;
    11'b00000110010: data <= 32'h35fb3bc8;
    11'b00000110011: data <= 32'hb95b35f1;
    11'b00000110100: data <= 32'h25e834a6;
    11'b00000110101: data <= 32'h3a243837;
    11'b00000110110: data <= 32'h3510b4ab;
    11'b00000110111: data <= 32'hb5d6c046;
    11'b00000111000: data <= 32'ha0f2c1d8;
    11'b00000111001: data <= 32'h3a77bd7b;
    11'b00000111010: data <= 32'h39fa3aa8;
    11'b00000111011: data <= 32'haec93cd0;
    11'b00000111100: data <= 32'hb92daf3f;
    11'b00000111101: data <= 32'hba5dba88;
    11'b00000111110: data <= 32'hbdab26ee;
    11'b00000111111: data <= 32'hc0863ab1;
    11'b00001000000: data <= 32'hbf31344c;
    11'b00001000001: data <= 32'h3432b970;
    11'b00001000010: data <= 32'h3f7fb637;
    11'b00001000011: data <= 32'h3d2d3b02;
    11'b00001000100: data <= 32'hb5843e72;
    11'b00001000101: data <= 32'hb9293dc7;
    11'b00001000110: data <= 32'h38873cdd;
    11'b00001000111: data <= 32'h3cc13c1f;
    11'b00001001000: data <= 32'h335b2789;
    11'b00001001001: data <= 32'hb98dbe6f;
    11'b00001001010: data <= 32'h2984c05a;
    11'b00001001011: data <= 32'h3e4ebb09;
    11'b00001001100: data <= 32'h3fc638e3;
    11'b00001001101: data <= 32'h3b4035f4;
    11'b00001001110: data <= 32'hb196bb75;
    11'b00001001111: data <= 32'hb988bc6b;
    11'b00001010000: data <= 32'hbd1330ce;
    11'b00001010001: data <= 32'hbfbe3a12;
    11'b00001010010: data <= 32'hbe84b71c;
    11'b00001010011: data <= 32'hb161bf49;
    11'b00001010100: data <= 32'h3abdbd4c;
    11'b00001010101: data <= 32'h32b338a9;
    11'b00001010110: data <= 32'hbb1c3f57;
    11'b00001010111: data <= 32'hb8e43eec;
    11'b00001011000: data <= 32'h38ff3d45;
    11'b00001011001: data <= 32'h39d93cac;
    11'b00001011010: data <= 32'hb96e38e2;
    11'b00001011011: data <= 32'hbdc2b81b;
    11'b00001011100: data <= 32'ha1fabc17;
    11'b00001011101: data <= 32'h404eb442;
    11'b00001011110: data <= 32'h414b383c;
    11'b00001011111: data <= 32'h3d732b96;
    11'b00001100000: data <= 32'h30ebbaf6;
    11'b00001100001: data <= 32'hae48b883;
    11'b00001100010: data <= 32'hb45a392a;
    11'b00001100011: data <= 32'hbb3c38e4;
    11'b00001100100: data <= 32'hbc8cbd26;
    11'b00001100101: data <= 32'hb6dfc1b0;
    11'b00001100110: data <= 32'h32d8c008;
    11'b00001100111: data <= 32'hb1133329;
    11'b00001101000: data <= 32'hba063da6;
    11'b00001101001: data <= 32'hb5ce3c03;
    11'b00001101010: data <= 32'h35f53872;
    11'b00001101011: data <= 32'hb26e3b5c;
    11'b00001101100: data <= 32'hbf593c83;
    11'b00001101101: data <= 32'hc06f36ec;
    11'b00001101110: data <= 32'hb42db495;
    11'b00001101111: data <= 32'h401dad10;
    11'b00001110000: data <= 32'h40ac3711;
    11'b00001110001: data <= 32'h3bb03498;
    11'b00001110010: data <= 32'h3179a9df;
    11'b00001110011: data <= 32'h3931381c;
    11'b00001110100: data <= 32'h3b5d3d66;
    11'b00001110101: data <= 32'h2cf63949;
    11'b00001110110: data <= 32'hba46be58;
    11'b00001110111: data <= 32'hb818c208;
    11'b00001111000: data <= 32'h3457c001;
    11'b00001111001: data <= 32'h365897c6;
    11'b00001111010: data <= 32'h2c753885;
    11'b00001111011: data <= 32'h3050b484;
    11'b00001111100: data <= 32'h31e6b81d;
    11'b00001111101: data <= 32'hbadd388b;
    11'b00001111110: data <= 32'hc0e23d7e;
    11'b00001111111: data <= 32'hc113397e;
    11'b00010000000: data <= 32'hb8bdb782;
    11'b00010000001: data <= 32'h3d2ab889;
    11'b00010000010: data <= 32'h3cae3250;
    11'b00010000011: data <= 32'ha52d3981;
    11'b00010000100: data <= 32'haa763adc;
    11'b00010000101: data <= 32'h3ca73d99;
    11'b00010000110: data <= 32'h3e4b3f78;
    11'b00010000111: data <= 32'h34f03bc2;
    11'b00010001000: data <= 32'hbba7bc40;
    11'b00010001001: data <= 32'hb888c056;
    11'b00010001010: data <= 32'h3a44bd1b;
    11'b00010001011: data <= 32'h3d9421cd;
    11'b00010001100: data <= 32'h3c2cb332;
    11'b00010001101: data <= 32'h3952bd45;
    11'b00010001110: data <= 32'h3554bc82;
    11'b00010001111: data <= 32'hb983380d;
    11'b00010010000: data <= 32'hc0103d87;
    11'b00010010001: data <= 32'hc0593395;
    11'b00010010010: data <= 32'hba7dbd8d;
    11'b00010010011: data <= 32'h34e4bdd5;
    11'b00010010100: data <= 32'haf98b1fe;
    11'b00010010101: data <= 32'hbb273a82;
    11'b00010010110: data <= 32'hb3423c60;
    11'b00010010111: data <= 32'h3d233dbf;
    11'b00010011000: data <= 32'h3d853f6d;
    11'b00010011001: data <= 32'hb5aa3d7f;
    11'b00010011010: data <= 32'hbe93a245;
    11'b00010011011: data <= 32'hb9deba9a;
    11'b00010011100: data <= 32'h3cdfb55b;
    11'b00010011101: data <= 32'h400b312a;
    11'b00010011110: data <= 32'h3dd1b89d;
    11'b00010011111: data <= 32'h3b30be14;
    11'b00010100000: data <= 32'h3a5dbad8;
    11'b00010100001: data <= 32'h345b3b62;
    11'b00010100010: data <= 32'hbaa23d6c;
    11'b00010100011: data <= 32'hbd74b6d9;
    11'b00010100100: data <= 32'hba9ec09d;
    11'b00010100101: data <= 32'hb574c03d;
    11'b00010100110: data <= 32'hb9feb808;
    11'b00010100111: data <= 32'hbc343784;
    11'b00010101000: data <= 32'had5c3631;
    11'b00010101001: data <= 32'h3c9c3832;
    11'b00010101010: data <= 32'h39383d40;
    11'b00010101011: data <= 32'hbd8a3e94;
    11'b00010101100: data <= 32'hc0ce3b7a;
    11'b00010101101: data <= 32'hbbea3178;
    11'b00010101110: data <= 32'h3c983171;
    11'b00010101111: data <= 32'h3eda32c4;
    11'b00010110000: data <= 32'h3b68b75e;
    11'b00010110001: data <= 32'h393fbb5d;
    11'b00010110010: data <= 32'h3d3c2c7d;
    11'b00010110011: data <= 32'h3dd13e73;
    11'b00010110100: data <= 32'h367f3dcf;
    11'b00010110101: data <= 32'hb961b9a6;
    11'b00010110110: data <= 32'hb9e7c0ee;
    11'b00010110111: data <= 32'hb613c002;
    11'b00010111000: data <= 32'hb700b81d;
    11'b00010111001: data <= 32'hb68eb16d;
    11'b00010111010: data <= 32'h3654bb13;
    11'b00010111011: data <= 32'h3c2dba50;
    11'b00010111100: data <= 32'h2b9638e6;
    11'b00010111101: data <= 32'hbfd93ec0;
    11'b00010111110: data <= 32'hc14d3d10;
    11'b00010111111: data <= 32'hbc9e33df;
    11'b00011000000: data <= 32'h3872ae91;
    11'b00011000001: data <= 32'h387814c5;
    11'b00011000010: data <= 32'hb490b12c;
    11'b00011000011: data <= 32'h2d81afb0;
    11'b00011000100: data <= 32'h3e683b4e;
    11'b00011000101: data <= 32'h4055402c;
    11'b00011000110: data <= 32'h3b403e98;
    11'b00011000111: data <= 32'hb8bfb517;
    11'b00011001000: data <= 32'hb9dbbe82;
    11'b00011001001: data <= 32'h2511bc47;
    11'b00011001010: data <= 32'h36c2b145;
    11'b00011001011: data <= 32'h3805b9d5;
    11'b00011001100: data <= 32'h3b43bfde;
    11'b00011001101: data <= 32'h3c88beb8;
    11'b00011001110: data <= 32'h3045343e;
    11'b00011001111: data <= 32'hbe3c3e6b;
    11'b00011010000: data <= 32'hc0343b6f;
    11'b00011010001: data <= 32'hbc3eb807;
    11'b00011010010: data <= 32'hb270bb42;
    11'b00011010011: data <= 32'hba26b615;
    11'b00011010100: data <= 32'hbdc7a67a;
    11'b00011010101: data <= 32'hb6803169;
    11'b00011010110: data <= 32'h3e633ba6;
    11'b00011010111: data <= 32'h402a3fb5;
    11'b00011011000: data <= 32'h370b3f19;
    11'b00011011001: data <= 32'hbca7381f;
    11'b00011011010: data <= 32'hbb30b401;
    11'b00011011011: data <= 32'h36ce312a;
    11'b00011011100: data <= 32'h3c3e3536;
    11'b00011011101: data <= 32'h3b54bb69;
    11'b00011011110: data <= 32'h3c1ec08a;
    11'b00011011111: data <= 32'h3d74be86;
    11'b00011100000: data <= 32'h3b2d383c;
    11'b00011100001: data <= 32'hb5453e46;
    11'b00011100010: data <= 32'hbc083523;
    11'b00011100011: data <= 32'hb9c4bd96;
    11'b00011100100: data <= 32'hb959be43;
    11'b00011100101: data <= 32'hbdfcb8fc;
    11'b00011100110: data <= 32'hbf67b20d;
    11'b00011100111: data <= 32'hb745b5de;
    11'b00011101000: data <= 32'h3dc02675;
    11'b00011101001: data <= 32'h3db83c77;
    11'b00011101010: data <= 32'hb83f3ebf;
    11'b00011101011: data <= 32'hbfa23d0f;
    11'b00011101100: data <= 32'hbc723ab4;
    11'b00011101101: data <= 32'h37c53b8a;
    11'b00011101110: data <= 32'h3b2438e0;
    11'b00011101111: data <= 32'h360aba14;
    11'b00011110000: data <= 32'h3862bf0b;
    11'b00011110001: data <= 32'h3e21ba64;
    11'b00011110010: data <= 32'h3f7f3cc2;
    11'b00011110011: data <= 32'h3bf13e94;
    11'b00011110100: data <= 32'ha4d9a913;
    11'b00011110101: data <= 32'hb5aebea8;
    11'b00011110110: data <= 32'hb909bdcb;
    11'b00011110111: data <= 32'hbd24b6dd;
    11'b00011111000: data <= 32'hbd5bb816;
    11'b00011111001: data <= 32'ha73cbdbd;
    11'b00011111010: data <= 32'h3d4cbd79;
    11'b00011111011: data <= 32'h3a5b2ea4;
    11'b00011111100: data <= 32'hbcc13dac;
    11'b00011111101: data <= 32'hc0543df5;
    11'b00011111110: data <= 32'hbc723c17;
    11'b00011111111: data <= 32'h318e3ab7;
    11'b00100000000: data <= 32'hac5b37c6;
    11'b00100000001: data <= 32'hbb3fb75c;
    11'b00100000010: data <= 32'hb564bba0;
    11'b00100000011: data <= 32'h3df32e26;
    11'b00100000100: data <= 32'h40e83eb7;
    11'b00100000101: data <= 32'h3e6e3edd;
    11'b00100000110: data <= 32'h34562ed9;
    11'b00100000111: data <= 32'hb30cbc06;
    11'b00100001000: data <= 32'hb31ab733;
    11'b00100001001: data <= 32'hb72b334b;
    11'b00100001010: data <= 32'hb682b9c5;
    11'b00100001011: data <= 32'h3804c0bb;
    11'b00100001100: data <= 32'h3d4fc0c2;
    11'b00100001101: data <= 32'h395ab7e0;
    11'b00100001110: data <= 32'hbb9b3ca1;
    11'b00100001111: data <= 32'hbe443c83;
    11'b00100010000: data <= 32'hb9d23521;
    11'b00100010001: data <= 32'hb3882a87;
    11'b00100010010: data <= 32'hbcf02de7;
    11'b00100010011: data <= 32'hc060b453;
    11'b00100010100: data <= 32'hbc72b80e;
    11'b00100010101: data <= 32'h3d0b34a3;
    11'b00100010110: data <= 32'h40a53df6;
    11'b00100010111: data <= 32'h3cd73e53;
    11'b00100011000: data <= 32'hb3c238d5;
    11'b00100011001: data <= 32'hb6163295;
    11'b00100011010: data <= 32'h32d63b41;
    11'b00100011011: data <= 32'h34e63c1c;
    11'b00100011100: data <= 32'h3083b942;
    11'b00100011101: data <= 32'h38f1c134;
    11'b00100011110: data <= 32'h3d57c0d6;
    11'b00100011111: data <= 32'h3c78b544;
    11'b00100100000: data <= 32'h2f1c3c58;
    11'b00100100001: data <= 32'hb5983802;
    11'b00100100010: data <= 32'habbbb936;
    11'b00100100011: data <= 32'hb68ab9c2;
    11'b00100100100: data <= 32'hbf84b13a;
    11'b00100100101: data <= 32'hc168b411;
    11'b00100100110: data <= 32'hbd3bba0d;
    11'b00100100111: data <= 32'h3c1fb78c;
    11'b00100101000: data <= 32'h3e9d388c;
    11'b00100101001: data <= 32'h32243ca5;
    11'b00100101010: data <= 32'hbc4d3c25;
    11'b00100101011: data <= 32'hb8f03cc9;
    11'b00100101100: data <= 32'h369c3f45;
    11'b00100101101: data <= 32'h36423e08;
    11'b00100101110: data <= 32'hb359b607;
    11'b00100101111: data <= 32'h29c1c025;
    11'b00100110000: data <= 32'h3cb9be45;
    11'b00100110001: data <= 32'h3f0f3639;
    11'b00100110010: data <= 32'h3d4b3cc2;
    11'b00100110011: data <= 32'h3a4c2882;
    11'b00100110100: data <= 32'h3866bc8e;
    11'b00100110101: data <= 32'hb2c2ba25;
    11'b00100110110: data <= 32'hbe8f2e39;
    11'b00100110111: data <= 32'hc069b46a;
    11'b00100111000: data <= 32'hbae0bdfa;
    11'b00100111001: data <= 32'h3b7ebefb;
    11'b00100111010: data <= 32'h3b83b8d1;
    11'b00100111011: data <= 32'hb93b38da;
    11'b00100111100: data <= 32'hbdf73c3b;
    11'b00100111101: data <= 32'hb89e3d60;
    11'b00100111110: data <= 32'h35ec3f0d;
    11'b00100111111: data <= 32'hb3f93da2;
    11'b00101000000: data <= 32'hbd8aad14;
    11'b00101000001: data <= 32'hbbfebcd2;
    11'b00101000010: data <= 32'h3a92b81d;
    11'b00101000011: data <= 32'h40353c22;
    11'b00101000100: data <= 32'h3f913cfc;
    11'b00101000101: data <= 32'h3ca4aac5;
    11'b00101000110: data <= 32'h3a18ba49;
    11'b00101000111: data <= 32'h331b2e11;
    11'b00101001000: data <= 32'hba0f3b40;
    11'b00101001001: data <= 32'hbc96b108;
    11'b00101001010: data <= 32'hb1f0c050;
    11'b00101001011: data <= 32'h3b93c166;
    11'b00101001100: data <= 32'h38e8bd41;
    11'b00101001101: data <= 32'hb9a332cd;
    11'b00101001110: data <= 32'hbc273912;
    11'b00101001111: data <= 32'hab3c38d7;
    11'b00101010000: data <= 32'h34ac3b10;
    11'b00101010001: data <= 32'hbc843b24;
    11'b00101010010: data <= 32'hc1362d9a;
    11'b00101010011: data <= 32'hbfacb8be;
    11'b00101010100: data <= 32'h3684aa62;
    11'b00101010101: data <= 32'h3f793c00;
    11'b00101010110: data <= 32'h3dd83bfb;
    11'b00101010111: data <= 32'h38c12fcc;
    11'b00101011000: data <= 32'h381a3027;
    11'b00101011001: data <= 32'h390d3d89;
    11'b00101011010: data <= 32'h30453f7d;
    11'b00101011011: data <= 32'hb593308b;
    11'b00101011100: data <= 32'h2e45c080;
    11'b00101011101: data <= 32'h3af6c16a;
    11'b00101011110: data <= 32'h3a0ebc8e;
    11'b00101011111: data <= 32'h2b1f31f5;
    11'b00101100000: data <= 32'h2e92261d;
    11'b00101100001: data <= 32'h3a55b7a9;
    11'b00101100010: data <= 32'h3647af57;
    11'b00101100011: data <= 32'hbe633762;
    11'b00101100100: data <= 32'hc22f30fb;
    11'b00101100101: data <= 32'hc04ab87f;
    11'b00101100110: data <= 32'h3177b811;
    11'b00101100111: data <= 32'h3cc83165;
    11'b00101101000: data <= 32'h3596364a;
    11'b00101101001: data <= 32'hb6ff3409;
    11'b00101101010: data <= 32'h2e883b53;
    11'b00101101011: data <= 32'h3ad6408b;
    11'b00101101100: data <= 32'h378340db;
    11'b00101101101: data <= 32'hb6af37b6;
    11'b00101101110: data <= 32'hb5dbbec3;
    11'b00101101111: data <= 32'h3855bf1d;
    11'b00101110000: data <= 32'h3c58b410;
    11'b00101110001: data <= 32'h3c283738;
    11'b00101110010: data <= 32'h3ce1b725;
    11'b00101110011: data <= 32'h3e15bcc2;
    11'b00101110100: data <= 32'h39a4b757;
    11'b00101110101: data <= 32'hbd3338bc;
    11'b00101110110: data <= 32'hc10f3498;
    11'b00101110111: data <= 32'hbe45bbd3;
    11'b00101111000: data <= 32'h32ecbe22;
    11'b00101111001: data <= 32'h37c7bbd8;
    11'b00101111010: data <= 32'hb991b514;
    11'b00101111011: data <= 32'hbc912ead;
    11'b00101111100: data <= 32'ha0183bcf;
    11'b00101111101: data <= 32'h3b804057;
    11'b00101111110: data <= 32'h309a407c;
    11'b00101111111: data <= 32'hbd3d3963;
    11'b00110000000: data <= 32'hbd86baa2;
    11'b00110000001: data <= 32'h1629b860;
    11'b00110000010: data <= 32'h3cd5395a;
    11'b00110000011: data <= 32'h3df73965;
    11'b00110000100: data <= 32'h3e42b90e;
    11'b00110000101: data <= 32'h3eccbc8d;
    11'b00110000110: data <= 32'h3c4e3027;
    11'b00110000111: data <= 32'hb6ab3d6e;
    11'b00110001000: data <= 32'hbd4138c7;
    11'b00110001001: data <= 32'hb909bd8d;
    11'b00110001010: data <= 32'h3679c0b0;
    11'b00110001011: data <= 32'h2dbfbeb8;
    11'b00110001100: data <= 32'hbc23b9dc;
    11'b00110001101: data <= 32'hbbcab4f5;
    11'b00110001110: data <= 32'h37343327;
    11'b00110001111: data <= 32'h3c333ca0;
    11'b00110010000: data <= 32'hb75a3df4;
    11'b00110010001: data <= 32'hc0ba3946;
    11'b00110010010: data <= 32'hc099b163;
    11'b00110010011: data <= 32'hb7c3321c;
    11'b00110010100: data <= 32'h3b6a3b76;
    11'b00110010101: data <= 32'h3c1d381a;
    11'b00110010110: data <= 32'h3b1fb91a;
    11'b00110010111: data <= 32'h3cfdb81c;
    11'b00110011000: data <= 32'h3d433cef;
    11'b00110011001: data <= 32'h380a40a9;
    11'b00110011010: data <= 32'hb41f3c0d;
    11'b00110011011: data <= 32'ha911bd88;
    11'b00110011100: data <= 32'h3717c099;
    11'b00110011101: data <= 32'h2c77bdb1;
    11'b00110011110: data <= 32'hb898b8d0;
    11'b00110011111: data <= 32'ha8beba32;
    11'b00110100000: data <= 32'h3d3bbb0f;
    11'b00110100001: data <= 32'h3d35ad37;
    11'b00110100010: data <= 32'hba4339fa;
    11'b00110100011: data <= 32'hc18f38ae;
    11'b00110100100: data <= 32'hc0f119a3;
    11'b00110100101: data <= 32'hb8ef28d0;
    11'b00110100110: data <= 32'h35cf353b;
    11'b00110100111: data <= 32'haeb7adff;
    11'b00110101000: data <= 32'hb5c9b978;
    11'b00110101001: data <= 32'h38402db4;
    11'b00110101010: data <= 32'h3d7f4011;
    11'b00110101011: data <= 32'h3ba741b8;
    11'b00110101100: data <= 32'ha57c3d36;
    11'b00110101101: data <= 32'hb409bb1e;
    11'b00110101110: data <= 32'h302ebd61;
    11'b00110101111: data <= 32'h32b2b572;
    11'b00110110000: data <= 32'h322faa0f;
    11'b00110110001: data <= 32'h3bd1bc48;
    11'b00110110010: data <= 32'h4012bebf;
    11'b00110110011: data <= 32'h3e7bb9d3;
    11'b00110110100: data <= 32'hb80e38cf;
    11'b00110110101: data <= 32'hc05f3962;
    11'b00110110110: data <= 32'hbee4b322;
    11'b00110110111: data <= 32'hb4eeb9f5;
    11'b00110111000: data <= 32'hb195b99c;
    11'b00110111001: data <= 32'hbceaba99;
    11'b00110111010: data <= 32'hbd74bb1f;
    11'b00110111011: data <= 32'h2fef3000;
    11'b00110111100: data <= 32'h3d883f95;
    11'b00110111101: data <= 32'h3a7f4113;
    11'b00110111110: data <= 32'hb9323d13;
    11'b00110111111: data <= 32'hbc7eb1ff;
    11'b00111000000: data <= 32'hb70ba9a9;
    11'b00111000001: data <= 32'h33433afe;
    11'b00111000010: data <= 32'h389d37d3;
    11'b00111000011: data <= 32'h3d20bc9c;
    11'b00111000100: data <= 32'h403bbf35;
    11'b00111000101: data <= 32'h3f40b6b7;
    11'b00111000110: data <= 32'h33a33cc9;
    11'b00111000111: data <= 32'hbb423c0c;
    11'b00111001000: data <= 32'hb808b7ea;
    11'b00111001001: data <= 32'h327abdc9;
    11'b00111001010: data <= 32'hb718bd6a;
    11'b00111001011: data <= 32'hbee1bcb9;
    11'b00111001100: data <= 32'hbdf5bcba;
    11'b00111001101: data <= 32'h361db828;
    11'b00111001110: data <= 32'h3e0c3a9d;
    11'b00111001111: data <= 32'h35e33e13;
    11'b00111010000: data <= 32'hbe3c3b77;
    11'b00111010001: data <= 32'hbff13543;
    11'b00111010010: data <= 32'hbb3c3aaf;
    11'b00111010011: data <= 32'h216e3dc8;
    11'b00111010100: data <= 32'h31f03879;
    11'b00111010101: data <= 32'h3878bc9e;
    11'b00111010110: data <= 32'h3db7bd66;
    11'b00111010111: data <= 32'h3efb3813;
    11'b00111011000: data <= 32'h3c064034;
    11'b00111011001: data <= 32'h347a3dbc;
    11'b00111011010: data <= 32'h3683b800;
    11'b00111011011: data <= 32'h380bbdbd;
    11'b00111011100: data <= 32'hb6f3bc38;
    11'b00111011101: data <= 32'hbdbfbad2;
    11'b00111011110: data <= 32'hba0cbd79;
    11'b00111011111: data <= 32'h3c9ebde4;
    11'b00111100000: data <= 32'h3f28b83f;
    11'b00111100001: data <= 32'h2d393731;
    11'b00111100010: data <= 32'hbfe33882;
    11'b00111100011: data <= 32'hc03e3716;
    11'b00111100100: data <= 32'hbb0a3ae3;
    11'b00111100101: data <= 32'hb5133c49;
    11'b00111100110: data <= 32'hba732bca;
    11'b00111100111: data <= 32'hba6bbcf2;
    11'b00111101000: data <= 32'h3630ba93;
    11'b00111101001: data <= 32'h3df23d19;
    11'b00111101010: data <= 32'h3d7e4133;
    11'b00111101011: data <= 32'h398d3e72;
    11'b00111101100: data <= 32'h374eb238;
    11'b00111101101: data <= 32'h3556b8d0;
    11'b00111101110: data <= 32'hb549300f;
    11'b00111101111: data <= 32'hba3623de;
    11'b00111110000: data <= 32'h322dbd5a;
    11'b00111110001: data <= 32'h3f6fc057;
    11'b00111110010: data <= 32'h4014bd69;
    11'b00111110011: data <= 32'h33082250;
    11'b00111110100: data <= 32'hbde9378e;
    11'b00111110101: data <= 32'hbd2433b5;
    11'b00111110110: data <= 32'hb47c32c2;
    11'b00111110111: data <= 32'hb8443084;
    11'b00111111000: data <= 32'hbf3fb928;
    11'b00111111001: data <= 32'hbfe7bda8;
    11'b00111111010: data <= 32'hb564b996;
    11'b00111111011: data <= 32'h3d193cda;
    11'b00111111100: data <= 32'h3cee4069;
    11'b00111111101: data <= 32'h32f03d44;
    11'b00111111110: data <= 32'hb4803282;
    11'b00111111111: data <= 32'hb271389f;
    11'b01000000000: data <= 32'hb50a3e09;
    11'b01000000001: data <= 32'hb5a63b19;
    11'b01000000010: data <= 32'h386abca8;
    11'b01000000011: data <= 32'h3f8bc088;
    11'b01000000100: data <= 32'h4005bcd5;
    11'b01000000101: data <= 32'h398036ff;
    11'b01000000110: data <= 32'hb5163a07;
    11'b01000000111: data <= 32'h2e2fa078;
    11'b01000001000: data <= 32'h389eb7cb;
    11'b01000001001: data <= 32'hb823b856;
    11'b01000001010: data <= 32'hc086bbc0;
    11'b01000001011: data <= 32'hc08dbe20;
    11'b01000001100: data <= 32'hb497bc67;
    11'b01000001101: data <= 32'h3d433422;
    11'b01000001110: data <= 32'h3a8a3c23;
    11'b01000001111: data <= 32'hb937390f;
    11'b01000010000: data <= 32'hbc9736a3;
    11'b01000010001: data <= 32'hb9313d9a;
    11'b01000010010: data <= 32'hb6824089;
    11'b01000010011: data <= 32'hb85a3cd1;
    11'b01000010100: data <= 32'hac1abc2b;
    11'b01000010101: data <= 32'h3c40bf5c;
    11'b01000010110: data <= 32'h3e6bb599;
    11'b01000010111: data <= 32'h3c903d45;
    11'b01000011000: data <= 32'h3a673caa;
    11'b01000011001: data <= 32'h3cd3ae0d;
    11'b01000011010: data <= 32'h3caab90c;
    11'b01000011011: data <= 32'hb586b573;
    11'b01000011100: data <= 32'hbffeb83a;
    11'b01000011101: data <= 32'hbe90bda0;
    11'b01000011110: data <= 32'h36dabef8;
    11'b01000011111: data <= 32'h3e55bc16;
    11'b01000100000: data <= 32'h37c6b3c2;
    11'b01000100001: data <= 32'hbcb7ab82;
    11'b01000100010: data <= 32'hbd7a353a;
    11'b01000100011: data <= 32'hb8523dbd;
    11'b01000100100: data <= 32'hb7594009;
    11'b01000100101: data <= 32'hbcf63a68;
    11'b01000100110: data <= 32'hbd5dbc69;
    11'b01000100111: data <= 32'hb1f9bd2c;
    11'b01000101000: data <= 32'h3bfe37dc;
    11'b01000101001: data <= 32'h3d143f8f;
    11'b01000101010: data <= 32'h3cd93d25;
    11'b01000101011: data <= 32'h3da3a572;
    11'b01000101100: data <= 32'h3c89ac5f;
    11'b01000101101: data <= 32'hb25d3a09;
    11'b01000101110: data <= 32'hbd59384f;
    11'b01000101111: data <= 32'hb935bc11;
    11'b01000110000: data <= 32'h3cc4c059;
    11'b01000110001: data <= 32'h3f32bf50;
    11'b01000110010: data <= 32'h36f7bae2;
    11'b01000110011: data <= 32'hbb67b56c;
    11'b01000110100: data <= 32'hb8f82a96;
    11'b01000110101: data <= 32'h33ce3a5d;
    11'b01000110110: data <= 32'hb5143c55;
    11'b01000110111: data <= 32'hbfda2af3;
    11'b01000111000: data <= 32'hc0fbbd10;
    11'b01000111001: data <= 32'hbc75bc18;
    11'b01000111010: data <= 32'h38643922;
    11'b01000111011: data <= 32'h3c123e57;
    11'b01000111100: data <= 32'h39ff3aa2;
    11'b01000111101: data <= 32'h39a0283a;
    11'b01000111110: data <= 32'h38af3a96;
    11'b01000111111: data <= 32'hb1c74036;
    11'b01001000000: data <= 32'hba733e88;
    11'b01001000001: data <= 32'haf10b87a;
    11'b01001000010: data <= 32'h3d41c03d;
    11'b01001000011: data <= 32'h3e8cbecc;
    11'b01001000100: data <= 32'h38acb809;
    11'b01001000101: data <= 32'haa6aad43;
    11'b01001000110: data <= 32'h39ceb279;
    11'b01001000111: data <= 32'h3d5725fd;
    11'b01001001000: data <= 32'h241033f4;
    11'b01001001001: data <= 32'hc075b5e6;
    11'b01001001010: data <= 32'hc19cbd23;
    11'b01001001011: data <= 32'hbcb0bc8e;
    11'b01001001100: data <= 32'h3827a8d0;
    11'b01001001101: data <= 32'h38ad374a;
    11'b01001001110: data <= 32'hb159ade9;
    11'b01001001111: data <= 32'hb480ae3e;
    11'b01001010000: data <= 32'h29363dbd;
    11'b01001010001: data <= 32'hb29e41c2;
    11'b01001010010: data <= 32'hb9fd4030;
    11'b01001010011: data <= 32'hb767b512;
    11'b01001010100: data <= 32'h385abe9b;
    11'b01001010101: data <= 32'h3c02ba7d;
    11'b01001010110: data <= 32'h39763757;
    11'b01001010111: data <= 32'h3ab036ac;
    11'b01001011000: data <= 32'h3f68b539;
    11'b01001011001: data <= 32'h4036b545;
    11'b01001011010: data <= 32'h35c3327d;
    11'b01001011011: data <= 32'hbf941a29;
    11'b01001011100: data <= 32'hc04ebb9a;
    11'b01001011101: data <= 32'hb68fbdb4;
    11'b01001011110: data <= 32'h3ad0bc48;
    11'b01001011111: data <= 32'h3368bab4;
    11'b01001100000: data <= 32'hbaedbc00;
    11'b01001100001: data <= 32'hb9dab68a;
    11'b01001100010: data <= 32'h2c343d7a;
    11'b01001100011: data <= 32'had1f4141;
    11'b01001100100: data <= 32'hbc693ebe;
    11'b01001100101: data <= 32'hbdefb69c;
    11'b01001100110: data <= 32'hb9bfbc5c;
    11'b01001100111: data <= 32'h30ed317e;
    11'b01001101000: data <= 32'h38573cf5;
    11'b01001101001: data <= 32'h3c7a3912;
    11'b01001101010: data <= 32'h4022b660;
    11'b01001101011: data <= 32'h403bad82;
    11'b01001101100: data <= 32'h38133c28;
    11'b01001101101: data <= 32'hbcdd3c4c;
    11'b01001101110: data <= 32'hbc31b4e0;
    11'b01001101111: data <= 32'h3852be36;
    11'b01001110000: data <= 32'h3cb1bee4;
    11'b01001110001: data <= 32'h2c62bdee;
    11'b01001110010: data <= 32'hbb3dbd7d;
    11'b01001110011: data <= 32'hb3b1b9e0;
    11'b01001110100: data <= 32'h3ab7399f;
    11'b01001110101: data <= 32'h350d3e68;
    11'b01001110110: data <= 32'hbdfe3a3a;
    11'b01001110111: data <= 32'hc0e9b97a;
    11'b01001111000: data <= 32'hbebdb9e3;
    11'b01001111001: data <= 32'hb70238b2;
    11'b01001111010: data <= 32'h31f33cc2;
    11'b01001111011: data <= 32'h38e93290;
    11'b01001111100: data <= 32'h3d30b8af;
    11'b01001111101: data <= 32'h3dc3377e;
    11'b01001111110: data <= 32'h36d24065;
    11'b01001111111: data <= 32'hb902406e;
    11'b01010000000: data <= 32'hb44e3569;
    11'b01010000001: data <= 32'h3b53bd5c;
    11'b01010000010: data <= 32'h3c3fbe1d;
    11'b01010000011: data <= 32'h9bbabc5b;
    11'b01010000100: data <= 32'hb5dcbc22;
    11'b01010000101: data <= 32'h3b34bb41;
    11'b01010000110: data <= 32'h3fedaf31;
    11'b01010000111: data <= 32'h3af63872;
    11'b01010001000: data <= 32'hbe3c2ec7;
    11'b01010001001: data <= 32'hc15eba38;
    11'b01010001010: data <= 32'hbeebb942;
    11'b01010001011: data <= 32'hb6fe33a0;
    11'b01010001100: data <= 32'hb25f346f;
    11'b01010001101: data <= 32'hb56cba1e;
    11'b01010001110: data <= 32'h301bbbb2;
    11'b01010001111: data <= 32'h393f3aae;
    11'b01010010000: data <= 32'h34dd41bb;
    11'b01010010001: data <= 32'hb67b4160;
    11'b01010010010: data <= 32'hb4d238d6;
    11'b01010010011: data <= 32'h3601bb04;
    11'b01010010100: data <= 32'h363cb8d2;
    11'b01010010101: data <= 32'hb14027d0;
    11'b01010010110: data <= 32'h33dcb502;
    11'b01010010111: data <= 32'h3fa1bb5f;
    11'b01010011000: data <= 32'h4194b8c8;
    11'b01010011001: data <= 32'h3d2c328c;
    11'b01010011010: data <= 32'hbcbb337e;
    11'b01010011011: data <= 32'hbff3b6d4;
    11'b01010011100: data <= 32'hbab8b97a;
    11'b01010011101: data <= 32'h2d95b7f8;
    11'b01010011110: data <= 32'hb711bb12;
    11'b01010011111: data <= 32'hbc94beee;
    11'b01010100000: data <= 32'hb8e1bd9e;
    11'b01010100001: data <= 32'h36ce3974;
    11'b01010100010: data <= 32'h36b7411f;
    11'b01010100011: data <= 32'hb818405e;
    11'b01010100100: data <= 32'hbc0c35ab;
    11'b01010100101: data <= 32'hb9e9b6a2;
    11'b01010100110: data <= 32'hb8453781;
    11'b01010100111: data <= 32'hb7ba3c53;
    11'b01010101000: data <= 32'h36553157;
    11'b01010101001: data <= 32'h4021bba0;
    11'b01010101010: data <= 32'h4179b8a7;
    11'b01010101011: data <= 32'h3d5639c9;
    11'b01010101100: data <= 32'hb8a83c8e;
    11'b01010101101: data <= 32'hba6f34c4;
    11'b01010101110: data <= 32'h35c7b8c4;
    11'b01010101111: data <= 32'h3964bbcd;
    11'b01010110000: data <= 32'hb850bddb;
    11'b01010110001: data <= 32'hbd8dc02a;
    11'b01010110010: data <= 32'hb704beb4;
    11'b01010110011: data <= 32'h3c0c2c16;
    11'b01010110100: data <= 32'h3b193ddc;
    11'b01010110101: data <= 32'hb9563c30;
    11'b01010110110: data <= 32'hbf17b1ab;
    11'b01010110111: data <= 32'hbe88b0a6;
    11'b01010111000: data <= 32'hbc923c44;
    11'b01010111001: data <= 32'hbac43d67;
    11'b01010111010: data <= 32'hae43aadd;
    11'b01010111011: data <= 32'h3cebbcc7;
    11'b01010111100: data <= 32'h3f73b46c;
    11'b01010111101: data <= 32'h3c073e92;
    11'b01010111110: data <= 32'had914064;
    11'b01010111111: data <= 32'h30673bed;
    11'b01011000000: data <= 32'h3c38b515;
    11'b01011000001: data <= 32'h3a59ba05;
    11'b01011000010: data <= 32'hb924bc0c;
    11'b01011000011: data <= 32'hbc64be52;
    11'b01011000100: data <= 32'h3716be88;
    11'b01011000101: data <= 32'h401eb93b;
    11'b01011000110: data <= 32'h3e0f345e;
    11'b01011000111: data <= 32'hb8e22b75;
    11'b01011001000: data <= 32'hbfbab82d;
    11'b01011001001: data <= 32'hbe7fabec;
    11'b01011001010: data <= 32'hbc163bb0;
    11'b01011001011: data <= 32'hbc3a39b8;
    11'b01011001100: data <= 32'hbbb4bb4f;
    11'b01011001101: data <= 32'hac6bbea3;
    11'b01011001110: data <= 32'h3a29ac6c;
    11'b01011001111: data <= 32'h38ea4068;
    11'b01011010000: data <= 32'h2f16413e;
    11'b01011010001: data <= 32'h35703cbc;
    11'b01011010010: data <= 32'h3a7a2603;
    11'b01011010011: data <= 32'h34082ec2;
    11'b01011010100: data <= 32'hbb293328;
    11'b01011010101: data <= 32'hb96cb88f;
    11'b01011010110: data <= 32'h3d40bd7b;
    11'b01011010111: data <= 32'h41a5bc5d;
    11'b01011011000: data <= 32'h3fa3b4d0;
    11'b01011011001: data <= 32'hb4cfb005;
    11'b01011011010: data <= 32'hbd1ab54c;
    11'b01011011011: data <= 32'hb90c9c6a;
    11'b01011011100: data <= 32'hb375370a;
    11'b01011011101: data <= 32'hbc1db47d;
    11'b01011011110: data <= 32'hbed0bf5a;
    11'b01011011111: data <= 32'hbc11c03a;
    11'b01011100000: data <= 32'h32cbb2c3;
    11'b01011100001: data <= 32'h384d3fa7;
    11'b01011100010: data <= 32'h2c92400d;
    11'b01011100011: data <= 32'hb07a399e;
    11'b01011100100: data <= 32'haf19337f;
    11'b01011100101: data <= 32'hb9003c6c;
    11'b01011100110: data <= 32'hbd0e3de2;
    11'b01011100111: data <= 32'hb88d33e3;
    11'b01011101000: data <= 32'h3dd1bcb6;
    11'b01011101001: data <= 32'h4164bc79;
    11'b01011101010: data <= 32'h3f0ba53d;
    11'b01011101011: data <= 32'h2d133873;
    11'b01011101100: data <= 32'hb12f355c;
    11'b01011101101: data <= 32'h3a0c312f;
    11'b01011101110: data <= 32'h398b2a98;
    11'b01011101111: data <= 32'hbb02ba8f;
    11'b01011110000: data <= 32'hbfdac044;
    11'b01011110001: data <= 32'hbc58c07e;
    11'b01011110010: data <= 32'h3862b92f;
    11'b01011110011: data <= 32'h3b653b05;
    11'b01011110100: data <= 32'h1ef139b8;
    11'b01011110101: data <= 32'hba2cb144;
    11'b01011110110: data <= 32'hbb7f339e;
    11'b01011110111: data <= 32'hbccb3ecb;
    11'b01011111000: data <= 32'hbe273fed;
    11'b01011111001: data <= 32'hbb6c34df;
    11'b01011111010: data <= 32'h395bbd3d;
    11'b01011111011: data <= 32'h3ea7bb3b;
    11'b01011111100: data <= 32'h3c7339e7;
    11'b01011111101: data <= 32'h34d73e13;
    11'b01011111110: data <= 32'h3a163c04;
    11'b01011111111: data <= 32'h3ec43672;
    11'b01100000000: data <= 32'h3c79321b;
    11'b01100000001: data <= 32'hbab2b676;
    11'b01100000010: data <= 32'hbf07bdfd;
    11'b01100000011: data <= 32'hb639bfa2;
    11'b01100000100: data <= 32'h3de3bc65;
    11'b01100000101: data <= 32'h3e22b48f;
    11'b01100000110: data <= 32'h2c7eb821;
    11'b01100000111: data <= 32'hbbb5bab9;
    11'b01100001000: data <= 32'hbb9630a0;
    11'b01100001001: data <= 32'hbbc33ea7;
    11'b01100001010: data <= 32'hbdfb3e33;
    11'b01100001011: data <= 32'hbe2db66d;
    11'b01100001100: data <= 32'hb8bfbefe;
    11'b01100001101: data <= 32'h354fb9e3;
    11'b01100001110: data <= 32'h35e83d26;
    11'b01100001111: data <= 32'h34a83fc9;
    11'b01100010000: data <= 32'h3c133c78;
    11'b01100010001: data <= 32'h3ead384e;
    11'b01100010010: data <= 32'h3a1c3aa2;
    11'b01100010011: data <= 32'hbc343a5a;
    11'b01100010100: data <= 32'hbd98b41f;
    11'b01100010101: data <= 32'h36debd23;
    11'b01100010110: data <= 32'h4071bd33;
    11'b01100010111: data <= 32'h3f7ebb32;
    11'b01100011000: data <= 32'h3338bb87;
    11'b01100011001: data <= 32'hb7d4baff;
    11'b01100011010: data <= 32'h20933083;
    11'b01100011011: data <= 32'h27d23cdf;
    11'b01100011100: data <= 32'hbc71391f;
    11'b01100011101: data <= 32'hc010bd2e;
    11'b01100011110: data <= 32'hbe45c059;
    11'b01100011111: data <= 32'hb7b6ba31;
    11'b01100100000: data <= 32'h269e3c8d;
    11'b01100100001: data <= 32'h31193d88;
    11'b01100100010: data <= 32'h38f6372a;
    11'b01100100011: data <= 32'h3af0369a;
    11'b01100100100: data <= 32'habb93e4b;
    11'b01100100101: data <= 32'hbda0401d;
    11'b01100100110: data <= 32'hbcec3a9c;
    11'b01100100111: data <= 32'h3965ba4e;
    11'b01100101000: data <= 32'h403fbccb;
    11'b01100101001: data <= 32'h3e43b998;
    11'b01100101010: data <= 32'h34cbb691;
    11'b01100101011: data <= 32'h3608b4aa;
    11'b01100101100: data <= 32'h3d9f34d1;
    11'b01100101101: data <= 32'h3ceb3a7f;
    11'b01100101110: data <= 32'hb8fe2883;
    11'b01100101111: data <= 32'hc041be7a;
    11'b01100110000: data <= 32'hbed8c05c;
    11'b01100110001: data <= 32'hb546bb8c;
    11'b01100110010: data <= 32'h34a93554;
    11'b01100110011: data <= 32'h2d4c2c43;
    11'b01100110100: data <= 32'h1c6db987;
    11'b01100110101: data <= 32'h22372bf1;
    11'b01100110110: data <= 32'hb9463fe7;
    11'b01100110111: data <= 32'hbe5e4145;
    11'b01100111000: data <= 32'hbd783c63;
    11'b01100111001: data <= 32'h2e5aba0a;
    11'b01100111010: data <= 32'h3c5dbba3;
    11'b01100111011: data <= 32'h393a252c;
    11'b01100111100: data <= 32'h311f3859;
    11'b01100111101: data <= 32'h3c5b3654;
    11'b01100111110: data <= 32'h40d037cb;
    11'b01100111111: data <= 32'h3f953a39;
    11'b01101000000: data <= 32'hb6023441;
    11'b01101000001: data <= 32'hbf77bbee;
    11'b01101000010: data <= 32'hbc45be64;
    11'b01101000011: data <= 32'h3864bc24;
    11'b01101000100: data <= 32'h3b35b8dd;
    11'b01101000101: data <= 32'h2f80bce9;
    11'b01101000110: data <= 32'hb505be8a;
    11'b01101000111: data <= 32'hb100b48f;
    11'b01101001000: data <= 32'hb73a3f6d;
    11'b01101001001: data <= 32'hbd574089;
    11'b01101001010: data <= 32'hbe91378f;
    11'b01101001011: data <= 32'hbb81bcae;
    11'b01101001100: data <= 32'hb4d0ba2c;
    11'b01101001101: data <= 32'hb612393c;
    11'b01101001110: data <= 32'hb0a93c66;
    11'b01101001111: data <= 32'h3cf13851;
    11'b01101010000: data <= 32'h40e93726;
    11'b01101010001: data <= 32'h3ea53c6a;
    11'b01101010010: data <= 32'hb8423cf7;
    11'b01101010011: data <= 32'hbdfb34d3;
    11'b01101010100: data <= 32'hb25ab962;
    11'b01101010101: data <= 32'h3d97bb46;
    11'b01101010110: data <= 32'h3d1ebc56;
    11'b01101010111: data <= 32'h305fbef0;
    11'b01101011000: data <= 32'haf4abf53;
    11'b01101011001: data <= 32'h38b2b62b;
    11'b01101011010: data <= 32'h38ba3d92;
    11'b01101011011: data <= 32'hb9363d57;
    11'b01101011100: data <= 32'hbf1fb7db;
    11'b01101011101: data <= 32'hbf01be8b;
    11'b01101011110: data <= 32'hbcd3b9ad;
    11'b01101011111: data <= 32'hbb6e39e9;
    11'b01101100000: data <= 32'hb6be39e4;
    11'b01101100001: data <= 32'h3a74b10d;
    11'b01101100010: data <= 32'h3ea028ae;
    11'b01101100011: data <= 32'h3a663df8;
    11'b01101100100: data <= 32'hbb6640a7;
    11'b01101100101: data <= 32'hbd093dee;
    11'b01101100110: data <= 32'h33c42c8a;
    11'b01101100111: data <= 32'h3df3b8e7;
    11'b01101101000: data <= 32'h3bb0baad;
    11'b01101101001: data <= 32'haa60bced;
    11'b01101101010: data <= 32'h3677bcff;
    11'b01101101011: data <= 32'h3f31b277;
    11'b01101101100: data <= 32'h3f8f3b89;
    11'b01101101101: data <= 32'h2f5d388f;
    11'b01101101110: data <= 32'hbe8bbbea;
    11'b01101101111: data <= 32'hbf4abe9a;
    11'b01101110000: data <= 32'hbc6ab934;
    11'b01101110001: data <= 32'hb9b13443;
    11'b01101110010: data <= 32'hb800b640;
    11'b01101110011: data <= 32'h3120bd94;
    11'b01101110100: data <= 32'h3968b8ed;
    11'b01101110101: data <= 32'h29563e76;
    11'b01101110110: data <= 32'hbc8f41a0;
    11'b01101110111: data <= 32'hbcd03f4c;
    11'b01101111000: data <= 32'ha5b3327b;
    11'b01101111001: data <= 32'h392ab544;
    11'b01101111010: data <= 32'ha95cadb9;
    11'b01101111011: data <= 32'hb803b1ea;
    11'b01101111100: data <= 32'h3a7bb6cb;
    11'b01101111101: data <= 32'h41602799;
    11'b01101111110: data <= 32'h414b3a06;
    11'b01101111111: data <= 32'h381c3821;
    11'b01110000000: data <= 32'hbd28b871;
    11'b01110000001: data <= 32'hbc98bbf2;
    11'b01110000010: data <= 32'hb140b6e7;
    11'b01110000011: data <= 32'h1f1bb59e;
    11'b01110000100: data <= 32'hb69fbe41;
    11'b01110000101: data <= 32'hb46dc0e6;
    11'b01110000110: data <= 32'h3406bca5;
    11'b01110000111: data <= 32'h2abf3d75;
    11'b01110001000: data <= 32'hbaa540cf;
    11'b01110001001: data <= 32'hbcb83cad;
    11'b01110001010: data <= 32'hb9d2b48d;
    11'b01110001011: data <= 32'hb8eab226;
    11'b01110001100: data <= 32'hbcce3915;
    11'b01110001101: data <= 32'hbc3338c6;
    11'b01110001110: data <= 32'h3a3ead58;
    11'b01110001111: data <= 32'h4161a870;
    11'b01110010000: data <= 32'h40d43a75;
    11'b01110010001: data <= 32'h35413ca4;
    11'b01110010010: data <= 32'hbb9338c3;
    11'b01110010011: data <= 32'hb2aa2c34;
    11'b01110010100: data <= 32'h3b0da678;
    11'b01110010101: data <= 32'h38a0b8e4;
    11'b01110010110: data <= 32'hb643c007;
    11'b01110010111: data <= 32'hb511c15c;
    11'b01110011000: data <= 32'h3961bd22;
    11'b01110011001: data <= 32'h3b863b39;
    11'b01110011010: data <= 32'ha4173da5;
    11'b01110011011: data <= 32'hbc0f28c8;
    11'b01110011100: data <= 32'hbd2abb78;
    11'b01110011101: data <= 32'hbdd2b0f8;
    11'b01110011110: data <= 32'hbf4a3b6a;
    11'b01110011111: data <= 32'hbd9d3856;
    11'b01110100000: data <= 32'h3518b8e8;
    11'b01110100001: data <= 32'h3f59b87e;
    11'b01110100010: data <= 32'h3da73b0f;
    11'b01110100011: data <= 32'hb35b3fe1;
    11'b01110100100: data <= 32'hb9ff3ed0;
    11'b01110100101: data <= 32'h368e3b52;
    11'b01110100110: data <= 32'h3d0e3682;
    11'b01110100111: data <= 32'h3709b4a0;
    11'b01110101000: data <= 32'hb960bdda;
    11'b01110101001: data <= 32'haee2bffd;
    11'b01110101010: data <= 32'h3e5cbbb0;
    11'b01110101011: data <= 32'h405037f1;
    11'b01110101100: data <= 32'h3b0e37eb;
    11'b01110101101: data <= 32'hb971b9ea;
    11'b01110101110: data <= 32'hbcfebc8f;
    11'b01110101111: data <= 32'hbd3da716;
    11'b01110110000: data <= 32'hbe2d39fe;
    11'b01110110001: data <= 32'hbd88b489;
    11'b01110110010: data <= 32'hb49bbf08;
    11'b01110110011: data <= 32'h39d1bd71;
    11'b01110110100: data <= 32'h364b3a2b;
    11'b01110110101: data <= 32'hb92f409a;
    11'b01110110110: data <= 32'hb93b4002;
    11'b01110110111: data <= 32'h36bd3c20;
    11'b01110111000: data <= 32'h39d33920;
    11'b01110111001: data <= 32'hb75636e8;
    11'b01110111010: data <= 32'hbd1cb4e7;
    11'b01110111011: data <= 32'h2828bb73;
    11'b01110111100: data <= 32'h4097b82a;
    11'b01110111101: data <= 32'h41c034bb;
    11'b01110111110: data <= 32'h3d3d31f4;
    11'b01110111111: data <= 32'hb538b8eb;
    11'b01111000000: data <= 32'hb894b8d6;
    11'b01111000001: data <= 32'hb46e3572;
    11'b01111000010: data <= 32'hb8eb36b1;
    11'b01111000011: data <= 32'hbc5fbcfa;
    11'b01111000100: data <= 32'hb9b5c18d;
    11'b01111000101: data <= 32'h2c8abfea;
    11'b01111000110: data <= 32'h2de3374d;
    11'b01111000111: data <= 32'hb7c03f71;
    11'b01111001000: data <= 32'hb7ef3d14;
    11'b01111001001: data <= 32'h22d935e8;
    11'b01111001010: data <= 32'hb4c838bf;
    11'b01111001011: data <= 32'hbe543c87;
    11'b01111001100: data <= 32'hbfbe3978;
    11'b01111001101: data <= 32'haf67b474;
    11'b01111001110: data <= 32'h4076b6a1;
    11'b01111001111: data <= 32'h412733aa;
    11'b01111010000: data <= 32'h3bef383e;
    11'b01111010001: data <= 32'hb05e3485;
    11'b01111010010: data <= 32'h3578369e;
    11'b01111010011: data <= 32'h3ba63b17;
    11'b01111010100: data <= 32'h34323533;
    11'b01111010101: data <= 32'hbb05be68;
    11'b01111010110: data <= 32'hbaaec1ea;
    11'b01111010111: data <= 32'h325ac008;
    11'b01111011000: data <= 32'h39ab2ec1;
    11'b01111011001: data <= 32'h346c3b17;
    11'b01111011010: data <= 32'hb180a811;
    11'b01111011011: data <= 32'hb575b895;
    11'b01111011100: data <= 32'hbc1536c7;
    11'b01111011101: data <= 32'hc0583de8;
    11'b01111011110: data <= 32'hc0833b4a;
    11'b01111011111: data <= 32'hb81db829;
    11'b01111100000: data <= 32'h3d8abaec;
    11'b01111100001: data <= 32'h3db230da;
    11'b01111100010: data <= 32'h31153c66;
    11'b01111100011: data <= 32'hb0d23cfc;
    11'b01111100100: data <= 32'h3bef3cfd;
    11'b01111100101: data <= 32'h3e703d5b;
    11'b01111100110: data <= 32'h36d13918;
    11'b01111100111: data <= 32'hbc39bc2a;
    11'b01111101000: data <= 32'hba3ec049;
    11'b01111101001: data <= 32'h3ad5bdc9;
    11'b01111101010: data <= 32'h3f06ae20;
    11'b01111101011: data <= 32'h3cabaa09;
    11'b01111101100: data <= 32'h336bbc45;
    11'b01111101101: data <= 32'hb410bc61;
    11'b01111101110: data <= 32'hbac636b8;
    11'b01111101111: data <= 32'hbf283dc0;
    11'b01111110000: data <= 32'hc00e35c2;
    11'b01111110001: data <= 32'hbb76bde3;
    11'b01111110010: data <= 32'h3445bea2;
    11'b01111110011: data <= 32'h30feac5c;
    11'b01111110100: data <= 32'hb8ad3d58;
    11'b01111110101: data <= 32'hb2d63e00;
    11'b01111110110: data <= 32'h3c7d3d26;
    11'b01111110111: data <= 32'h3d6b3daa;
    11'b01111111000: data <= 32'hb41a3ccd;
    11'b01111111001: data <= 32'hbe952fa3;
    11'b01111111010: data <= 32'hba34bac1;
    11'b01111111011: data <= 32'h3daeb969;
    11'b01111111100: data <= 32'h40d0af3e;
    11'b01111111101: data <= 32'h3e30b749;
    11'b01111111110: data <= 32'h37c2bced;
    11'b01111111111: data <= 32'h34e0ba68;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    