
module memory_rom_4(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'hbc8fbc6d;
    11'b00000000001: data <= 32'hb8d8b85f;
    11'b00000000010: data <= 32'h396b3a16;
    11'b00000000011: data <= 32'h38253f36;
    11'b00000000100: data <= 32'hbcd33d04;
    11'b00000000101: data <= 32'hc0bab2f7;
    11'b00000000110: data <= 32'hbeafb8ad;
    11'b00000000111: data <= 32'hb3283847;
    11'b00000001000: data <= 32'h38803cf1;
    11'b00000001001: data <= 32'h3aff351c;
    11'b00000001010: data <= 32'h3d9bb9c3;
    11'b00000001011: data <= 32'h3e8d2623;
    11'b00000001100: data <= 32'h3a4f3f27;
    11'b00000001101: data <= 32'hb651402e;
    11'b00000001110: data <= 32'hb66134ca;
    11'b00000001111: data <= 32'h38efbe55;
    11'b00000010000: data <= 32'h3b28bf8f;
    11'b00000010001: data <= 32'haed6bd11;
    11'b00000010010: data <= 32'hb97fbc06;
    11'b00000010011: data <= 32'h363fbb6a;
    11'b00000010100: data <= 32'h3e98b359;
    11'b00000010101: data <= 32'h3b0238ee;
    11'b00000010110: data <= 32'hbe0037e6;
    11'b00000010111: data <= 32'hc1b1b509;
    11'b00000011000: data <= 32'hbfd2b66f;
    11'b00000011001: data <= 32'hb68c3631;
    11'b00000011010: data <= 32'h2b0f3894;
    11'b00000011011: data <= 32'hb094b679;
    11'b00000011100: data <= 32'h3307baf9;
    11'b00000011101: data <= 32'h3b3138d9;
    11'b00000011110: data <= 32'h3a4c4153;
    11'b00000011111: data <= 32'h27db4176;
    11'b00000100000: data <= 32'hb11a393d;
    11'b00000100001: data <= 32'h35e4bc7b;
    11'b00000100010: data <= 32'h37a8bc21;
    11'b00000100011: data <= 32'hacb9b42c;
    11'b00000100100: data <= 32'h2beab70d;
    11'b00000100101: data <= 32'h3dfabc96;
    11'b00000100110: data <= 32'h4103bbc5;
    11'b00000100111: data <= 32'h3d13a475;
    11'b00000101000: data <= 32'hbcfa35bc;
    11'b00000101001: data <= 32'hc0acb12a;
    11'b00000101010: data <= 32'hbd1cb847;
    11'b00000101011: data <= 32'hae6db5eb;
    11'b00000101100: data <= 32'hb699b865;
    11'b00000101101: data <= 32'hbcc1bd25;
    11'b00000101110: data <= 32'hba01bcb0;
    11'b00000101111: data <= 32'h37d63948;
    11'b00000110000: data <= 32'h3a88413a;
    11'b00000110001: data <= 32'hab3d40f5;
    11'b00000110010: data <= 32'hba1838f9;
    11'b00000110011: data <= 32'hb8a6b7ab;
    11'b00000110100: data <= 32'hb3fd323d;
    11'b00000110101: data <= 32'hb1993b54;
    11'b00000110110: data <= 32'h37412e64;
    11'b00000110111: data <= 32'h3f9dbce1;
    11'b00000111000: data <= 32'h415bbc69;
    11'b00000111001: data <= 32'h3de1347f;
    11'b00000111010: data <= 32'hb87c3c0d;
    11'b00000111011: data <= 32'hbc80350b;
    11'b00000111100: data <= 32'had7db96e;
    11'b00000111101: data <= 32'h36c1bc3e;
    11'b00000111110: data <= 32'hb947bd42;
    11'b00000111111: data <= 32'hbeaebf14;
    11'b00001000000: data <= 32'hbaedbdfd;
    11'b00001000001: data <= 32'h3a632cff;
    11'b00001000010: data <= 32'h3c353e7a;
    11'b00001000011: data <= 32'hb6403ded;
    11'b00001000100: data <= 32'hbe9b341d;
    11'b00001000101: data <= 32'hbe331a37;
    11'b00001000110: data <= 32'hbaeb3c3c;
    11'b00001000111: data <= 32'hb76a3de3;
    11'b00001001000: data <= 32'h2f1f2fec;
    11'b00001001001: data <= 32'h3d18bd38;
    11'b00001001010: data <= 32'h400db9d4;
    11'b00001001011: data <= 32'h3d723cce;
    11'b00001001100: data <= 32'h30e44008;
    11'b00001001101: data <= 32'h29823b21;
    11'b00001001110: data <= 32'h3a97b8ac;
    11'b00001001111: data <= 32'h3990bc4b;
    11'b00001010000: data <= 32'hb9bcbc79;
    11'b00001010001: data <= 32'hbdc7be08;
    11'b00001010010: data <= 32'hafc6bea0;
    11'b00001010011: data <= 32'h3eafba6d;
    11'b00001010100: data <= 32'h3de634bb;
    11'b00001010101: data <= 32'hb8963661;
    11'b00001010110: data <= 32'hc024af67;
    11'b00001010111: data <= 32'hbf243123;
    11'b00001011000: data <= 32'hbb7b3c89;
    11'b00001011001: data <= 32'hba5e3c53;
    11'b00001011010: data <= 32'hba7eb7b0;
    11'b00001011011: data <= 32'ha82ebe1d;
    11'b00001011100: data <= 32'h3bcab4b5;
    11'b00001011101: data <= 32'h3c463fe8;
    11'b00001011110: data <= 32'h3838413a;
    11'b00001011111: data <= 32'h37f83cb6;
    11'b00001100000: data <= 32'h3af4b3c0;
    11'b00001100001: data <= 32'h36d4b4a0;
    11'b00001100010: data <= 32'hba0a9590;
    11'b00001100011: data <= 32'hbaf7b92f;
    11'b00001100100: data <= 32'h3ad6be54;
    11'b00001100101: data <= 32'h40fabde4;
    11'b00001100110: data <= 32'h3f5fb85d;
    11'b00001100111: data <= 32'hb625aabf;
    11'b00001101000: data <= 32'hbe6db091;
    11'b00001101001: data <= 32'hbc0b2d90;
    11'b00001101010: data <= 32'hb5c83895;
    11'b00001101011: data <= 32'hbbd82f6a;
    11'b00001101100: data <= 32'hbf17bd4a;
    11'b00001101101: data <= 32'hbccdbf60;
    11'b00001101110: data <= 32'h3361b33c;
    11'b00001101111: data <= 32'h3b0d3fca;
    11'b00001110000: data <= 32'h37a9408f;
    11'b00001110001: data <= 32'h2ecb3b56;
    11'b00001110010: data <= 32'h2ed73083;
    11'b00001110011: data <= 32'hb40d3ad3;
    11'b00001110100: data <= 32'hbb363d75;
    11'b00001110101: data <= 32'hb81b3390;
    11'b00001110110: data <= 32'h3d08bda1;
    11'b00001110111: data <= 32'h4132be79;
    11'b00001111000: data <= 32'h3f71b776;
    11'b00001111001: data <= 32'h2ce4361e;
    11'b00001111010: data <= 32'hb7953444;
    11'b00001111011: data <= 32'h35c4202a;
    11'b00001111100: data <= 32'h380ea934;
    11'b00001111101: data <= 32'hbba8b8f5;
    11'b00001111110: data <= 32'hc07ebf0d;
    11'b00001111111: data <= 32'hbe29c012;
    11'b00010000000: data <= 32'h3495b902;
    11'b00010000001: data <= 32'h3c153c17;
    11'b00010000010: data <= 32'h32f03c77;
    11'b00010000011: data <= 32'hb95a32d3;
    11'b00010000100: data <= 32'hba703570;
    11'b00010000101: data <= 32'hbabd3ec4;
    11'b00010000110: data <= 32'hbc6e404c;
    11'b00010000111: data <= 32'hb9c1385b;
    11'b00010001000: data <= 32'h3980bd72;
    11'b00010001001: data <= 32'h3f31bd3f;
    11'b00010001010: data <= 32'h3db934f6;
    11'b00010001011: data <= 32'h380a3d32;
    11'b00010001100: data <= 32'h39423a99;
    11'b00010001101: data <= 32'h3e032c5d;
    11'b00010001110: data <= 32'h3c61b07f;
    11'b00010001111: data <= 32'hbac9b787;
    11'b00010010000: data <= 32'hc027bd84;
    11'b00010010001: data <= 32'hbbb3bf9e;
    11'b00010010010: data <= 32'h3c2bbced;
    11'b00010010011: data <= 32'h3db2b41a;
    11'b00010010100: data <= 32'h28c6b27b;
    11'b00010010101: data <= 32'hbc84b800;
    11'b00010010110: data <= 32'hbc4b34c0;
    11'b00010010111: data <= 32'hba903f3e;
    11'b00010011000: data <= 32'hbcc73fc8;
    11'b00010011001: data <= 32'hbd8d2dd6;
    11'b00010011010: data <= 32'hb88fbe38;
    11'b00010011011: data <= 32'h381cbb42;
    11'b00010011100: data <= 32'h3a3b3c57;
    11'b00010011101: data <= 32'h392f3fa9;
    11'b00010011110: data <= 32'h3c933c30;
    11'b00010011111: data <= 32'h3f0932d4;
    11'b00010100000: data <= 32'h3c1036bf;
    11'b00010100001: data <= 32'hbaae38c5;
    11'b00010100010: data <= 32'hbe33b4cf;
    11'b00010100011: data <= 32'ha5cebddd;
    11'b00010100100: data <= 32'h3f71be97;
    11'b00010100101: data <= 32'h3f02bc78;
    11'b00010100110: data <= 32'h2d12bb16;
    11'b00010100111: data <= 32'hbaceba16;
    11'b00010101000: data <= 32'hb593309a;
    11'b00010101001: data <= 32'haa1b3d39;
    11'b00010101010: data <= 32'hbc193c33;
    11'b00010101011: data <= 32'hc02bb9dc;
    11'b00010101100: data <= 32'hbefdbf65;
    11'b00010101101: data <= 32'hb7aab9e7;
    11'b00010101110: data <= 32'h350a3cd1;
    11'b00010101111: data <= 32'h37c23e85;
    11'b00010110000: data <= 32'h3a7e38e9;
    11'b00010110001: data <= 32'h3c66343f;
    11'b00010110010: data <= 32'h36183d32;
    11'b00010110011: data <= 32'hbbc63fda;
    11'b00010110100: data <= 32'hbc873ac3;
    11'b00010110101: data <= 32'h37eabbcf;
    11'b00010110110: data <= 32'h4009be90;
    11'b00010110111: data <= 32'h3e83bc63;
    11'b00010111000: data <= 32'h33bcb8b8;
    11'b00010111001: data <= 32'h2736b6e9;
    11'b00010111010: data <= 32'h3c132b18;
    11'b00010111011: data <= 32'h3c593956;
    11'b00010111100: data <= 32'hb9433386;
    11'b00010111101: data <= 32'hc0bfbce2;
    11'b00010111110: data <= 32'hc048bfbc;
    11'b00010111111: data <= 32'hb8c7bb08;
    11'b00011000000: data <= 32'h35453823;
    11'b00011000001: data <= 32'h326c3796;
    11'b00011000010: data <= 32'h290ab5a5;
    11'b00011000011: data <= 32'h309c2ebc;
    11'b00011000100: data <= 32'hb40c3fb7;
    11'b00011000101: data <= 32'hbc6e4199;
    11'b00011000110: data <= 32'hbc7e3d71;
    11'b00011000111: data <= 32'h3089ba0f;
    11'b00011001000: data <= 32'h3cf1bd28;
    11'b00011001001: data <= 32'h3b97b579;
    11'b00011001010: data <= 32'h34e9355a;
    11'b00011001011: data <= 32'h3b7d3119;
    11'b00011001100: data <= 32'h406c2cba;
    11'b00011001101: data <= 32'h3fa6365c;
    11'b00011001110: data <= 32'hb541320b;
    11'b00011001111: data <= 32'hc042baef;
    11'b00011010000: data <= 32'hbe64be4f;
    11'b00011010001: data <= 32'h3017bc85;
    11'b00011010010: data <= 32'h39f4b83e;
    11'b00011010011: data <= 32'h95d2bb28;
    11'b00011010100: data <= 32'hb862bd53;
    11'b00011010101: data <= 32'hb4bab27a;
    11'b00011010110: data <= 32'hb4633fc8;
    11'b00011010111: data <= 32'hbc014148;
    11'b00011011000: data <= 32'hbdd43bd2;
    11'b00011011001: data <= 32'hbb0dbb72;
    11'b00011011010: data <= 32'hae1abaf3;
    11'b00011011011: data <= 32'h22493833;
    11'b00011011100: data <= 32'h30b13c60;
    11'b00011011101: data <= 32'h3d2c36fa;
    11'b00011011110: data <= 32'h410c2c2b;
    11'b00011011111: data <= 32'h3fc9393f;
    11'b00011100000: data <= 32'hb41c3c18;
    11'b00011100001: data <= 32'hbe5533f8;
    11'b00011100010: data <= 32'hb8c3bac5;
    11'b00011100011: data <= 32'h3c40bcd9;
    11'b00011100100: data <= 32'h3c88bcf4;
    11'b00011100101: data <= 32'hace0be97;
    11'b00011100110: data <= 32'hb84dbf01;
    11'b00011100111: data <= 32'h3296b75a;
    11'b00011101000: data <= 32'h382a3da4;
    11'b00011101001: data <= 32'hb85d3ed6;
    11'b00011101010: data <= 32'hbf372c49;
    11'b00011101011: data <= 32'hbf8bbd23;
    11'b00011101100: data <= 32'hbcacb8ea;
    11'b00011101101: data <= 32'hb9423b01;
    11'b00011101110: data <= 32'hb1753c17;
    11'b00011101111: data <= 32'h3b5396fd;
    11'b00011110000: data <= 32'h3f6bb0c7;
    11'b00011110001: data <= 32'h3d0a3cba;
    11'b00011110010: data <= 32'hb71b4068;
    11'b00011110011: data <= 32'hbc6c3dec;
    11'b00011110100: data <= 32'h2fb9af0f;
    11'b00011110101: data <= 32'h3db3bc01;
    11'b00011110110: data <= 32'h3c18bc9b;
    11'b00011110111: data <= 32'hb0e4bd77;
    11'b00011111000: data <= 32'h9318bda8;
    11'b00011111001: data <= 32'h3d83b824;
    11'b00011111010: data <= 32'h3ef839d6;
    11'b00011111011: data <= 32'h2e3339cf;
    11'b00011111100: data <= 32'hbf5fb8ec;
    11'b00011111101: data <= 32'hc063bd9f;
    11'b00011111110: data <= 32'hbd4db863;
    11'b00011111111: data <= 32'hb97d381e;
    11'b00100000000: data <= 32'hb7532c46;
    11'b00100000001: data <= 32'h2f03bc33;
    11'b00100000010: data <= 32'h3a1ab8d2;
    11'b00100000011: data <= 32'h37293e1c;
    11'b00100000100: data <= 32'hb91341de;
    11'b00100000101: data <= 32'hbb65401d;
    11'b00100000110: data <= 32'h2cbc3298;
    11'b00100000111: data <= 32'h3ac5b8d4;
    11'b00100001000: data <= 32'h3461b5d0;
    11'b00100001001: data <= 32'hb630b565;
    11'b00100001010: data <= 32'h38ccb958;
    11'b00100001011: data <= 32'h40e7b6e9;
    11'b00100001100: data <= 32'h414d3527;
    11'b00100001101: data <= 32'h389c3656;
    11'b00100001110: data <= 32'hbe06b78e;
    11'b00100001111: data <= 32'hbe6fbbfc;
    11'b00100010000: data <= 32'hb838b80c;
    11'b00100010001: data <= 32'hb0c4b2ca;
    11'b00100010010: data <= 32'hb8bdbcb0;
    11'b00100010011: data <= 32'hb8b0c043;
    11'b00100010100: data <= 32'h2c13bc6f;
    11'b00100010101: data <= 32'h32af3d9e;
    11'b00100010110: data <= 32'hb8094174;
    11'b00100010111: data <= 32'hbbdc3e8a;
    11'b00100011000: data <= 32'hb8f9aa2b;
    11'b00100011001: data <= 32'hb580b39a;
    11'b00100011010: data <= 32'hba3b38b8;
    11'b00100011011: data <= 32'hba4d393f;
    11'b00100011100: data <= 32'h3a34b17e;
    11'b00100011101: data <= 32'h416ab6f6;
    11'b00100011110: data <= 32'h415c3549;
    11'b00100011111: data <= 32'h38ec3b3c;
    11'b00100100000: data <= 32'hbbed37d3;
    11'b00100100001: data <= 32'hb844b0b8;
    11'b00100100010: data <= 32'h38ebb50c;
    11'b00100100011: data <= 32'h3744b99b;
    11'b00100100100: data <= 32'hb916bf72;
    11'b00100100101: data <= 32'hba5cc12a;
    11'b00100100110: data <= 32'h33d3bd8d;
    11'b00100100111: data <= 32'h3aab3af3;
    11'b00100101000: data <= 32'h2bd03eea;
    11'b00100101001: data <= 32'hbc25385b;
    11'b00100101010: data <= 32'hbd80b8d5;
    11'b00100101011: data <= 32'hbd62a815;
    11'b00100101100: data <= 32'hbe123c86;
    11'b00100101101: data <= 32'hbcbd3b29;
    11'b00100101110: data <= 32'h35c3b6c2;
    11'b00100101111: data <= 32'h3fe9b9ec;
    11'b00100110000: data <= 32'h3f61387a;
    11'b00100110001: data <= 32'h33e63f3e;
    11'b00100110010: data <= 32'hb8903e92;
    11'b00100110011: data <= 32'h35943983;
    11'b00100110100: data <= 32'h3d1a2839;
    11'b00100110101: data <= 32'h3862b84c;
    11'b00100110110: data <= 32'hba3abe1b;
    11'b00100110111: data <= 32'hb860c046;
    11'b00100111000: data <= 32'h3c83bd30;
    11'b00100111001: data <= 32'h3fdc33d2;
    11'b00100111010: data <= 32'h3a9c38ce;
    11'b00100111011: data <= 32'hbb1ab6d1;
    11'b00100111100: data <= 32'hbe42bb8b;
    11'b00100111101: data <= 32'hbdd22c9b;
    11'b00100111110: data <= 32'hbdee3c2e;
    11'b00100111111: data <= 32'hbd78339a;
    11'b00101000000: data <= 32'hb666bd78;
    11'b00101000001: data <= 32'h3a12bd4f;
    11'b00101000010: data <= 32'h3a13396e;
    11'b00101000011: data <= 32'hb18040c6;
    11'b00101000100: data <= 32'hb60e405a;
    11'b00101000101: data <= 32'h387b3be9;
    11'b00101000110: data <= 32'h3c043616;
    11'b00101000111: data <= 32'had31333f;
    11'b00101001000: data <= 32'hbc95b634;
    11'b00101001001: data <= 32'hb26abc90;
    11'b00101001010: data <= 32'h4009bbd8;
    11'b00101001011: data <= 32'h41aab0c6;
    11'b00101001100: data <= 32'h3d5727bc;
    11'b00101001101: data <= 32'hb858b8c9;
    11'b00101001110: data <= 32'hbbd2b96f;
    11'b00101001111: data <= 32'hb88133a8;
    11'b00101010000: data <= 32'hb9d038b7;
    11'b00101010001: data <= 32'hbd21ba5a;
    11'b00101010010: data <= 32'hbc41c0d2;
    11'b00101010011: data <= 32'hb12cbf9d;
    11'b00101010100: data <= 32'h326037da;
    11'b00101010101: data <= 32'hb2d0404a;
    11'b00101010110: data <= 32'hb5493eb0;
    11'b00101010111: data <= 32'h30a03871;
    11'b00101011000: data <= 32'h29a8386a;
    11'b00101011001: data <= 32'hbc5f3c91;
    11'b00101011010: data <= 32'hbe9b3a76;
    11'b00101011011: data <= 32'hb081b523;
    11'b00101011100: data <= 32'h406bba49;
    11'b00101011101: data <= 32'h4198b315;
    11'b00101011110: data <= 32'h3cf5341c;
    11'b00101011111: data <= 32'hb1eb2f1f;
    11'b00101100000: data <= 32'h2c0d2fb2;
    11'b00101100001: data <= 32'h3a1d3878;
    11'b00101100010: data <= 32'h3236342e;
    11'b00101100011: data <= 32'hbc6dbd93;
    11'b00101100100: data <= 32'hbd4dc1a1;
    11'b00101100101: data <= 32'hb420c032;
    11'b00101100110: data <= 32'h38652c66;
    11'b00101100111: data <= 32'h34833cae;
    11'b00101101000: data <= 32'hb3c9369a;
    11'b00101101001: data <= 32'hb694b4df;
    11'b00101101010: data <= 32'hbac13839;
    11'b00101101011: data <= 32'hbf363ed8;
    11'b00101101100: data <= 32'hc0093d44;
    11'b00101101101: data <= 32'hb7dfb46d;
    11'b00101101110: data <= 32'h3df5bbf1;
    11'b00101101111: data <= 32'h3f3fb034;
    11'b00101110000: data <= 32'h38b63b7e;
    11'b00101110001: data <= 32'h1db13c7f;
    11'b00101110010: data <= 32'h3ba83b89;
    11'b00101110011: data <= 32'h3ec03b6e;
    11'b00101110100: data <= 32'h38d0369f;
    11'b00101110101: data <= 32'hbc7bbc36;
    11'b00101110110: data <= 32'hbcd2c07c;
    11'b00101110111: data <= 32'h3613bf08;
    11'b00101111000: data <= 32'h3e0fb567;
    11'b00101111001: data <= 32'h3c26292b;
    11'b00101111010: data <= 32'ha74bba80;
    11'b00101111011: data <= 32'hb87bbbc7;
    11'b00101111100: data <= 32'hbb723790;
    11'b00101111101: data <= 32'hbead3ef1;
    11'b00101111110: data <= 32'hbffa3b57;
    11'b00101111111: data <= 32'hbc3abc1e;
    11'b00110000000: data <= 32'h3460be42;
    11'b00110000001: data <= 32'h37afaf20;
    11'b00110000010: data <= 32'hb16c3db3;
    11'b00110000011: data <= 32'h21f13e78;
    11'b00110000100: data <= 32'h3d0c3cb2;
    11'b00110000101: data <= 32'h3ebd3c7e;
    11'b00110000110: data <= 32'h32283c10;
    11'b00110000111: data <= 32'hbdd62d3f;
    11'b00110001000: data <= 32'hbbd2bc0e;
    11'b00110001001: data <= 32'h3c92bc66;
    11'b00110001010: data <= 32'h40a6b830;
    11'b00110001011: data <= 32'h3e05b8d9;
    11'b00110001100: data <= 32'h3307bd0d;
    11'b00110001101: data <= 32'haddcbbad;
    11'b00110001110: data <= 32'ha92838b7;
    11'b00110001111: data <= 32'hb9a33da3;
    11'b00110010000: data <= 32'hbe5129b9;
    11'b00110010001: data <= 32'hbe01bffa;
    11'b00110010010: data <= 32'hb9a8c03e;
    11'b00110010011: data <= 32'hb5e1b41a;
    11'b00110010100: data <= 32'hb7e93d07;
    11'b00110010101: data <= 32'ha4f43c71;
    11'b00110010110: data <= 32'h3bd2387a;
    11'b00110010111: data <= 32'h3b4a3bee;
    11'b00110011000: data <= 32'hb9c53ed9;
    11'b00110011001: data <= 32'hbfd93d4d;
    11'b00110011010: data <= 32'hbb612e36;
    11'b00110011011: data <= 32'h3d76b8b8;
    11'b00110011100: data <= 32'h408fb7bc;
    11'b00110011101: data <= 32'h3d0bb80f;
    11'b00110011110: data <= 32'h34ffba25;
    11'b00110011111: data <= 32'h39f4b48a;
    11'b00110100000: data <= 32'h3d4e3b50;
    11'b00110100001: data <= 32'h380c3c80;
    11'b00110100010: data <= 32'hbc43b85e;
    11'b00110100011: data <= 32'hbe79c0c6;
    11'b00110100100: data <= 32'hbb62c068;
    11'b00110100101: data <= 32'hb41fb757;
    11'b00110100110: data <= 32'hb105376f;
    11'b00110100111: data <= 32'h2c65b1de;
    11'b00110101000: data <= 32'h37fab8a8;
    11'b00110101001: data <= 32'h2c6138f0;
    11'b00110101010: data <= 32'hbda94038;
    11'b00110101011: data <= 32'hc0813fc6;
    11'b00110101100: data <= 32'hbc6b367e;
    11'b00110101101: data <= 32'h3a65b8cd;
    11'b00110101110: data <= 32'h3d0eb60c;
    11'b00110101111: data <= 32'h35842ca7;
    11'b00110110000: data <= 32'h30ec313b;
    11'b00110110001: data <= 32'h3dce381b;
    11'b00110110010: data <= 32'h40b33cf9;
    11'b00110110011: data <= 32'h3ccb3ca4;
    11'b00110110100: data <= 32'hbabbb547;
    11'b00110110101: data <= 32'hbdd3bf2a;
    11'b00110110110: data <= 32'hb65dbe7c;
    11'b00110110111: data <= 32'h38b9b83b;
    11'b00110111000: data <= 32'h3876b791;
    11'b00110111001: data <= 32'h3454be05;
    11'b00110111010: data <= 32'h3489be36;
    11'b00110111011: data <= 32'haf1c3496;
    11'b00110111100: data <= 32'hbd134021;
    11'b00110111101: data <= 32'hc00b3ea7;
    11'b00110111110: data <= 32'hbd6eb241;
    11'b00110111111: data <= 32'hb33abc6d;
    11'b00111000000: data <= 32'hb119b5c5;
    11'b00111000001: data <= 32'hb9d738a8;
    11'b00111000010: data <= 32'hb0bf39bb;
    11'b00111000011: data <= 32'h3ea239ef;
    11'b00111000100: data <= 32'h40f13d16;
    11'b00111000101: data <= 32'h3bcd3df3;
    11'b00111000110: data <= 32'hbc5538fa;
    11'b00111000111: data <= 32'hbcf0b7a8;
    11'b00111001000: data <= 32'h359ab924;
    11'b00111001001: data <= 32'h3db5b61b;
    11'b00111001010: data <= 32'h3c1dbbfd;
    11'b00111001011: data <= 32'h3656c02b;
    11'b00111001100: data <= 32'h382bbf0c;
    11'b00111001101: data <= 32'h38e2344d;
    11'b00111001110: data <= 32'hb3673ef3;
    11'b00111001111: data <= 32'hbd2b3aab;
    11'b00111010000: data <= 32'hbdd1bc9f;
    11'b00111010001: data <= 32'hbc44beac;
    11'b00111010010: data <= 32'hbc90b6c4;
    11'b00111010011: data <= 32'hbd4138c7;
    11'b00111010100: data <= 32'hb5b235c0;
    11'b00111010101: data <= 32'h3d702c89;
    11'b00111010110: data <= 32'h3f0e3ac7;
    11'b00111010111: data <= 32'h2e573f58;
    11'b00111011000: data <= 32'hbe563ed9;
    11'b00111011001: data <= 32'hbc833a28;
    11'b00111011010: data <= 32'h39b03125;
    11'b00111011011: data <= 32'h3e0cafac;
    11'b00111011100: data <= 32'h39f7baef;
    11'b00111011101: data <= 32'h334cbeb5;
    11'b00111011110: data <= 32'h3c19bca4;
    11'b00111011111: data <= 32'h3f45389f;
    11'b00111100000: data <= 32'h3c763db6;
    11'b00111100001: data <= 32'hb758309e;
    11'b00111100010: data <= 32'hbd3abea2;
    11'b00111100011: data <= 32'hbce9beeb;
    11'b00111100100: data <= 32'hbc8fb670;
    11'b00111100101: data <= 32'hbc602f2c;
    11'b00111100110: data <= 32'hb4eeba34;
    11'b00111100111: data <= 32'h3af6bcce;
    11'b00111101000: data <= 32'h3ae0306e;
    11'b00111101001: data <= 32'hb97d3fc0;
    11'b00111101010: data <= 32'hbf7d4082;
    11'b00111101011: data <= 32'hbc843cd2;
    11'b00111101100: data <= 32'h36bd350d;
    11'b00111101101: data <= 32'h39372be2;
    11'b00111101110: data <= 32'hb4abb482;
    11'b00111101111: data <= 32'hb447b9be;
    11'b00111110000: data <= 32'h3da7b4b7;
    11'b00111110001: data <= 32'h417f3b5a;
    11'b00111110010: data <= 32'h3fcd3d4a;
    11'b00111110011: data <= 32'ha5a62f92;
    11'b00111110100: data <= 32'hbc1bbcdb;
    11'b00111110101: data <= 32'hb98dbc2a;
    11'b00111110110: data <= 32'hb4c1b0a4;
    11'b00111110111: data <= 32'hb576b7f8;
    11'b00111111000: data <= 32'had9fbff9;
    11'b00111111001: data <= 32'h386dc0a8;
    11'b00111111010: data <= 32'h3790b72d;
    11'b00111111011: data <= 32'hb9813ee9;
    11'b00111111100: data <= 32'hbe3c3fd2;
    11'b00111111101: data <= 32'hbc4c3920;
    11'b00111111110: data <= 32'hb472b21b;
    11'b00111111111: data <= 32'hb94a2c3e;
    11'b01000000000: data <= 32'hbe2334c4;
    11'b01000000001: data <= 32'hbae81ec5;
    11'b01000000010: data <= 32'h3da82cfc;
    11'b01000000011: data <= 32'h41ae3b27;
    11'b01000000100: data <= 32'h3f2d3d7e;
    11'b01000000101: data <= 32'hb3053a05;
    11'b01000000110: data <= 32'hba63a4a8;
    11'b01000000111: data <= 32'h2e8d2f09;
    11'b01000001000: data <= 32'h39683533;
    11'b01000001001: data <= 32'h343dba43;
    11'b01000001010: data <= 32'h2284c111;
    11'b01000001011: data <= 32'h386cc145;
    11'b01000001100: data <= 32'h3b24b87a;
    11'b01000001101: data <= 32'h332e3d77;
    11'b01000001110: data <= 32'hb94e3c5c;
    11'b01000001111: data <= 32'hbaa7b6c3;
    11'b01000010000: data <= 32'hbacbbafc;
    11'b01000010001: data <= 32'hbe631e9a;
    11'b01000010010: data <= 32'hc07e3815;
    11'b01000010011: data <= 32'hbcdeac81;
    11'b01000010100: data <= 32'h3c31b75a;
    11'b01000010101: data <= 32'h4035351b;
    11'b01000010110: data <= 32'h3ac73d83;
    11'b01000010111: data <= 32'hba8d3e36;
    11'b01000011000: data <= 32'hb9a13cb5;
    11'b01000011001: data <= 32'h38ff3c4a;
    11'b01000011010: data <= 32'h3c113a4a;
    11'b01000011011: data <= 32'h2feeb85d;
    11'b01000011100: data <= 32'hb47cc034;
    11'b01000011101: data <= 32'h39ccbfff;
    11'b01000011110: data <= 32'h3f33b1d0;
    11'b01000011111: data <= 32'h3e0a3c49;
    11'b01000100000: data <= 32'h35a6344f;
    11'b01000100001: data <= 32'hb6f6bca1;
    11'b01000100010: data <= 32'hbaecbc54;
    11'b01000100011: data <= 32'hbe4c2fdb;
    11'b01000100100: data <= 32'hc0113559;
    11'b01000100101: data <= 32'hbc8ebb3a;
    11'b01000100110: data <= 32'h388abea5;
    11'b01000100111: data <= 32'h3c5eb8ac;
    11'b01000101000: data <= 32'hb0af3cc3;
    11'b01000101001: data <= 32'hbd0a3fa7;
    11'b01000101010: data <= 32'hb91a3e61;
    11'b01000101011: data <= 32'h38ee3d1d;
    11'b01000101100: data <= 32'h37423be6;
    11'b01000101101: data <= 32'hbaa929ec;
    11'b01000101110: data <= 32'hbbc6bc3b;
    11'b01000101111: data <= 32'h3a63bb9c;
    11'b01000110000: data <= 32'h41093502;
    11'b01000110001: data <= 32'h40a83b6c;
    11'b01000110010: data <= 32'h3b13a0dd;
    11'b01000110011: data <= 32'hacfabc04;
    11'b01000110100: data <= 32'hb4cbb7d4;
    11'b01000110101: data <= 32'hb9533889;
    11'b01000110110: data <= 32'hbc872ab8;
    11'b01000110111: data <= 32'hba31bf8c;
    11'b01000111000: data <= 32'h338bc18b;
    11'b01000111001: data <= 32'h37b5bd39;
    11'b01000111010: data <= 32'hb6f03ac7;
    11'b01000111011: data <= 32'hbc3d3e34;
    11'b01000111100: data <= 32'hb6a23bd5;
    11'b01000111101: data <= 32'h33f0394d;
    11'b01000111110: data <= 32'hb8e03af4;
    11'b01000111111: data <= 32'hc01e3903;
    11'b01001000000: data <= 32'hbef1b069;
    11'b01001000001: data <= 32'h38e9b4d3;
    11'b01001000010: data <= 32'h410736be;
    11'b01001000011: data <= 32'h40453aae;
    11'b01001000100: data <= 32'h38fc34cd;
    11'b01001000101: data <= 32'h2beaac82;
    11'b01001000110: data <= 32'h37e93924;
    11'b01001000111: data <= 32'h379d3cec;
    11'b01001001000: data <= 32'hb4309847;
    11'b01001001001: data <= 32'hb82cc09b;
    11'b01001001010: data <= 32'h2feec21c;
    11'b01001001011: data <= 32'h38b9bd9b;
    11'b01001001100: data <= 32'h3295383c;
    11'b01001001101: data <= 32'hb237396f;
    11'b01001001110: data <= 32'h28c8b35a;
    11'b01001001111: data <= 32'hab4cb438;
    11'b01001010000: data <= 32'hbd96392d;
    11'b01001010001: data <= 32'hc1873b5b;
    11'b01001010010: data <= 32'hc0402cf9;
    11'b01001010011: data <= 32'h33b6b873;
    11'b01001010100: data <= 32'h3f06ae9e;
    11'b01001010101: data <= 32'h3c40390c;
    11'b01001010110: data <= 32'hb2393a75;
    11'b01001010111: data <= 32'h9de13ba3;
    11'b01001011000: data <= 32'h3c493e74;
    11'b01001011001: data <= 32'h3c5a3f1e;
    11'b01001011010: data <= 32'haf3d34b6;
    11'b01001011011: data <= 32'hb9ebbf54;
    11'b01001011100: data <= 32'h2e3dc0a2;
    11'b01001011101: data <= 32'h3cc1bab6;
    11'b01001011110: data <= 32'h3d34362a;
    11'b01001011111: data <= 32'h3ab7b1c4;
    11'b01001100000: data <= 32'h388bbcdd;
    11'b01001100001: data <= 32'h28fbba22;
    11'b01001100010: data <= 32'hbd46394b;
    11'b01001100011: data <= 32'hc0f33b5d;
    11'b01001100100: data <= 32'hbf9fb711;
    11'b01001100101: data <= 32'haf13be31;
    11'b01001100110: data <= 32'h39b8bc19;
    11'b01001100111: data <= 32'hb1423458;
    11'b01001101000: data <= 32'hbb703c06;
    11'b01001101001: data <= 32'hac293d30;
    11'b01001101010: data <= 32'h3cdd3f17;
    11'b01001101011: data <= 32'h3ab43f8f;
    11'b01001101100: data <= 32'hbaba3a52;
    11'b01001101101: data <= 32'hbdc3ba18;
    11'b01001101110: data <= 32'ha63fbc38;
    11'b01001101111: data <= 32'h3ed1aaeb;
    11'b01001110000: data <= 32'h400c3631;
    11'b01001110001: data <= 32'h3d6ab8b3;
    11'b01001110010: data <= 32'h3b24bd7d;
    11'b01001110011: data <= 32'h3868b6bb;
    11'b01001110100: data <= 32'hb6183c66;
    11'b01001110101: data <= 32'hbd883ac1;
    11'b01001110110: data <= 32'hbd0ebcc2;
    11'b01001110111: data <= 32'hb48fc117;
    11'b01001111000: data <= 32'h994abf04;
    11'b01001111001: data <= 32'hba0dae3c;
    11'b01001111010: data <= 32'hbbf93930;
    11'b01001111011: data <= 32'h3025392d;
    11'b01001111100: data <= 32'h3c373bf7;
    11'b01001111101: data <= 32'h28233e17;
    11'b01001111110: data <= 32'hbfc03cd8;
    11'b01001111111: data <= 32'hc07633de;
    11'b01010000000: data <= 32'hb494aecd;
    11'b01010000001: data <= 32'h3e9f3578;
    11'b01010000010: data <= 32'h3f27359d;
    11'b01010000011: data <= 32'h3bb7b7a2;
    11'b01010000100: data <= 32'h3a95b9b6;
    11'b01010000101: data <= 32'h3cca3883;
    11'b01010000110: data <= 32'h3aac3f35;
    11'b01010000111: data <= 32'hb3263b4a;
    11'b01010001000: data <= 32'hb9a7be12;
    11'b01010001001: data <= 32'hb4f4c18f;
    11'b01010001010: data <= 32'had15bf08;
    11'b01010001011: data <= 32'hb688b415;
    11'b01010001100: data <= 32'hb4d0ae61;
    11'b01010001101: data <= 32'h38f9b901;
    11'b01010001110: data <= 32'h3b3db28e;
    11'b01010001111: data <= 32'hb9063be8;
    11'b01010010000: data <= 32'hc12d3d8e;
    11'b01010010001: data <= 32'hc1213909;
    11'b01010010010: data <= 32'hb86dab33;
    11'b01010010011: data <= 32'h3be823c6;
    11'b01010010100: data <= 32'h39412f5b;
    11'b01010010101: data <= 32'haedbb0cd;
    11'b01010010110: data <= 32'h372a30cb;
    11'b01010010111: data <= 32'h3e913de4;
    11'b01010011000: data <= 32'h3e6340aa;
    11'b01010011001: data <= 32'h33ab3ca1;
    11'b01010011010: data <= 32'hb98fbc69;
    11'b01010011011: data <= 32'hb58ebff0;
    11'b01010011100: data <= 32'h3533bbbd;
    11'b01010011101: data <= 32'h37e5aeee;
    11'b01010011110: data <= 32'h3949ba8c;
    11'b01010011111: data <= 32'h3cacbeff;
    11'b01010100000: data <= 32'h3c06bc1d;
    11'b01010100001: data <= 32'hb88b39f1;
    11'b01010100010: data <= 32'hc07f3d7f;
    11'b01010100011: data <= 32'hc04d34ed;
    11'b01010100100: data <= 32'hb922ba9c;
    11'b01010100101: data <= 32'h2d76ba8a;
    11'b01010100110: data <= 32'hb993b487;
    11'b01010100111: data <= 32'hbcaaa037;
    11'b01010101000: data <= 32'h2e923795;
    11'b01010101001: data <= 32'h3ef63e5c;
    11'b01010101010: data <= 32'h3e2a4095;
    11'b01010101011: data <= 32'hb3b43db7;
    11'b01010101100: data <= 32'hbd21b114;
    11'b01010101101: data <= 32'hb825b8d7;
    11'b01010101110: data <= 32'h39ed3075;
    11'b01010101111: data <= 32'h3ca7325a;
    11'b01010110000: data <= 32'h3c8ebc9f;
    11'b01010110001: data <= 32'h3d8dc030;
    11'b01010110010: data <= 32'h3d5ebba1;
    11'b01010110011: data <= 32'h34273c27;
    11'b01010110100: data <= 32'hbc323d61;
    11'b01010110101: data <= 32'hbccbb4f3;
    11'b01010110110: data <= 32'hb801bef2;
    11'b01010110111: data <= 32'hb855be0e;
    11'b01010111000: data <= 32'hbde6b8be;
    11'b01010111001: data <= 32'hbe1db3d2;
    11'b01010111010: data <= 32'h2fbfadb2;
    11'b01010111011: data <= 32'h3e7539c3;
    11'b01010111100: data <= 32'h3b1b3e89;
    11'b01010111101: data <= 32'hbce03e25;
    11'b01010111110: data <= 32'hc01339f4;
    11'b01010111111: data <= 32'hba153837;
    11'b01011000000: data <= 32'h3a123ad7;
    11'b01011000001: data <= 32'h3be635fe;
    11'b01011000010: data <= 32'h3965bc40;
    11'b01011000011: data <= 32'h3c40be6c;
    11'b01011000100: data <= 32'h3ec5af96;
    11'b01011000101: data <= 32'h3d733ec9;
    11'b01011000110: data <= 32'h349c3db0;
    11'b01011000111: data <= 32'hb4d6b93e;
    11'b01011001000: data <= 32'hb46dc001;
    11'b01011001001: data <= 32'hb8edbdd5;
    11'b01011001010: data <= 32'hbd3db84d;
    11'b01011001011: data <= 32'hbc0fb9d0;
    11'b01011001100: data <= 32'h386ebd01;
    11'b01011001101: data <= 32'h3dfdb930;
    11'b01011001110: data <= 32'h34073a00;
    11'b01011001111: data <= 32'hbf823dbd;
    11'b01011010000: data <= 32'hc0a93c68;
    11'b01011010001: data <= 32'hbae33a2b;
    11'b01011010010: data <= 32'h351a39fb;
    11'b01011010011: data <= 32'ha956332d;
    11'b01011010100: data <= 32'hb86eba3c;
    11'b01011010101: data <= 32'h356fba6b;
    11'b01011010110: data <= 32'h3f583a32;
    11'b01011010111: data <= 32'h40284066;
    11'b01011011000: data <= 32'h3ba23e32;
    11'b01011011001: data <= 32'ha825b6c7;
    11'b01011011010: data <= 32'hb230bd32;
    11'b01011011011: data <= 32'hb416b836;
    11'b01011011100: data <= 32'hb803ab4e;
    11'b01011011101: data <= 32'hae26bc8e;
    11'b01011011110: data <= 32'h3c57c0a0;
    11'b01011011111: data <= 32'h3e19beba;
    11'b01011100000: data <= 32'h318032b9;
    11'b01011100001: data <= 32'hbe773d08;
    11'b01011100010: data <= 32'hbf2e3a87;
    11'b01011100011: data <= 32'hb91f2fea;
    11'b01011100100: data <= 32'hb48aa113;
    11'b01011100101: data <= 32'hbd4fb129;
    11'b01011100110: data <= 32'hbf4eb8d4;
    11'b01011100111: data <= 32'hb54ab61c;
    11'b01011101000: data <= 32'h3ef03baf;
    11'b01011101001: data <= 32'h40174021;
    11'b01011101010: data <= 32'h38f83e2f;
    11'b01011101011: data <= 32'hb80e3389;
    11'b01011101100: data <= 32'hb57720cb;
    11'b01011101101: data <= 32'h313c3a5c;
    11'b01011101110: data <= 32'h332038c7;
    11'b01011101111: data <= 32'h3709bcf7;
    11'b01011110000: data <= 32'h3cf5c155;
    11'b01011110001: data <= 32'h3e84bf1c;
    11'b01011110010: data <= 32'h39e8359b;
    11'b01011110011: data <= 32'hb7da3cbc;
    11'b01011110100: data <= 32'hb90f32dc;
    11'b01011110101: data <= 32'hb06cba6b;
    11'b01011110110: data <= 32'hb936b9fa;
    11'b01011110111: data <= 32'hc034b6ec;
    11'b01011111000: data <= 32'hc0c3b941;
    11'b01011111001: data <= 32'hb817b9b6;
    11'b01011111010: data <= 32'h3e22315a;
    11'b01011111011: data <= 32'h3dab3cd9;
    11'b01011111100: data <= 32'hb5643d2b;
    11'b01011111101: data <= 32'hbd203ae4;
    11'b01011111110: data <= 32'hb8853c85;
    11'b01011111111: data <= 32'h35133ee7;
    11'b01100000000: data <= 32'h33c23c12;
    11'b01100000001: data <= 32'h2ac7bc29;
    11'b01100000010: data <= 32'h39f2c069;
    11'b01100000011: data <= 32'h3e87bbf5;
    11'b01100000100: data <= 32'h3e3b3c01;
    11'b01100000101: data <= 32'h3a9f3d03;
    11'b01100000110: data <= 32'h37fcb33d;
    11'b01100000111: data <= 32'h35fcbcea;
    11'b01100001000: data <= 32'hb8a5ba2b;
    11'b01100001001: data <= 32'hbfddb39c;
    11'b01100001010: data <= 32'hbfd2ba8f;
    11'b01100001011: data <= 32'hafa0be62;
    11'b01100001100: data <= 32'h3da1bcb4;
    11'b01100001101: data <= 32'h39bf2d3a;
    11'b01100001110: data <= 32'hbc7e3aeb;
    11'b01100001111: data <= 32'hbe9b3c28;
    11'b01100010000: data <= 32'hb8783d9d;
    11'b01100010001: data <= 32'h311c3ef9;
    11'b01100010010: data <= 32'hb8253b99;
    11'b01100010011: data <= 32'hbc91b9e8;
    11'b01100010100: data <= 32'hb33fbd77;
    11'b01100010101: data <= 32'h3db39d89;
    11'b01100010110: data <= 32'h40203e53;
    11'b01100010111: data <= 32'h3e163d38;
    11'b01100011000: data <= 32'h3b76b395;
    11'b01100011001: data <= 32'h38b6ba34;
    11'b01100011010: data <= 32'hb1d52fa3;
    11'b01100011011: data <= 32'hbc9237ae;
    11'b01100011100: data <= 32'hbbcabaf8;
    11'b01100011101: data <= 32'h37adc0d9;
    11'b01100011110: data <= 32'h3d8dc078;
    11'b01100011111: data <= 32'h36f7b943;
    11'b01100100000: data <= 32'hbc5f3807;
    11'b01100100001: data <= 32'hbcac397f;
    11'b01100100010: data <= 32'hafac3a10;
    11'b01100100011: data <= 32'had7e3bb0;
    11'b01100100100: data <= 32'hbe3c381b;
    11'b01100100101: data <= 32'hc0e0b84c;
    11'b01100100110: data <= 32'hbc81ba3f;
    11'b01100100111: data <= 32'h3c5b3647;
    11'b01100101000: data <= 32'h3fb83e0a;
    11'b01100101001: data <= 32'h3cd03c70;
    11'b01100101010: data <= 32'h379c2d0a;
    11'b01100101011: data <= 32'h36b4348b;
    11'b01100101100: data <= 32'h34043dda;
    11'b01100101101: data <= 32'hb4a13d8c;
    11'b01100101110: data <= 32'hb3e3b992;
    11'b01100101111: data <= 32'h39b4c14c;
    11'b01100110000: data <= 32'h3d57c0b6;
    11'b01100110001: data <= 32'h3972b8a4;
    11'b01100110010: data <= 32'hb2f53694;
    11'b01100110011: data <= 32'h21842c7e;
    11'b01100110100: data <= 32'h392fb440;
    11'b01100110101: data <= 32'hb08d2b66;
    11'b01100110110: data <= 32'hc05c30dc;
    11'b01100110111: data <= 32'hc20fb783;
    11'b01100111000: data <= 32'hbdaaba90;
    11'b01100111001: data <= 32'h3a93b0dc;
    11'b01100111010: data <= 32'h3d193939;
    11'b01100111011: data <= 32'h318c38b3;
    11'b01100111100: data <= 32'hb6f735ef;
    11'b01100111101: data <= 32'h2e9b3ceb;
    11'b01100111110: data <= 32'h37de40e2;
    11'b01100111111: data <= 32'ha0c13fda;
    11'b01101000000: data <= 32'hb633b612;
    11'b01101000001: data <= 32'h336cc049;
    11'b01101000010: data <= 32'h3c52be18;
    11'b01101000011: data <= 32'h3c9d3186;
    11'b01101000100: data <= 32'h3b483881;
    11'b01101000101: data <= 32'h3cceb6e8;
    11'b01101000110: data <= 32'h3d70bb5c;
    11'b01101000111: data <= 32'h2e11b292;
    11'b01101001000: data <= 32'hbfea34f3;
    11'b01101001001: data <= 32'hc127b661;
    11'b01101001010: data <= 32'hbbb2bd6d;
    11'b01101001011: data <= 32'h3a13bd29;
    11'b01101001100: data <= 32'h383fb854;
    11'b01101001101: data <= 32'hba7baceb;
    11'b01101001110: data <= 32'hbc243559;
    11'b01101001111: data <= 32'h2a6e3dae;
    11'b01101010000: data <= 32'h384b40eb;
    11'b01101010001: data <= 32'hb6f63f85;
    11'b01101010010: data <= 32'hbd78af24;
    11'b01101010011: data <= 32'hba61bd0f;
    11'b01101010100: data <= 32'h38e3b5cf;
    11'b01101010101: data <= 32'h3d9c3bc2;
    11'b01101010110: data <= 32'h3e01398a;
    11'b01101010111: data <= 32'h3ea5b8e7;
    11'b01101011000: data <= 32'h3e75ba47;
    11'b01101011001: data <= 32'h37f63762;
    11'b01101011010: data <= 32'hbc793c4c;
    11'b01101011011: data <= 32'hbdceb1a1;
    11'b01101011100: data <= 32'hb136bf97;
    11'b01101011101: data <= 32'h3aa3c075;
    11'b01101011110: data <= 32'h2ee8bd54;
    11'b01101011111: data <= 32'hbc52b848;
    11'b01101100000: data <= 32'hba44ac72;
    11'b01101100001: data <= 32'h382539de;
    11'b01101100010: data <= 32'h38813e40;
    11'b01101100011: data <= 32'hbcac3d13;
    11'b01101100100: data <= 32'hc10e9d47;
    11'b01101100101: data <= 32'hbf12b887;
    11'b01101100110: data <= 32'h2fe83511;
    11'b01101100111: data <= 32'h3cac3c8d;
    11'b01101101000: data <= 32'h3c8937de;
    11'b01101101001: data <= 32'h3c7eb875;
    11'b01101101010: data <= 32'h3d3ba97b;
    11'b01101101011: data <= 32'h3abf3ea0;
    11'b01101101100: data <= 32'hb18c4021;
    11'b01101101101: data <= 32'hb761323b;
    11'b01101101110: data <= 32'h3517bfe4;
    11'b01101101111: data <= 32'h3a63c094;
    11'b01101110000: data <= 32'h2f28bcd6;
    11'b01101110001: data <= 32'hb836b851;
    11'b01101110010: data <= 32'h337eb8f3;
    11'b01101110011: data <= 32'h3d81b5db;
    11'b01101110100: data <= 32'h39e636b4;
    11'b01101110101: data <= 32'hbe663942;
    11'b01101110110: data <= 32'hc21922de;
    11'b01101110111: data <= 32'hc019b636;
    11'b01101111000: data <= 32'haf122e1b;
    11'b01101111001: data <= 32'h3864375b;
    11'b01101111010: data <= 32'h28c0af87;
    11'b01101111011: data <= 32'h951eb829;
    11'b01101111100: data <= 32'h39fe3973;
    11'b01101111101: data <= 32'h3c0c411f;
    11'b01101111110: data <= 32'h34c14156;
    11'b01101111111: data <= 32'hb47f384a;
    11'b01110000000: data <= 32'h28aabddb;
    11'b01110000001: data <= 32'h378abd94;
    11'b01110000010: data <= 32'h3513b45c;
    11'b01110000011: data <= 32'h35a2b136;
    11'b01110000100: data <= 32'h3d5fbc26;
    11'b01110000101: data <= 32'h404cbcbe;
    11'b01110000110: data <= 32'h3c39b11c;
    11'b01110000111: data <= 32'hbd6d38be;
    11'b01110001000: data <= 32'hc113303b;
    11'b01110001001: data <= 32'hbdc7b93e;
    11'b01110001010: data <= 32'h25adba2d;
    11'b01110001011: data <= 32'haf28b924;
    11'b01110001100: data <= 32'hbc5ebaf5;
    11'b01110001101: data <= 32'hbb44b986;
    11'b01110001110: data <= 32'h374a3a52;
    11'b01110001111: data <= 32'h3c4d410b;
    11'b01110010000: data <= 32'h303140f3;
    11'b01110010001: data <= 32'hbbc6392f;
    11'b01110010010: data <= 32'hbb15b947;
    11'b01110010011: data <= 32'hae93aea6;
    11'b01110010100: data <= 32'h362f3a8f;
    11'b01110010101: data <= 32'h3a9a330a;
    11'b01110010110: data <= 32'h3f04bcd5;
    11'b01110010111: data <= 32'h40adbd2e;
    11'b01110011000: data <= 32'h3d673294;
    11'b01110011001: data <= 32'hb86a3ceb;
    11'b01110011010: data <= 32'hbd2c3766;
    11'b01110011011: data <= 32'hb5dbbbdc;
    11'b01110011100: data <= 32'h35a0be3a;
    11'b01110011101: data <= 32'hb804bd8e;
    11'b01110011110: data <= 32'hbe5ebd40;
    11'b01110011111: data <= 32'hbbbfbc2c;
    11'b01110100000: data <= 32'h3a283053;
    11'b01110100001: data <= 32'h3cce3e16;
    11'b01110100010: data <= 32'hb5db3e6f;
    11'b01110100011: data <= 32'hbfcc37fe;
    11'b01110100100: data <= 32'hbf3fa133;
    11'b01110100101: data <= 32'hb8f33a56;
    11'b01110100110: data <= 32'h309c3d3e;
    11'b01110100111: data <= 32'h375c326a;
    11'b01110101000: data <= 32'h3c83bcf0;
    11'b01110101001: data <= 32'h3f3fba68;
    11'b01110101010: data <= 32'h3dd53cc4;
    11'b01110101011: data <= 32'h35584057;
    11'b01110101100: data <= 32'hae6d3b2f;
    11'b01110101101: data <= 32'h3725bbf3;
    11'b01110101110: data <= 32'h383cbe5c;
    11'b01110101111: data <= 32'hb877bcc7;
    11'b01110110000: data <= 32'hbd2abc8f;
    11'b01110110001: data <= 32'hb1d4bd8a;
    11'b01110110010: data <= 32'h3e47bb3b;
    11'b01110110011: data <= 32'h3ddc3208;
    11'b01110110100: data <= 32'hb97e394b;
    11'b01110110101: data <= 32'hc0d33484;
    11'b01110110110: data <= 32'hc0123284;
    11'b01110110111: data <= 32'hb9ce3a9b;
    11'b01110111000: data <= 32'hb4f93b1b;
    11'b01110111001: data <= 32'hb8acb556;
    11'b01110111010: data <= 32'hb170bd36;
    11'b01110111011: data <= 32'h3b64b33a;
    11'b01110111100: data <= 32'h3d7d4005;
    11'b01110111101: data <= 32'h3a874177;
    11'b01110111110: data <= 32'h355a3ca7;
    11'b01110111111: data <= 32'h3728b8cd;
    11'b01111000000: data <= 32'h34dbb9dd;
    11'b01111000001: data <= 32'hb766ae8b;
    11'b01111000010: data <= 32'hb8bdb73d;
    11'b01111000011: data <= 32'h3a89be2b;
    11'b01111000100: data <= 32'h40a1bedc;
    11'b01111000101: data <= 32'h3f06b922;
    11'b01111000110: data <= 32'hb810349e;
    11'b01111000111: data <= 32'hbfb03447;
    11'b01111001000: data <= 32'hbd302917;
    11'b01111001001: data <= 32'hb4f9313f;
    11'b01111001010: data <= 32'hb9bfad04;
    11'b01111001011: data <= 32'hbec4bc45;
    11'b01111001100: data <= 32'hbd4bbdf7;
    11'b01111001101: data <= 32'h34caae83;
    11'b01111001110: data <= 32'h3d113fe9;
    11'b01111001111: data <= 32'h39e840db;
    11'b01111010000: data <= 32'hb02f3c1f;
    11'b01111010001: data <= 32'hb4f0a779;
    11'b01111010010: data <= 32'hb4033842;
    11'b01111010011: data <= 32'hb72f3ceb;
    11'b01111010100: data <= 32'hb0d2346b;
    11'b01111010101: data <= 32'h3cdebe0d;
    11'b01111010110: data <= 32'h40d8bf93;
    11'b01111010111: data <= 32'h3f6ab822;
    11'b01111011000: data <= 32'h2deb39cf;
    11'b01111011001: data <= 32'hb99f3884;
    11'b01111011010: data <= 32'h2266b28f;
    11'b01111011011: data <= 32'h35efb85f;
    11'b01111011100: data <= 32'hbb12ba61;
    11'b01111011101: data <= 32'hc07dbdd3;
    11'b01111011110: data <= 32'hbe8abecb;
    11'b01111011111: data <= 32'h3614b8b5;
    11'b01111100000: data <= 32'h3d573c00;
    11'b01111100001: data <= 32'h35633d63;
    11'b01111100010: data <= 32'hbbf93844;
    11'b01111100011: data <= 32'hbcc13618;
    11'b01111100100: data <= 32'hb9e73dde;
    11'b01111100101: data <= 32'hb8cd3ff0;
    11'b01111100110: data <= 32'hb6383833;
    11'b01111100111: data <= 32'h38e7bdcf;
    11'b01111101000: data <= 32'h3ecebdfd;
    11'b01111101001: data <= 32'h3e833539;
    11'b01111101010: data <= 32'h39df3e64;
    11'b01111101011: data <= 32'h38273be6;
    11'b01111101100: data <= 32'h3c66b41e;
    11'b01111101101: data <= 32'h3acfb94d;
    11'b01111101110: data <= 32'hba91b8f8;
    11'b01111101111: data <= 32'hc013bc7d;
    11'b01111110000: data <= 32'hbc14bef4;
    11'b01111110001: data <= 32'h3c53bd8e;
    11'b01111110010: data <= 32'h3e5fb5aa;
    11'b01111110011: data <= 32'h24482f98;
    11'b01111110100: data <= 32'hbe02a43c;
    11'b01111110101: data <= 32'hbdb53718;
    11'b01111110110: data <= 32'hb9c13e5e;
    11'b01111110111: data <= 32'hba5e3f0a;
    11'b01111111000: data <= 32'hbcd82fc5;
    11'b01111111001: data <= 32'hb997be0a;
    11'b01111111010: data <= 32'h3847bba2;
    11'b01111111011: data <= 32'h3cc03c99;
    11'b01111111100: data <= 32'h3c244055;
    11'b01111111101: data <= 32'h3c293ca6;
    11'b01111111110: data <= 32'h3d4facba;
    11'b01111111111: data <= 32'h3a5a98e5;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    