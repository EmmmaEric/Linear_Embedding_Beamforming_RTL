
module memory_rom_0(
CLK, rst,
Addr, CEB, Q
);

input CLK, rst;
input [10:0] Addr;
input CEB;		
output [31:0] Q;

(*rom_style = "block" *) reg [31:0] data;

always @(posedge CLK) begin
if (rst) begin
    data <= 32'd0;
end else begin
if (CEB)
case(Addr)
    11'b00000000000: data <= 32'h2f99be57;
    11'b00000000001: data <= 32'h2837ba70;
    11'b00000000010: data <= 32'hb0f63c11;
    11'b00000000011: data <= 32'hbc3e3e30;
    11'b00000000100: data <= 32'hbef3b073;
    11'b00000000101: data <= 32'hbd5bbfd8;
    11'b00000000110: data <= 32'hb8efbe99;
    11'b00000000111: data <= 32'hb87131cf;
    11'b00000001000: data <= 32'hb8b33ce5;
    11'b00000001001: data <= 32'h35283afb;
    11'b00000001010: data <= 32'h3dd138f2;
    11'b00000001011: data <= 32'h3c153d1e;
    11'b00000001100: data <= 32'hbb0e3f00;
    11'b00000001101: data <= 32'hbf6e3c1b;
    11'b00000001110: data <= 32'hb789afb5;
    11'b00000001111: data <= 32'h3e7cb850;
    11'b00000010000: data <= 32'h400ab82d;
    11'b00000010001: data <= 32'h3b2fbb2b;
    11'b00000010010: data <= 32'h355bbcae;
    11'b00000010011: data <= 32'h3bbcb489;
    11'b00000010100: data <= 32'h3cea3c81;
    11'b00000010101: data <= 32'h2ce23c3d;
    11'b00000010110: data <= 32'hbd61bacf;
    11'b00000010111: data <= 32'hbe4fc0c9;
    11'b00000011000: data <= 32'hbb80bf00;
    11'b00000011001: data <= 32'hb878ab78;
    11'b00000011010: data <= 32'hb670367e;
    11'b00000011011: data <= 32'h3330b5fa;
    11'b00000011100: data <= 32'h3a7cb622;
    11'b00000011101: data <= 32'h2e6a3c5c;
    11'b00000011110: data <= 32'hbe35409f;
    11'b00000011111: data <= 32'hc0263f0d;
    11'b00000100000: data <= 32'hb8bd349c;
    11'b00000100001: data <= 32'h3c69b6f6;
    11'b00000100010: data <= 32'h3c61b4a9;
    11'b00000100011: data <= 32'h30c6b32c;
    11'b00000100100: data <= 32'h362ab374;
    11'b00000100101: data <= 32'h3f6336bd;
    11'b00000100110: data <= 32'h40b13d3b;
    11'b00000100111: data <= 32'h3a7e3ba7;
    11'b00000101000: data <= 32'hbc52b9e9;
    11'b00000101001: data <= 32'hbd78bf9b;
    11'b00000101010: data <= 32'hb665bd44;
    11'b00000101011: data <= 32'h3314b4f9;
    11'b00000101100: data <= 32'h310ab967;
    11'b00000101101: data <= 32'h335ebef6;
    11'b00000101110: data <= 32'h36babd45;
    11'b00000101111: data <= 32'hb2723a82;
    11'b00000110000: data <= 32'hbdf9409a;
    11'b00000110001: data <= 32'hbfc23e21;
    11'b00000110010: data <= 32'hbba8b24b;
    11'b00000110011: data <= 32'h9565ba04;
    11'b00000110100: data <= 32'hb507abec;
    11'b00000110101: data <= 32'hba86373e;
    11'b00000110110: data <= 32'h33333698;
    11'b00000110111: data <= 32'h4054397c;
    11'b00000111000: data <= 32'h411c3d6d;
    11'b00000111001: data <= 32'h39ac3d38;
    11'b00000111010: data <= 32'hbc9232b3;
    11'b00000111011: data <= 32'hbba3b952;
    11'b00000111100: data <= 32'h379ab7f6;
    11'b00000111101: data <= 32'h3c57b5b6;
    11'b00000111110: data <= 32'h38adbd6e;
    11'b00000111111: data <= 32'h34adc0d6;
    11'b00001000000: data <= 32'h38cabe72;
    11'b00001000001: data <= 32'h3724396b;
    11'b00001000010: data <= 32'hb8a23f60;
    11'b00001000011: data <= 32'hbd903915;
    11'b00001000100: data <= 32'hbd01bc72;
    11'b00001000101: data <= 32'hbbf4bcbc;
    11'b00001000110: data <= 32'hbd7b2531;
    11'b00001000111: data <= 32'hbdb238ae;
    11'b00001001000: data <= 32'ha1bf312d;
    11'b00001001001: data <= 32'h3f4d30b8;
    11'b00001001010: data <= 32'h3f653c64;
    11'b00001001011: data <= 32'hac353f43;
    11'b00001001100: data <= 32'hbdd03d9b;
    11'b00001001101: data <= 32'hb92d38cb;
    11'b00001001110: data <= 32'h3bde3420;
    11'b00001001111: data <= 32'h3d11b108;
    11'b00001010000: data <= 32'h3654bd19;
    11'b00001010001: data <= 32'h33a1c026;
    11'b00001010010: data <= 32'h3ccfbc91;
    11'b00001010011: data <= 32'h3ebd3a3e;
    11'b00001010100: data <= 32'h39a83d46;
    11'b00001010101: data <= 32'hb970b255;
    11'b00001010110: data <= 32'hbcf2bead;
    11'b00001010111: data <= 32'hbd10bd0b;
    11'b00001011000: data <= 32'hbde2224e;
    11'b00001011001: data <= 32'hbd582cce;
    11'b00001011010: data <= 32'hb079bb7e;
    11'b00001011011: data <= 32'h3ca2bbfb;
    11'b00001011100: data <= 32'h3aba3893;
    11'b00001011101: data <= 32'hbac6402e;
    11'b00001011110: data <= 32'hbeae4025;
    11'b00001011111: data <= 32'hb89c3c85;
    11'b00001100000: data <= 32'h39f93816;
    11'b00001100001: data <= 32'h37d33078;
    11'b00001100010: data <= 32'hb7c4b8b1;
    11'b00001100011: data <= 32'haa62bc55;
    11'b00001100100: data <= 32'h3f19b58d;
    11'b00001100101: data <= 32'h41723bce;
    11'b00001100110: data <= 32'h3e593c3f;
    11'b00001100111: data <= 32'hb2dbb56c;
    11'b00001101000: data <= 32'hbb59bd4f;
    11'b00001101001: data <= 32'hb9b1b9b6;
    11'b00001101010: data <= 32'hb9612dbc;
    11'b00001101011: data <= 32'hb9b8b984;
    11'b00001101100: data <= 32'haf2cc06e;
    11'b00001101101: data <= 32'h3935c030;
    11'b00001101110: data <= 32'h350a2a2e;
    11'b00001101111: data <= 32'hbb853fb7;
    11'b00001110000: data <= 32'hbdc73f48;
    11'b00001110001: data <= 32'hb90b394b;
    11'b00001110010: data <= 32'ha9323184;
    11'b00001110011: data <= 32'hba9a35a2;
    11'b00001110100: data <= 32'hbe8031ab;
    11'b00001110101: data <= 32'hb7f2b3d4;
    11'b00001110110: data <= 32'h3f9a2c93;
    11'b00001110111: data <= 32'h41cf3bba;
    11'b00001111000: data <= 32'h3e243c83;
    11'b00001111001: data <= 32'hb40934c2;
    11'b00001111010: data <= 32'hb80ab22f;
    11'b00001111011: data <= 32'h334d3493;
    11'b00001111100: data <= 32'h35a835c0;
    11'b00001111101: data <= 32'hb06fbc94;
    11'b00001111110: data <= 32'had07c1b8;
    11'b00001111111: data <= 32'h38a8c0f3;
    11'b00010000000: data <= 32'h394bb146;
    11'b00010000001: data <= 32'hb0723dc4;
    11'b00010000010: data <= 32'hb9c33afa;
    11'b00010000011: data <= 32'hb8b9b61f;
    11'b00010000100: data <= 32'hba3fb659;
    11'b00010000101: data <= 32'hbf623705;
    11'b00010000110: data <= 32'hc0b73829;
    11'b00010000111: data <= 32'hbae9b2ae;
    11'b00010001000: data <= 32'h3dfeb56e;
    11'b00010001001: data <= 32'h404f3864;
    11'b00010001010: data <= 32'h39523d33;
    11'b00010001011: data <= 32'hb96e3cde;
    11'b00010001100: data <= 32'hb2973c22;
    11'b00010001101: data <= 32'h3b4f3ccc;
    11'b00010001110: data <= 32'h3a6d39f4;
    11'b00010001111: data <= 32'hb1f4bbb9;
    11'b00010010000: data <= 32'hb43ac0f7;
    11'b00010010001: data <= 32'h3ad9bfcb;
    11'b00010010010: data <= 32'h3e75263d;
    11'b00010010011: data <= 32'h3c693b6f;
    11'b00010010100: data <= 32'h3198af11;
    11'b00010010101: data <= 32'hb572bcc2;
    11'b00010010110: data <= 32'hbb5db905;
    11'b00010010111: data <= 32'hbfb03842;
    11'b00010011000: data <= 32'hc0833520;
    11'b00010011001: data <= 32'hbb92bc10;
    11'b00010011010: data <= 32'h3ab5bdb7;
    11'b00010011011: data <= 32'h3c15b198;
    11'b00010011100: data <= 32'hb5863d33;
    11'b00010011101: data <= 32'hbc393ee4;
    11'b00010011110: data <= 32'hac143e31;
    11'b00010011111: data <= 32'h3bb43df3;
    11'b00010100000: data <= 32'h35133c2e;
    11'b00010100001: data <= 32'hbbfbb452;
    11'b00010100010: data <= 32'hba04bd8b;
    11'b00010100011: data <= 32'h3c80bb95;
    11'b00010100100: data <= 32'h40eb3620;
    11'b00010100101: data <= 32'h3fe43905;
    11'b00010100110: data <= 32'h39ccb81c;
    11'b00010100111: data <= 32'h28dabc8e;
    11'b00010101000: data <= 32'hb563b157;
    11'b00010101001: data <= 32'hbc273a65;
    11'b00010101010: data <= 32'hbdd9b010;
    11'b00010101011: data <= 32'hba1ac029;
    11'b00010101100: data <= 32'h34ebc10a;
    11'b00010101101: data <= 32'h3418ba9c;
    11'b00010101110: data <= 32'hb9d63c14;
    11'b00010101111: data <= 32'hbb833da8;
    11'b00010110000: data <= 32'h2af43c0f;
    11'b00010110001: data <= 32'h37f43c11;
    11'b00010110010: data <= 32'hba203c7d;
    11'b00010110011: data <= 32'hc0443806;
    11'b00010110100: data <= 32'hbd72b552;
    11'b00010110101: data <= 32'h3c54b3b0;
    11'b00010110110: data <= 32'h411c380a;
    11'b00010110111: data <= 32'h3f81385f;
    11'b00010111000: data <= 32'h38d2b245;
    11'b00010111001: data <= 32'h359fb402;
    11'b00010111010: data <= 32'h38e03a9b;
    11'b00010111011: data <= 32'h31b03d09;
    11'b00010111100: data <= 32'hb8d6b5ec;
    11'b00010111101: data <= 32'hb89bc13b;
    11'b00010111110: data <= 32'h2fb5c1c0;
    11'b00010111111: data <= 32'h34abbc07;
    11'b00011000000: data <= 32'hb21238b6;
    11'b00011000001: data <= 32'hb37a373f;
    11'b00011000010: data <= 32'h34c7b24e;
    11'b00011000011: data <= 32'h1c7031e0;
    11'b00011000100: data <= 32'hbea03c2c;
    11'b00011000101: data <= 32'hc1b83b7b;
    11'b00011000110: data <= 32'hbf0016b8;
    11'b00011000111: data <= 32'h397eb5fe;
    11'b00011001000: data <= 32'h3f20301d;
    11'b00011001001: data <= 32'h3ae43816;
    11'b00011001010: data <= 32'habf53732;
    11'b00011001011: data <= 32'h37bb3a9c;
    11'b00011001100: data <= 32'h3d713f02;
    11'b00011001101: data <= 32'h3b493edf;
    11'b00011001110: data <= 32'hb5cab0b3;
    11'b00011001111: data <= 32'hb98cc066;
    11'b00011010000: data <= 32'h324dc075;
    11'b00011010001: data <= 32'h3b9eb8ea;
    11'b00011010010: data <= 32'h3b0e336d;
    11'b00011010011: data <= 32'h397eb8a5;
    11'b00011010100: data <= 32'h395ebd17;
    11'b00011010101: data <= 32'ha959b58d;
    11'b00011010110: data <= 32'hbeb93c28;
    11'b00011010111: data <= 32'hc1573b4f;
    11'b00011011000: data <= 32'hbeb0b808;
    11'b00011011001: data <= 32'h3121bd17;
    11'b00011011010: data <= 32'h38d3b8fa;
    11'b00011011011: data <= 32'hb6703599;
    11'b00011011100: data <= 32'hb9f33a85;
    11'b00011011101: data <= 32'h38043d1c;
    11'b00011011110: data <= 32'h3e443ff1;
    11'b00011011111: data <= 32'h39d93fa4;
    11'b00011100000: data <= 32'hbbad3723;
    11'b00011100001: data <= 32'hbccbbc40;
    11'b00011100010: data <= 32'h347dbbf2;
    11'b00011100011: data <= 32'h3e7729f5;
    11'b00011100100: data <= 32'h3eb22caf;
    11'b00011100101: data <= 32'h3cdcbc7b;
    11'b00011100110: data <= 32'h3c00be1e;
    11'b00011100111: data <= 32'h37a9afeb;
    11'b00011101000: data <= 32'hba133d3a;
    11'b00011101001: data <= 32'hbea8394e;
    11'b00011101010: data <= 32'hbccbbd6b;
    11'b00011101011: data <= 32'hb2e6c08a;
    11'b00011101100: data <= 32'hb478bd20;
    11'b00011101101: data <= 32'hbc632bd3;
    11'b00011101110: data <= 32'hbb1c3831;
    11'b00011101111: data <= 32'h38c639a4;
    11'b00011110000: data <= 32'h3d323d56;
    11'b00011110001: data <= 32'haf603ee5;
    11'b00011110010: data <= 32'hbff13c3f;
    11'b00011110011: data <= 32'hbf592dfb;
    11'b00011110100: data <= 32'h31a02654;
    11'b00011110101: data <= 32'h3ebd3749;
    11'b00011110110: data <= 32'h3e252998;
    11'b00011110111: data <= 32'h3b9abbf8;
    11'b00011111000: data <= 32'h3c5bbb31;
    11'b00011111001: data <= 32'h3d1d39eb;
    11'b00011111010: data <= 32'h385f3f39;
    11'b00011111011: data <= 32'hb8023832;
    11'b00011111100: data <= 32'hb9a3bf4a;
    11'b00011111101: data <= 32'hb524c12a;
    11'b00011111110: data <= 32'hb6dcbd70;
    11'b00011111111: data <= 32'hbaafb23d;
    11'b00100000000: data <= 32'hb565b4ff;
    11'b00100000001: data <= 32'h3b12b8b1;
    11'b00100000010: data <= 32'h3b8f32aa;
    11'b00100000011: data <= 32'hbb383d4e;
    11'b00100000100: data <= 32'hc1553d8b;
    11'b00100000101: data <= 32'hc05338cf;
    11'b00100000110: data <= 32'hae4f3207;
    11'b00100000111: data <= 32'h3c06343a;
    11'b00100001000: data <= 32'h372ea699;
    11'b00100001001: data <= 32'h22b9b81c;
    11'b00100001010: data <= 32'h3b3e295b;
    11'b00100001011: data <= 32'h3f9d3e79;
    11'b00100001100: data <= 32'h3dc3407b;
    11'b00100001101: data <= 32'h2b393974;
    11'b00100001110: data <= 32'hb8cfbde1;
    11'b00100001111: data <= 32'hb425bf7c;
    11'b00100010000: data <= 32'h2aa7b9c6;
    11'b00100010001: data <= 32'h2c62b40b;
    11'b00100010010: data <= 32'h3837bcda;
    11'b00100010011: data <= 32'h3d10bf40;
    11'b00100010100: data <= 32'h3b15b931;
    11'b00100010101: data <= 32'hbbab3c44;
    11'b00100010110: data <= 32'hc0d83d69;
    11'b00100010111: data <= 32'hbf813488;
    11'b00100011000: data <= 32'hb5a6b815;
    11'b00100011001: data <= 32'ha93bb6a1;
    11'b00100011010: data <= 32'hbba8b313;
    11'b00100011011: data <= 32'hbc02b1e7;
    11'b00100011100: data <= 32'h392037e5;
    11'b00100011101: data <= 32'h40233f3d;
    11'b00100011110: data <= 32'h3dcd4089;
    11'b00100011111: data <= 32'hb4fa3c29;
    11'b00100100000: data <= 32'hbc08b744;
    11'b00100100001: data <= 32'hb312b800;
    11'b00100100010: data <= 32'h391c3460;
    11'b00100100011: data <= 32'h3aa3aedc;
    11'b00100100100: data <= 32'h3c1bbec1;
    11'b00100100101: data <= 32'h3deac085;
    11'b00100100110: data <= 32'h3cdeb97c;
    11'b00100100111: data <= 32'hb09f3cd0;
    11'b00100101000: data <= 32'hbd2c3c95;
    11'b00100101001: data <= 32'hbc4eb756;
    11'b00100101010: data <= 32'hb6a0bdc8;
    11'b00100101011: data <= 32'hbabfbc33;
    11'b00100101100: data <= 32'hbf60b70b;
    11'b00100101101: data <= 32'hbdbfb566;
    11'b00100101110: data <= 32'h388c21d7;
    11'b00100101111: data <= 32'h3f573c37;
    11'b00100110000: data <= 32'h39e63f1c;
    11'b00100110001: data <= 32'hbcf93d5f;
    11'b00100110010: data <= 32'hbe7e38e0;
    11'b00100110011: data <= 32'hb4bf39b1;
    11'b00100110100: data <= 32'h3a5a3c00;
    11'b00100110101: data <= 32'h3a172c53;
    11'b00100110110: data <= 32'h396bbe55;
    11'b00100110111: data <= 32'h3d31bf20;
    11'b00100111000: data <= 32'h3edf2a90;
    11'b00100111001: data <= 32'h3c403eae;
    11'b00100111010: data <= 32'h2bf53c08;
    11'b00100111011: data <= 32'hb3b1bbba;
    11'b00100111100: data <= 32'hb475bf38;
    11'b00100111101: data <= 32'hbbf2bc44;
    11'b00100111110: data <= 32'hbf03b788;
    11'b00100111111: data <= 32'hbc30bb39;
    11'b00101000000: data <= 32'h3a73bcb9;
    11'b00101000001: data <= 32'h3e02b41e;
    11'b00101000010: data <= 32'haa633c18;
    11'b00101000011: data <= 32'hbfce3d93;
    11'b00101000100: data <= 32'hbfa13c66;
    11'b00101000101: data <= 32'hb6463c41;
    11'b00101000110: data <= 32'h35983c0d;
    11'b00101000111: data <= 32'hb3612cbb;
    11'b00101001000: data <= 32'hb6e9bc89;
    11'b00101001001: data <= 32'h3a11bb01;
    11'b00101001010: data <= 32'h40193b7d;
    11'b00101001011: data <= 32'h3fb0402a;
    11'b00101001100: data <= 32'h3a973c22;
    11'b00101001101: data <= 32'h2f0bba78;
    11'b00101001110: data <= 32'haeb9bcba;
    11'b00101001111: data <= 32'hb862b464;
    11'b00101010000: data <= 32'hbb57b1f5;
    11'b00101010001: data <= 32'hb276be03;
    11'b00101010010: data <= 32'h3cb6c0b8;
    11'b00101010011: data <= 32'h3d6abd52;
    11'b00101010100: data <= 32'hb432379f;
    11'b00101010101: data <= 32'hbf283cd5;
    11'b00101010110: data <= 32'hbdf53a80;
    11'b00101010111: data <= 32'hb5453774;
    11'b00101011000: data <= 32'hb66d362c;
    11'b00101011001: data <= 32'hbe55af4f;
    11'b00101011010: data <= 32'hbeafba08;
    11'b00101011011: data <= 32'h317cb4e6;
    11'b00101011100: data <= 32'h400c3cd2;
    11'b00101011101: data <= 32'h3fd04003;
    11'b00101011110: data <= 32'h38b33c6e;
    11'b00101011111: data <= 32'hb290acca;
    11'b00101100000: data <= 32'haa673031;
    11'b00101100001: data <= 32'h2b883b94;
    11'b00101100010: data <= 32'hace434e5;
    11'b00101100011: data <= 32'h35e4bf05;
    11'b00101100100: data <= 32'h3d47c1a3;
    11'b00101100101: data <= 32'h3dc6be1c;
    11'b00101100110: data <= 32'h34a2379c;
    11'b00101100111: data <= 32'hb9c63bb4;
    11'b00101101000: data <= 32'hb77f2c88;
    11'b00101101001: data <= 32'ha799b817;
    11'b00101101010: data <= 32'hbba5b4f3;
    11'b00101101011: data <= 32'hc0f3b4ae;
    11'b00101101100: data <= 32'hc096b9af;
    11'b00101101101: data <= 32'had86b867;
    11'b00101101110: data <= 32'h3ee23823;
    11'b00101101111: data <= 32'h3d013d3d;
    11'b00101110000: data <= 32'hb59e3c31;
    11'b00101110001: data <= 32'hbadf39cc;
    11'b00101110010: data <= 32'haec73d60;
    11'b00101110011: data <= 32'h35d93f8f;
    11'b00101110100: data <= 32'h2c2239b6;
    11'b00101110101: data <= 32'h2e1ebe30;
    11'b00101110110: data <= 32'h3babc0b7;
    11'b00101110111: data <= 32'h3e61ba8d;
    11'b00101111000: data <= 32'h3ce63ba3;
    11'b00101111001: data <= 32'h390b3a87;
    11'b00101111010: data <= 32'h38dbb865;
    11'b00101111011: data <= 32'h3625bc34;
    11'b00101111100: data <= 32'hbbc2b689;
    11'b00101111101: data <= 32'hc0d0b19b;
    11'b00101111110: data <= 32'hbfe2bb9d;
    11'b00101111111: data <= 32'h301ebde2;
    11'b00110000000: data <= 32'h3d83ba44;
    11'b00110000001: data <= 32'h361b34da;
    11'b00110000010: data <= 32'hbcd73a43;
    11'b00110000011: data <= 32'hbcec3c30;
    11'b00110000100: data <= 32'hadab3ee6;
    11'b00110000101: data <= 32'h32c44005;
    11'b00110000110: data <= 32'hb94f3a49;
    11'b00110000111: data <= 32'hbbf3bc4f;
    11'b00110001000: data <= 32'h3140bd94;
    11'b00110001001: data <= 32'h3e5531fa;
    11'b00110001010: data <= 32'h3f8d3dd0;
    11'b00110001011: data <= 32'h3db33a13;
    11'b00110001100: data <= 32'h3c70b92a;
    11'b00110001101: data <= 32'h3964b96f;
    11'b00110001110: data <= 32'hb7cc359f;
    11'b00110001111: data <= 32'hbe2535aa;
    11'b00110010000: data <= 32'hbc25bcc9;
    11'b00110010001: data <= 32'h38a7c0dd;
    11'b00110010010: data <= 32'h3cb4bf92;
    11'b00110010011: data <= 32'haa37b702;
    11'b00110010100: data <= 32'hbd2436d4;
    11'b00110010101: data <= 32'hbade3994;
    11'b00110010110: data <= 32'h325f3c73;
    11'b00110010111: data <= 32'hb1fe3d55;
    11'b00110011000: data <= 32'hbf253843;
    11'b00110011001: data <= 32'hc08ab952;
    11'b00110011010: data <= 32'hb934b921;
    11'b00110011011: data <= 32'h3d583972;
    11'b00110011100: data <= 32'h3f503dc4;
    11'b00110011101: data <= 32'h3cc53918;
    11'b00110011110: data <= 32'h3a50b40b;
    11'b00110011111: data <= 32'h398a3661;
    11'b00110100000: data <= 32'h30843e6f;
    11'b00110100001: data <= 32'hb8593c64;
    11'b00110100010: data <= 32'hb41abcbc;
    11'b00110100011: data <= 32'h3a70c18c;
    11'b00110100100: data <= 32'h3c67c038;
    11'b00110100101: data <= 32'h31c9b7ba;
    11'b00110100110: data <= 32'hb75131a8;
    11'b00110100111: data <= 32'h321eac3a;
    11'b00110101000: data <= 32'h3a1f22d4;
    11'b00110101001: data <= 32'hb7193730;
    11'b00110101010: data <= 32'hc1133424;
    11'b00110101011: data <= 32'hc1dbb7df;
    11'b00110101100: data <= 32'hbc03b8b0;
    11'b00110101101: data <= 32'h3bd73390;
    11'b00110101110: data <= 32'h3c6039d5;
    11'b00110101111: data <= 32'h311d34ed;
    11'b00110110000: data <= 32'ha6583340;
    11'b00110110001: data <= 32'h384c3dd1;
    11'b00110110010: data <= 32'h385c4135;
    11'b00110110011: data <= 32'hb0233e9a;
    11'b00110110100: data <= 32'hb485bafc;
    11'b00110110101: data <= 32'h3734c088;
    11'b00110110110: data <= 32'h3bf1bd55;
    11'b00110110111: data <= 32'h3a422fbf;
    11'b00110111000: data <= 32'h39c82fc5;
    11'b00110111001: data <= 32'h3d55ba12;
    11'b00110111010: data <= 32'h3d7aba2b;
    11'b00110111011: data <= 32'hb4e52e9a;
    11'b00110111100: data <= 32'hc0d1357f;
    11'b00110111101: data <= 32'hc121b7ef;
    11'b00110111110: data <= 32'hb9a3bcad;
    11'b00110111111: data <= 32'h39acbb06;
    11'b00111000000: data <= 32'h315bb59e;
    11'b00111000001: data <= 32'hbb58b200;
    11'b00111000010: data <= 32'hb91c359d;
    11'b00111000011: data <= 32'h37f23f09;
    11'b00111000100: data <= 32'h38cb416d;
    11'b00111000101: data <= 32'hb8373ec1;
    11'b00111000110: data <= 32'hbcafb724;
    11'b00111000111: data <= 32'hb6a1bd03;
    11'b00111001000: data <= 32'h39c9b03d;
    11'b00111001001: data <= 32'h3cd43ad4;
    11'b00111001010: data <= 32'h3db63094;
    11'b00111001011: data <= 32'h3f6ebc21;
    11'b00111001100: data <= 32'h3ebab9c1;
    11'b00111001101: data <= 32'h317e3930;
    11'b00111001110: data <= 32'hbdf53b6f;
    11'b00111001111: data <= 32'hbdd8b78b;
    11'b00111010000: data <= 32'ha84fbf72;
    11'b00111010001: data <= 32'h38c9bf89;
    11'b00111010010: data <= 32'hb69ebc92;
    11'b00111010011: data <= 32'hbd33b900;
    11'b00111010100: data <= 32'hb7eaa8dd;
    11'b00111010101: data <= 32'h3a8f3c64;
    11'b00111010110: data <= 32'h377f3f98;
    11'b00111010111: data <= 32'hbd703cf8;
    11'b00111011000: data <= 32'hc0a8b021;
    11'b00111011001: data <= 32'hbd36b5f0;
    11'b00111011010: data <= 32'h356f3940;
    11'b00111011011: data <= 32'h3c3e3c55;
    11'b00111011100: data <= 32'h3c9320e6;
    11'b00111011101: data <= 32'h3dbfbb2f;
    11'b00111011110: data <= 32'h3e2e2b2f;
    11'b00111011111: data <= 32'h39b03f19;
    11'b00111100000: data <= 32'hb6363f0c;
    11'b00111100001: data <= 32'hb668b468;
    11'b00111100010: data <= 32'h3715c024;
    11'b00111100011: data <= 32'h3851c017;
    11'b00111100100: data <= 32'hb6d2bc83;
    11'b00111100101: data <= 32'hba44ba27;
    11'b00111100110: data <= 32'h368ab9da;
    11'b00111100111: data <= 32'h3decae02;
    11'b00111101000: data <= 32'h36e23a05;
    11'b00111101001: data <= 32'hbfc439ac;
    11'b00111101010: data <= 32'hc1db8ccd;
    11'b00111101011: data <= 32'hbe8badff;
    11'b00111101100: data <= 32'h2852383b;
    11'b00111101101: data <= 32'h35e3384a;
    11'b00111101110: data <= 32'h2772b691;
    11'b00111101111: data <= 32'h362bb949;
    11'b00111110000: data <= 32'h3c893b4a;
    11'b00111110001: data <= 32'h3c31416a;
    11'b00111110010: data <= 32'h334140ab;
    11'b00111110011: data <= 32'haeaa298f;
    11'b00111110100: data <= 32'h3476be46;
    11'b00111110101: data <= 32'h35adbcc6;
    11'b00111110110: data <= 32'had2bb519;
    11'b00111110111: data <= 32'h3173b8b0;
    11'b00111111000: data <= 32'h3df0bd61;
    11'b00111111001: data <= 32'h4048bc3c;
    11'b00111111010: data <= 32'h390e2d4f;
    11'b00111111011: data <= 32'hbf1f389b;
    11'b00111111100: data <= 32'hc0fe2a2f;
    11'b00111111101: data <= 32'hbcadb6ac;
    11'b00111111110: data <= 32'ha767b55b;
    11'b00111111111: data <= 32'hb7aeb77f;
    11'b01000000000: data <= 32'hbcd8bbed;
    11'b01000000001: data <= 32'hb864b937;
    11'b01000000010: data <= 32'h3ad13c9a;
    11'b01000000011: data <= 32'h3c814184;
    11'b01000000100: data <= 32'h2d6f407e;
    11'b01000000101: data <= 32'hb9c334d2;
    11'b01000000110: data <= 32'hb7e5b900;
    11'b01000000111: data <= 32'ha45e30fd;
    11'b01000001000: data <= 32'h31e439ce;
    11'b01000001001: data <= 32'h3a38b4ea;
    11'b01000001010: data <= 32'h3fd9be76;
    11'b01000001011: data <= 32'h40c0bd02;
    11'b01000001100: data <= 32'h3be83565;
    11'b01000001101: data <= 32'hbb523c2e;
    11'b01000001110: data <= 32'hbd0831bf;
    11'b01000001111: data <= 32'hb26bbb50;
    11'b01000010000: data <= 32'h2ff3bcd8;
    11'b01000010001: data <= 32'hbc24bce5;
    11'b01000010010: data <= 32'hbf51bd9b;
    11'b01000010011: data <= 32'hb9b3bbca;
    11'b01000010100: data <= 32'h3c1f382e;
    11'b01000010101: data <= 32'h3c603f4c;
    11'b01000010110: data <= 32'hb83b3e1b;
    11'b01000010111: data <= 32'hbee135bb;
    11'b01000011000: data <= 32'hbd6532eb;
    11'b01000011001: data <= 32'hb6b93cb0;
    11'b01000011010: data <= 32'h2a233d1d;
    11'b01000011011: data <= 32'h3806b440;
    11'b01000011100: data <= 32'h3dc4be3f;
    11'b01000011101: data <= 32'h4000b9ae;
    11'b01000011110: data <= 32'h3d223d1c;
    11'b01000011111: data <= 32'h30693f5e;
    11'b01000100000: data <= 32'h259536e9;
    11'b01000100001: data <= 32'h38e8bc52;
    11'b01000100010: data <= 32'h3457bd6c;
    11'b01000100011: data <= 32'hbc70bc86;
    11'b01000100100: data <= 32'hbe37bd68;
    11'b01000100101: data <= 32'ha575bdce;
    11'b01000100110: data <= 32'h3e94b8f4;
    11'b01000100111: data <= 32'h3c8c3787;
    11'b01000101000: data <= 32'hbc17392d;
    11'b01000101001: data <= 32'hc08e3411;
    11'b01000101010: data <= 32'hbe813847;
    11'b01000101011: data <= 32'hb8ac3d2d;
    11'b01000101100: data <= 32'hb7863bc9;
    11'b01000101101: data <= 32'hb888b8f7;
    11'b01000101110: data <= 32'h3259bdaf;
    11'b01000101111: data <= 32'h3cfc24f2;
    11'b01000110000: data <= 32'h3d79404a;
    11'b01000110001: data <= 32'h3a2f40c1;
    11'b01000110010: data <= 32'h3897394a;
    11'b01000110011: data <= 32'h39c6b9a6;
    11'b01000110100: data <= 32'h31b2b851;
    11'b01000110101: data <= 32'hbaefb0c7;
    11'b01000110110: data <= 32'hba10babf;
    11'b01000110111: data <= 32'h3bbdbf39;
    11'b01000111000: data <= 32'h4091be59;
    11'b01000111001: data <= 32'h3d32b755;
    11'b01000111010: data <= 32'hbb8732b9;
    11'b01000111011: data <= 32'hbf7931ab;
    11'b01000111100: data <= 32'hbc0a34f5;
    11'b01000111101: data <= 32'hb59d38eb;
    11'b01000111110: data <= 32'hbc422d29;
    11'b01000111111: data <= 32'hbf32bcc1;
    11'b01001000000: data <= 32'hbbf5bdab;
    11'b01001000001: data <= 32'h391134b2;
    11'b01001000010: data <= 32'h3d22406a;
    11'b01001000011: data <= 32'h39c04056;
    11'b01001000100: data <= 32'h3153394b;
    11'b01001000101: data <= 32'h2dfa1c03;
    11'b01001000110: data <= 32'hb1c93a61;
    11'b01001000111: data <= 32'hb9243c99;
    11'b01001001000: data <= 32'hb110b2df;
    11'b01001001001: data <= 32'h3dc9bf86;
    11'b01001001010: data <= 32'h40dbbf6a;
    11'b01001001011: data <= 32'h3dc6b6f0;
    11'b01001001100: data <= 32'hb48937fa;
    11'b01001001101: data <= 32'hb9253483;
    11'b01001001110: data <= 32'h3291afa7;
    11'b01001001111: data <= 32'h3120b2d4;
    11'b01001010000: data <= 32'hbd9cb951;
    11'b01001010001: data <= 32'hc0f3be2a;
    11'b01001010010: data <= 32'hbda0be50;
    11'b01001010011: data <= 32'h38bcb118;
    11'b01001010100: data <= 32'h3ccd3d27;
    11'b01001010101: data <= 32'h31fe3cdd;
    11'b01001010110: data <= 32'hb9fb35d1;
    11'b01001010111: data <= 32'hb9e338e7;
    11'b01001011000: data <= 32'hb86f3f73;
    11'b01001011001: data <= 32'hb95f3fdf;
    11'b01001011010: data <= 32'hb4b02d89;
    11'b01001011011: data <= 32'h3b8cbefc;
    11'b01001011100: data <= 32'h3f61bd98;
    11'b01001011101: data <= 32'h3d993634;
    11'b01001011110: data <= 32'h38433cfb;
    11'b01001011111: data <= 32'h3970382f;
    11'b01001100000: data <= 32'h3d33b584;
    11'b01001100001: data <= 32'h38d5b75c;
    11'b01001100010: data <= 32'hbd75b8bd;
    11'b01001100011: data <= 32'hc094bd46;
    11'b01001100100: data <= 32'hbaecbefc;
    11'b01001100101: data <= 32'h3c82bc46;
    11'b01001100110: data <= 32'h3cf4ae8b;
    11'b01001100111: data <= 32'hb53029e3;
    11'b01001101000: data <= 32'hbd7aac71;
    11'b01001101001: data <= 32'hbc233a4e;
    11'b01001101010: data <= 32'hb8ac4026;
    11'b01001101011: data <= 32'hbb5c3f61;
    11'b01001101100: data <= 32'hbc93b0f5;
    11'b01001101101: data <= 32'hb542be63;
    11'b01001101110: data <= 32'h3a68b974;
    11'b01001101111: data <= 32'h3c863d24;
    11'b01001110000: data <= 32'h3bfc3f33;
    11'b01001110001: data <= 32'h3d48393e;
    11'b01001110010: data <= 32'h3e80b22d;
    11'b01001110011: data <= 32'h3952310e;
    11'b01001110100: data <= 32'hbc65368b;
    11'b01001110101: data <= 32'hbe1eb840;
    11'b01001110110: data <= 32'h2fa8bef3;
    11'b01001110111: data <= 32'h3f1ebf61;
    11'b01001111000: data <= 32'h3d59bc7a;
    11'b01001111001: data <= 32'hb6b4b923;
    11'b01001111010: data <= 32'hbc8ab590;
    11'b01001111011: data <= 32'hb68b382a;
    11'b01001111100: data <= 32'hadfe3dcd;
    11'b01001111101: data <= 32'hbca23bec;
    11'b01001111110: data <= 32'hc058b9ce;
    11'b01001111111: data <= 32'hbe6ebe39;
    11'b01010000000: data <= 32'hadebb468;
    11'b01010000001: data <= 32'h3a633dfe;
    11'b01010000010: data <= 32'h3afe3e5f;
    11'b01010000011: data <= 32'h3be136df;
    11'b01010000100: data <= 32'h3c4b31bf;
    11'b01010000101: data <= 32'h35333d27;
    11'b01010000110: data <= 32'hbada3f2a;
    11'b01010000111: data <= 32'hbab2365f;
    11'b01010001000: data <= 32'h39cebe17;
    11'b01010001001: data <= 32'h3fc2c007;
    11'b01010001010: data <= 32'h3d2abcb7;
    11'b01010001011: data <= 32'hac8ab799;
    11'b01010001100: data <= 32'haf19b4b4;
    11'b01010001101: data <= 32'h3b122d32;
    11'b01010001110: data <= 32'h39d43886;
    11'b01010001111: data <= 32'hbcb33092;
    11'b01010010000: data <= 32'hc174bc6e;
    11'b01010010001: data <= 32'hc03bbe44;
    11'b01010010010: data <= 32'hb4ceb739;
    11'b01010010011: data <= 32'h38f93a30;
    11'b01010010100: data <= 32'h35433896;
    11'b01010010101: data <= 32'h29fdb1c4;
    11'b01010010110: data <= 32'h317f3732;
    11'b01010010111: data <= 32'had78406d;
    11'b01010011000: data <= 32'hba31416e;
    11'b01010011001: data <= 32'hb9db3b46;
    11'b01010011010: data <= 32'h3693bcfe;
    11'b01010011011: data <= 32'h3d38be21;
    11'b01010011100: data <= 32'h3b92b5c8;
    11'b01010011101: data <= 32'h366134f7;
    11'b01010011110: data <= 32'h3c3ca4d1;
    11'b01010011111: data <= 32'h4030b30f;
    11'b01010100000: data <= 32'h3db12f85;
    11'b01010100001: data <= 32'hbb99287a;
    11'b01010100010: data <= 32'hc0febad7;
    11'b01010100011: data <= 32'hbe68bdd4;
    11'b01010100100: data <= 32'h3376bc11;
    11'b01010100101: data <= 32'h3970b74d;
    11'b01010100110: data <= 32'hb382b9c2;
    11'b01010100111: data <= 32'hb9eabb30;
    11'b01010101000: data <= 32'hb4b83650;
    11'b01010101001: data <= 32'haf0740ba;
    11'b01010101010: data <= 32'hba3e4149;
    11'b01010101011: data <= 32'hbd0239b6;
    11'b01010101100: data <= 32'hb98bbc5f;
    11'b01010101101: data <= 32'h3063ba37;
    11'b01010101110: data <= 32'h35df3954;
    11'b01010101111: data <= 32'h38c43c12;
    11'b01010110000: data <= 32'h3e80302c;
    11'b01010110001: data <= 32'h40ffb45a;
    11'b01010110010: data <= 32'h3e5236d5;
    11'b01010110011: data <= 32'hb9293ae6;
    11'b01010110100: data <= 32'hbed029e9;
    11'b01010110101: data <= 32'hb823bc7f;
    11'b01010110110: data <= 32'h3c14bdfb;
    11'b01010110111: data <= 32'h3a7abd8a;
    11'b01010111000: data <= 32'hb7ebbe0e;
    11'b01010111001: data <= 32'hba4bbd4e;
    11'b01010111010: data <= 32'h30dd2a1e;
    11'b01010111011: data <= 32'h379d3ed5;
    11'b01010111100: data <= 32'hb9953ee3;
    11'b01010111101: data <= 32'hbfdc286a;
    11'b01010111110: data <= 32'hbf7cbc5d;
    11'b01010111111: data <= 32'hbb15b39a;
    11'b01011000000: data <= 32'hb1633c8a;
    11'b01011000001: data <= 32'h35913bf0;
    11'b01011000010: data <= 32'h3d05b15d;
    11'b01011000011: data <= 32'h3fa8b28f;
    11'b01011000100: data <= 32'h3ca83cf0;
    11'b01011000101: data <= 32'hb70d4043;
    11'b01011000110: data <= 32'hbb3e3c7b;
    11'b01011000111: data <= 32'h351fb94a;
    11'b01011001000: data <= 32'h3d74bdfb;
    11'b01011001001: data <= 32'h39c0bd9f;
    11'b01011001010: data <= 32'hb6dbbd67;
    11'b01011001011: data <= 32'had58bcf8;
    11'b01011001100: data <= 32'h3d4bb5e0;
    11'b01011001101: data <= 32'h3dcc39eb;
    11'b01011001110: data <= 32'hb6e33958;
    11'b01011001111: data <= 32'hc09fb842;
    11'b01011010000: data <= 32'hc0aabc56;
    11'b01011010001: data <= 32'hbc8bb11f;
    11'b01011010010: data <= 32'hb5e539cc;
    11'b01011010011: data <= 32'hb2542ea3;
    11'b01011010100: data <= 32'h33f9bb6a;
    11'b01011010101: data <= 32'h3aafb3b7;
    11'b01011010110: data <= 32'h38983fae;
    11'b01011010111: data <= 32'hb5dc4202;
    11'b01011011000: data <= 32'hb89e3ed8;
    11'b01011011001: data <= 32'h34fbb4e4;
    11'b01011011010: data <= 32'h3afebbd5;
    11'b01011011011: data <= 32'h3388b83e;
    11'b01011011100: data <= 32'hb469b6c7;
    11'b01011011101: data <= 32'h3a99ba6e;
    11'b01011011110: data <= 32'h40f5b924;
    11'b01011011111: data <= 32'h40842e63;
    11'b01011100000: data <= 32'hac5d343a;
    11'b01011100001: data <= 32'hc003b714;
    11'b01011100010: data <= 32'hbf13badb;
    11'b01011100011: data <= 32'hb7f8b68c;
    11'b01011100100: data <= 32'hb1a2b343;
    11'b01011100101: data <= 32'hb9d3bc85;
    11'b01011100110: data <= 32'hb99bbf27;
    11'b01011100111: data <= 32'h2d8db7bf;
    11'b01011101000: data <= 32'h35ec3fd8;
    11'b01011101001: data <= 32'hb48a41c7;
    11'b01011101010: data <= 32'hba543dd0;
    11'b01011101011: data <= 32'hb804b3d8;
    11'b01011101100: data <= 32'hb33bb406;
    11'b01011101101: data <= 32'hb810391b;
    11'b01011101110: data <= 32'hb4fa3863;
    11'b01011101111: data <= 32'h3cfeb766;
    11'b01011110000: data <= 32'h41b2ba02;
    11'b01011110001: data <= 32'h40cb2fcb;
    11'b01011110010: data <= 32'h320a3a57;
    11'b01011110011: data <= 32'hbce73602;
    11'b01011110100: data <= 32'hb87db5a2;
    11'b01011110101: data <= 32'h3840b8f6;
    11'b01011110110: data <= 32'h30d0bbdd;
    11'b01011110111: data <= 32'hbc12bf98;
    11'b01011111000: data <= 32'hbc0dc07e;
    11'b01011111001: data <= 32'h3358bab1;
    11'b01011111010: data <= 32'h3ad03d2f;
    11'b01011111011: data <= 32'ha8523f71;
    11'b01011111100: data <= 32'hbcda3875;
    11'b01011111101: data <= 32'hbdecb6f4;
    11'b01011111110: data <= 32'hbcea34c0;
    11'b01011111111: data <= 32'hbc7e3d67;
    11'b01100000000: data <= 32'hb8f73aa2;
    11'b01100000001: data <= 32'h3ac2b90f;
    11'b01100000010: data <= 32'h4059baad;
    11'b01100000011: data <= 32'h3f333907;
    11'b01100000100: data <= 32'h32f53f5c;
    11'b01100000101: data <= 32'hb6e83db9;
    11'b01100000110: data <= 32'h3801336d;
    11'b01100000111: data <= 32'h3cbbb803;
    11'b01100001000: data <= 32'h32c2bb8c;
    11'b01100001001: data <= 32'hbc51beac;
    11'b01100001010: data <= 32'hb8e5c00d;
    11'b01100001011: data <= 32'h3ca4bc69;
    11'b01100001100: data <= 32'h3f343561;
    11'b01100001101: data <= 32'h362538ce;
    11'b01100001110: data <= 32'hbd90b50c;
    11'b01100001111: data <= 32'hbf6bb8cf;
    11'b01100010000: data <= 32'hbdbc37a1;
    11'b01100010001: data <= 32'hbcf33cf3;
    11'b01100010010: data <= 32'hbc3c3258;
    11'b01100010011: data <= 32'hb0f7bd6c;
    11'b01100010100: data <= 32'h3b47bc27;
    11'b01100010101: data <= 32'h3b4c3c6d;
    11'b01100010110: data <= 32'h2e704133;
    11'b01100010111: data <= 32'ha6a33ffb;
    11'b01100011000: data <= 32'h3a453876;
    11'b01100011001: data <= 32'h3bc0a9ab;
    11'b01100011010: data <= 32'hb2f6ac24;
    11'b01100011011: data <= 32'hbc66b89c;
    11'b01100011100: data <= 32'h2baabd3c;
    11'b01100011101: data <= 32'h405dbcb7;
    11'b01100011110: data <= 32'h4133b5bb;
    11'b01100011111: data <= 32'h3a28ad9b;
    11'b01100100000: data <= 32'hbc5fb82a;
    11'b01100100001: data <= 32'hbd17b746;
    11'b01100100010: data <= 32'hb941365e;
    11'b01100100011: data <= 32'hba61385b;
    11'b01100100100: data <= 32'hbd93bb0d;
    11'b01100100101: data <= 32'hbc91c070;
    11'b01100100110: data <= 32'haf4ebd69;
    11'b01100100111: data <= 32'h36513c69;
    11'b01100101000: data <= 32'h2c9c40e6;
    11'b01100101001: data <= 32'had3f3e81;
    11'b01100101010: data <= 32'h33da3696;
    11'b01100101011: data <= 32'h29c63810;
    11'b01100101100: data <= 32'hbbc23c85;
    11'b01100101101: data <= 32'hbcfc3943;
    11'b01100101110: data <= 32'h3646b923;
    11'b01100101111: data <= 32'h4100bc94;
    11'b01100110000: data <= 32'h4150b79a;
    11'b01100110001: data <= 32'h3af330e9;
    11'b01100110010: data <= 32'hb7532e0f;
    11'b01100110011: data <= 32'ha9432af8;
    11'b01100110100: data <= 32'h38f43543;
    11'b01100110101: data <= 32'hb09fad10;
    11'b01100110110: data <= 32'hbe11be5a;
    11'b01100110111: data <= 32'hbe49c142;
    11'b01100111000: data <= 32'hb443be67;
    11'b01100111001: data <= 32'h3927385e;
    11'b01100111010: data <= 32'h34f33d96;
    11'b01100111011: data <= 32'hb57f3804;
    11'b01100111100: data <= 32'hb884ae26;
    11'b01100111101: data <= 32'hbb103b01;
    11'b01100111110: data <= 32'hbe443fc5;
    11'b01100111111: data <= 32'hbe093cf4;
    11'b01101000000: data <= 32'h2b3eb867;
    11'b01101000001: data <= 32'h3f35bcc3;
    11'b01101000010: data <= 32'h3f6db054;
    11'b01101000011: data <= 32'h38c83c01;
    11'b01101000100: data <= 32'h30df3c3b;
    11'b01101000101: data <= 32'h3c6e3929;
    11'b01101000110: data <= 32'h3e4c3748;
    11'b01101000111: data <= 32'h3296ac21;
    11'b01101001000: data <= 32'hbe0abd53;
    11'b01101001001: data <= 32'hbd56c079;
    11'b01101001010: data <= 32'h3703be65;
    11'b01101001011: data <= 32'h3deab388;
    11'b01101001100: data <= 32'h39fa2b8d;
    11'b01101001101: data <= 32'hb771b968;
    11'b01101001110: data <= 32'hbb5cb89b;
    11'b01101001111: data <= 32'hbc3e3baa;
    11'b01101010000: data <= 32'hbe333ff2;
    11'b01101010001: data <= 32'hbee23ad8;
    11'b01101010010: data <= 32'hba3ebc86;
    11'b01101010011: data <= 32'h377cbdaa;
    11'b01101010100: data <= 32'h395733fd;
    11'b01101010101: data <= 32'h30ce3ed0;
    11'b01101010110: data <= 32'h36f33e5f;
    11'b01101010111: data <= 32'h3e283b0d;
    11'b01101011000: data <= 32'h3e8539ea;
    11'b01101011001: data <= 32'haa533967;
    11'b01101011010: data <= 32'hbe2eb1c1;
    11'b01101011011: data <= 32'hba40bcee;
    11'b01101011100: data <= 32'h3d77bd58;
    11'b01101011101: data <= 32'h407bba48;
    11'b01101011110: data <= 32'h3c54ba2c;
    11'b01101011111: data <= 32'hb490bcb2;
    11'b01101100000: data <= 32'hb722b91c;
    11'b01101100001: data <= 32'hb3743b04;
    11'b01101100010: data <= 32'hbac73db8;
    11'b01101100011: data <= 32'hbee7ae61;
    11'b01101100100: data <= 32'hbe6fbfcf;
    11'b01101100101: data <= 32'hb986bed9;
    11'b01101100110: data <= 32'hb13a34f9;
    11'b01101100111: data <= 32'hb00a3e83;
    11'b01101101000: data <= 32'h35a53cb8;
    11'b01101101001: data <= 32'h3c9a380c;
    11'b01101101010: data <= 32'h3ae73bdf;
    11'b01101101011: data <= 32'hb9f43ed6;
    11'b01101101100: data <= 32'hbeca3cb8;
    11'b01101101101: data <= 32'hb6e5b39f;
    11'b01101101110: data <= 32'h3eecbc13;
    11'b01101101111: data <= 32'h4088bacc;
    11'b01101110000: data <= 32'h3beeb981;
    11'b01101110001: data <= 32'h2ceeb9fe;
    11'b01101110010: data <= 32'h390db2b8;
    11'b01101110011: data <= 32'h3ca53aa1;
    11'b01101110100: data <= 32'h30733aa2;
    11'b01101110101: data <= 32'hbe25ba93;
    11'b01101110110: data <= 32'hbfd6c0ae;
    11'b01101110111: data <= 32'hbc05bf40;
    11'b01101111000: data <= 32'hb084a301;
    11'b01101111001: data <= 32'h98d139b7;
    11'b01101111010: data <= 32'h2f6caab9;
    11'b01101111011: data <= 32'h3664b547;
    11'b01101111100: data <= 32'haa833c17;
    11'b01101111101: data <= 32'hbd5040d7;
    11'b01101111110: data <= 32'hbf6e3fb4;
    11'b01101111111: data <= 32'hb8a32f6c;
    11'b01110000000: data <= 32'h3c9fbb47;
    11'b01110000001: data <= 32'h3d7ab834;
    11'b01110000010: data <= 32'h36832c94;
    11'b01110000011: data <= 32'h35b13154;
    11'b01110000100: data <= 32'h3ea935f1;
    11'b01110000101: data <= 32'h40913b28;
    11'b01110000110: data <= 32'h3a4539a1;
    11'b01110000111: data <= 32'hbd55b963;
    11'b01110001000: data <= 32'hbee2bf7a;
    11'b01110001001: data <= 32'hb694be18;
    11'b01110001010: data <= 32'h38e1b78f;
    11'b01110001011: data <= 32'h36b4b803;
    11'b01110001100: data <= 32'ha80fbd99;
    11'b01110001101: data <= 32'haa69bc86;
    11'b01110001110: data <= 32'hb51f3af6;
    11'b01110001111: data <= 32'hbd0640e3;
    11'b01110010000: data <= 32'hbf463eb1;
    11'b01110010001: data <= 32'hbc73b57d;
    11'b01110010010: data <= 32'hab0dbc67;
    11'b01110010011: data <= 32'h21ceb064;
    11'b01110010100: data <= 32'hb6213a98;
    11'b01110010101: data <= 32'h35e53a2f;
    11'b01110010110: data <= 32'h401e389a;
    11'b01110010111: data <= 32'h40f93bc7;
    11'b01110011000: data <= 32'h39883cac;
    11'b01110011001: data <= 32'hbd3835ae;
    11'b01110011010: data <= 32'hbcb3b99f;
    11'b01110011011: data <= 32'h3840bb44;
    11'b01110011100: data <= 32'h3db0b9d0;
    11'b01110011101: data <= 32'h39ebbd1f;
    11'b01110011110: data <= 32'ha1f6c021;
    11'b01110011111: data <= 32'h31eebd9b;
    11'b01110100000: data <= 32'h36313988;
    11'b01110100001: data <= 32'hb6893f96;
    11'b01110100010: data <= 32'hbde639e1;
    11'b01110100011: data <= 32'hbe84bcbf;
    11'b01110100100: data <= 32'hbc98bd92;
    11'b01110100101: data <= 32'hbc05293b;
    11'b01110100110: data <= 32'hbb4c3b9a;
    11'b01110100111: data <= 32'h30cf37a1;
    11'b01110101000: data <= 32'h3eb62d01;
    11'b01110101001: data <= 32'h3f133b1a;
    11'b01110101010: data <= 32'h1b363f8c;
    11'b01110101011: data <= 32'hbdd53e8f;
    11'b01110101100: data <= 32'hb9f337d7;
    11'b01110101101: data <= 32'h3c3cb4ba;
    11'b01110101110: data <= 32'h3e3bb8e6;
    11'b01110101111: data <= 32'h386ebcca;
    11'b01110110000: data <= 32'h2aa9bee3;
    11'b01110110001: data <= 32'h3ba5bc11;
    11'b01110110010: data <= 32'h3ecb3919;
    11'b01110110011: data <= 32'h3a423cf9;
    11'b01110110100: data <= 32'hbba8af73;
    11'b01110110101: data <= 32'hbf0cbeb8;
    11'b01110110110: data <= 32'hbdd3bdb5;
    11'b01110110111: data <= 32'hbc64a593;
    11'b01110111000: data <= 32'hbb083537;
    11'b01110111001: data <= 32'haf10b959;
    11'b01110111010: data <= 32'h3b2cbbad;
    11'b01110111011: data <= 32'h3a1138a1;
    11'b01110111100: data <= 32'hb96b40b2;
    11'b01110111101: data <= 32'hbe5040bd;
    11'b01110111110: data <= 32'hb95c3bef;
    11'b01110111111: data <= 32'h3a07a994;
    11'b01111000000: data <= 32'h3a05b38e;
    11'b01111000001: data <= 32'hb318b6c4;
    11'b01111000010: data <= 32'ha617b9f6;
    11'b01111000011: data <= 32'h3ee1b5a6;
    11'b01111000100: data <= 32'h4199397f;
    11'b01111000101: data <= 32'h3e6a3b7c;
    11'b01111000110: data <= 32'hb877b2e2;
    11'b01111000111: data <= 32'hbdbdbd3c;
    11'b01111001000: data <= 32'hbad7bbb9;
    11'b01111001001: data <= 32'hb52eb036;
    11'b01111001010: data <= 32'hb666b8e1;
    11'b01111001011: data <= 32'hb426bff6;
    11'b01111001100: data <= 32'h34d8bfda;
    11'b01111001101: data <= 32'h344131cf;
    11'b01111001110: data <= 32'hb9ba407e;
    11'b01111001111: data <= 32'hbd94403a;
    11'b01111010000: data <= 32'hbaf63865;
    11'b01111010001: data <= 32'hb18eb419;
    11'b01111010010: data <= 32'hb89a30db;
    11'b01111010011: data <= 32'hbcee370e;
    11'b01111010100: data <= 32'hb4be2b70;
    11'b01111010101: data <= 32'h3fd2a7b3;
    11'b01111010110: data <= 32'h4201393d;
    11'b01111010111: data <= 32'h3e463c60;
    11'b01111011000: data <= 32'hb810383d;
    11'b01111011001: data <= 32'hbb09b1cd;
    11'b01111011010: data <= 32'h3183afa5;
    11'b01111011011: data <= 32'h3940ac55;
    11'b01111011100: data <= 32'h2979bccc;
    11'b01111011101: data <= 32'hb50cc152;
    11'b01111011110: data <= 32'h3439c0ab;
    11'b01111011111: data <= 32'h398fac64;
    11'b01111100000: data <= 32'h2d173eae;
    11'b01111100001: data <= 32'hba963c71;
    11'b01111100010: data <= 32'hbc30b6e9;
    11'b01111100011: data <= 32'hbc38b952;
    11'b01111100100: data <= 32'hbe6a360c;
    11'b01111100101: data <= 32'hbfa03a73;
    11'b01111100110: data <= 32'hb91d27f9;
    11'b01111100111: data <= 32'h3e14b750;
    11'b01111101000: data <= 32'h407935b9;
    11'b01111101001: data <= 32'h3a3a3ddc;
    11'b01111101010: data <= 32'hba1a3e56;
    11'b01111101011: data <= 32'hb6b43c1c;
    11'b01111101100: data <= 32'h3b42396e;
    11'b01111101101: data <= 32'h3c323333;
    11'b01111101110: data <= 32'haafabc27;
    11'b01111101111: data <= 32'hb703c093;
    11'b01111110000: data <= 32'h398bbf8d;
    11'b01111110001: data <= 32'h3f0ca9d3;
    11'b01111110010: data <= 32'h3d223bfc;
    11'b01111110011: data <= 32'hadab2d10;
    11'b01111110100: data <= 32'hbb9cbcad;
    11'b01111110101: data <= 32'hbd05ba71;
    11'b01111110110: data <= 32'hbebf378c;
    11'b01111110111: data <= 32'hbf713811;
    11'b01111111000: data <= 32'hbaddbae5;
    11'b01111111001: data <= 32'h39c5be01;
    11'b01111111010: data <= 32'h3c49b1fd;
    11'b01111111011: data <= 32'hb03e3ea1;
    11'b01111111100: data <= 32'hbc03405c;
    11'b01111111101: data <= 32'hb3073e27;
    11'b01111111110: data <= 32'h3b473bc4;
    11'b01111111111: data <= 32'h380438d8;
    11'b10000000000: data <= 32'd0;
    11'b10000000001: data <= 32'd0;
    11'b10000000010: data <= 32'd0;
    11'b10000000011: data <= 32'd0;
    11'b10000000100: data <= 32'd0;
    11'b10000000101: data <= 32'd0;
    11'b10000000110: data <= 32'd0;
    11'b10000000111: data <= 32'd0;
    11'b10000001000: data <= 32'd0;
    11'b10000001001: data <= 32'd0;
    11'b10000001010: data <= 32'd0;
    11'b10000001011: data <= 32'd0;
    11'b10000001100: data <= 32'd0;
    11'b10000001101: data <= 32'd0;
    11'b10000001110: data <= 32'd0;
    11'b10000001111: data <= 32'd0;
    11'b10000010000: data <= 32'd0;
    11'b10000010001: data <= 32'd0;
    11'b10000010010: data <= 32'd0;
    11'b10000010011: data <= 32'd0;
    11'b10000010100: data <= 32'd0;
    11'b10000010101: data <= 32'd0;
    11'b10000010110: data <= 32'd0;
    11'b10000010111: data <= 32'd0;
    11'b10000011000: data <= 32'd0;
    11'b10000011001: data <= 32'd0;
    11'b10000011010: data <= 32'd0;
    11'b10000011011: data <= 32'd0;
    11'b10000011100: data <= 32'd0;
    11'b10000011101: data <= 32'd0;
    11'b10000011110: data <= 32'd0;
    11'b10000011111: data <= 32'd0;
    11'b10000100000: data <= 32'd0;
    11'b10000100001: data <= 32'd0;
    11'b10000100010: data <= 32'd0;
    11'b10000100011: data <= 32'd0;
    11'b10000100100: data <= 32'd0;
    11'b10000100101: data <= 32'd0;
    11'b10000100110: data <= 32'd0;
    11'b10000100111: data <= 32'd0;
    11'b10000101000: data <= 32'd0;
    11'b10000101001: data <= 32'd0;
    11'b10000101010: data <= 32'd0;
    11'b10000101011: data <= 32'd0;
    11'b10000101100: data <= 32'd0;
    11'b10000101101: data <= 32'd0;
    11'b10000101110: data <= 32'd0;
    11'b10000101111: data <= 32'd0;
    11'b10000110000: data <= 32'd0;
    11'b10000110001: data <= 32'd0;
    11'b10000110010: data <= 32'd0;
    11'b10000110011: data <= 32'd0;
    11'b10000110100: data <= 32'd0;
    11'b10000110101: data <= 32'd0;
    11'b10000110110: data <= 32'd0;
    11'b10000110111: data <= 32'd0;
    11'b10000111000: data <= 32'd0;
    11'b10000111001: data <= 32'd0;
    11'b10000111010: data <= 32'd0;
    11'b10000111011: data <= 32'd0;
    11'b10000111100: data <= 32'd0;
    11'b10000111101: data <= 32'd0;
    11'b10000111110: data <= 32'd0;
    11'b10000111111: data <= 32'd0;
    11'b10001000000: data <= 32'd0;
    11'b10001000001: data <= 32'd0;
    11'b10001000010: data <= 32'd0;
    11'b10001000011: data <= 32'd0;
    11'b10001000100: data <= 32'd0;
    11'b10001000101: data <= 32'd0;
    11'b10001000110: data <= 32'd0;
    11'b10001000111: data <= 32'd0;
    11'b10001001000: data <= 32'd0;
    11'b10001001001: data <= 32'd0;
    11'b10001001010: data <= 32'd0;
    11'b10001001011: data <= 32'd0;
    11'b10001001100: data <= 32'd0;
    11'b10001001101: data <= 32'd0;
    11'b10001001110: data <= 32'd0;
    11'b10001001111: data <= 32'd0;
    11'b10001010000: data <= 32'd0;
    11'b10001010001: data <= 32'd0;
    11'b10001010010: data <= 32'd0;
    11'b10001010011: data <= 32'd0;
    11'b10001010100: data <= 32'd0;
    11'b10001010101: data <= 32'd0;
    11'b10001010110: data <= 32'd0;
    11'b10001010111: data <= 32'd0;
    11'b10001011000: data <= 32'd0;
    11'b10001011001: data <= 32'd0;
    11'b10001011010: data <= 32'd0;
    11'b10001011011: data <= 32'd0;
    11'b10001011100: data <= 32'd0;
    11'b10001011101: data <= 32'd0;
    11'b10001011110: data <= 32'd0;
    11'b10001011111: data <= 32'd0;
    11'b10001100000: data <= 32'd0;
    11'b10001100001: data <= 32'd0;
    11'b10001100010: data <= 32'd0;
    11'b10001100011: data <= 32'd0;
    11'b10001100100: data <= 32'd0;
    11'b10001100101: data <= 32'd0;
    11'b10001100110: data <= 32'd0;
    11'b10001100111: data <= 32'd0;
    11'b10001101000: data <= 32'd0;
    11'b10001101001: data <= 32'd0;
    11'b10001101010: data <= 32'd0;
    11'b10001101011: data <= 32'd0;
    11'b10001101100: data <= 32'd0;
    11'b10001101101: data <= 32'd0;
    11'b10001101110: data <= 32'd0;
    11'b10001101111: data <= 32'd0;
    11'b10001110000: data <= 32'd0;
    11'b10001110001: data <= 32'd0;
    11'b10001110010: data <= 32'd0;
    11'b10001110011: data <= 32'd0;
    11'b10001110100: data <= 32'd0;
    11'b10001110101: data <= 32'd0;
    11'b10001110110: data <= 32'd0;
    11'b10001110111: data <= 32'd0;
    11'b10001111000: data <= 32'd0;
    11'b10001111001: data <= 32'd0;
    11'b10001111010: data <= 32'd0;
    11'b10001111011: data <= 32'd0;
    11'b10001111100: data <= 32'd0;
    11'b10001111101: data <= 32'd0;
    11'b10001111110: data <= 32'd0;
    11'b10001111111: data <= 32'd0;
    11'b10010000000: data <= 32'd0;
    11'b10010000001: data <= 32'd0;
    11'b10010000010: data <= 32'd0;
    11'b10010000011: data <= 32'd0;
    11'b10010000100: data <= 32'd0;
    11'b10010000101: data <= 32'd0;
    11'b10010000110: data <= 32'd0;
    11'b10010000111: data <= 32'd0;
    11'b10010001000: data <= 32'd0;
    11'b10010001001: data <= 32'd0;
    11'b10010001010: data <= 32'd0;
    11'b10010001011: data <= 32'd0;
    11'b10010001100: data <= 32'd0;
    11'b10010001101: data <= 32'd0;
    11'b10010001110: data <= 32'd0;
    11'b10010001111: data <= 32'd0;
    11'b10010010000: data <= 32'd0;
    11'b10010010001: data <= 32'd0;
    11'b10010010010: data <= 32'd0;
    11'b10010010011: data <= 32'd0;
    11'b10010010100: data <= 32'd0;
    11'b10010010101: data <= 32'd0;
    11'b10010010110: data <= 32'd0;
    11'b10010010111: data <= 32'd0;
    11'b10010011000: data <= 32'd0;
    11'b10010011001: data <= 32'd0;
    11'b10010011010: data <= 32'd0;
    11'b10010011011: data <= 32'd0;
    11'b10010011100: data <= 32'd0;
    11'b10010011101: data <= 32'd0;
    11'b10010011110: data <= 32'd0;
    11'b10010011111: data <= 32'd0;
    11'b10010100000: data <= 32'd0;
    11'b10010100001: data <= 32'd0;
    11'b10010100010: data <= 32'd0;
    11'b10010100011: data <= 32'd0;
    11'b10010100100: data <= 32'd0;
    11'b10010100101: data <= 32'd0;
    11'b10010100110: data <= 32'd0;
    11'b10010100111: data <= 32'd0;
    11'b10010101000: data <= 32'd0;
    11'b10010101001: data <= 32'd0;
    11'b10010101010: data <= 32'd0;
    11'b10010101011: data <= 32'd0;
    11'b10010101100: data <= 32'd0;
    11'b10010101101: data <= 32'd0;
    11'b10010101110: data <= 32'd0;
    11'b10010101111: data <= 32'd0;
    11'b10010110000: data <= 32'd0;
    11'b10010110001: data <= 32'd0;
    11'b10010110010: data <= 32'd0;
    11'b10010110011: data <= 32'd0;
    11'b10010110100: data <= 32'd0;
    11'b10010110101: data <= 32'd0;
    11'b10010110110: data <= 32'd0;
    11'b10010110111: data <= 32'd0;
    11'b10010111000: data <= 32'd0;
    11'b10010111001: data <= 32'd0;
    11'b10010111010: data <= 32'd0;
    11'b10010111011: data <= 32'd0;
    11'b10010111100: data <= 32'd0;
    11'b10010111101: data <= 32'd0;
    11'b10010111110: data <= 32'd0;
    11'b10010111111: data <= 32'd0;
    11'b10011000000: data <= 32'd0;
    11'b10011000001: data <= 32'd0;
    11'b10011000010: data <= 32'd0;
    11'b10011000011: data <= 32'd0;
    11'b10011000100: data <= 32'd0;
    11'b10011000101: data <= 32'd0;
    11'b10011000110: data <= 32'd0;
    11'b10011000111: data <= 32'd0;
    11'b10011001000: data <= 32'd0;
    11'b10011001001: data <= 32'd0;
    11'b10011001010: data <= 32'd0;
    11'b10011001011: data <= 32'd0;
    11'b10011001100: data <= 32'd0;
    11'b10011001101: data <= 32'd0;
    11'b10011001110: data <= 32'd0;
    11'b10011001111: data <= 32'd0;
    11'b10011010000: data <= 32'd0;
    11'b10011010001: data <= 32'd0;
    11'b10011010010: data <= 32'd0;
    11'b10011010011: data <= 32'd0;
    11'b10011010100: data <= 32'd0;
    11'b10011010101: data <= 32'd0;
    11'b10011010110: data <= 32'd0;
    11'b10011010111: data <= 32'd0;
    11'b10011011000: data <= 32'd0;
    11'b10011011001: data <= 32'd0;
    11'b10011011010: data <= 32'd0;
    11'b10011011011: data <= 32'd0;
    11'b10011011100: data <= 32'd0;
    11'b10011011101: data <= 32'd0;
    11'b10011011110: data <= 32'd0;
    11'b10011011111: data <= 32'd0;
    11'b10011100000: data <= 32'd0;
    11'b10011100001: data <= 32'd0;
    11'b10011100010: data <= 32'd0;
    11'b10011100011: data <= 32'd0;
    11'b10011100100: data <= 32'd0;
    11'b10011100101: data <= 32'd0;
    11'b10011100110: data <= 32'd0;
    11'b10011100111: data <= 32'd0;
    11'b10011101000: data <= 32'd0;
    11'b10011101001: data <= 32'd0;
    11'b10011101010: data <= 32'd0;
    11'b10011101011: data <= 32'd0;
    11'b10011101100: data <= 32'd0;
    11'b10011101101: data <= 32'd0;
    11'b10011101110: data <= 32'd0;
    11'b10011101111: data <= 32'd0;
    11'b10011110000: data <= 32'd0;
    11'b10011110001: data <= 32'd0;
    11'b10011110010: data <= 32'd0;
    11'b10011110011: data <= 32'd0;
    11'b10011110100: data <= 32'd0;
    11'b10011110101: data <= 32'd0;
    11'b10011110110: data <= 32'd0;
    11'b10011110111: data <= 32'd0;
    11'b10011111000: data <= 32'd0;
    11'b10011111001: data <= 32'd0;
    11'b10011111010: data <= 32'd0;
    11'b10011111011: data <= 32'd0;
    11'b10011111100: data <= 32'd0;
    11'b10011111101: data <= 32'd0;
    11'b10011111110: data <= 32'd0;
    11'b10011111111: data <= 32'd0;
    11'b10100000000: data <= 32'd0;
    11'b10100000001: data <= 32'd0;
    11'b10100000010: data <= 32'd0;
    11'b10100000011: data <= 32'd0;
    11'b10100000100: data <= 32'd0;
    11'b10100000101: data <= 32'd0;
    11'b10100000110: data <= 32'd0;
    11'b10100000111: data <= 32'd0;
    11'b10100001000: data <= 32'd0;
    11'b10100001001: data <= 32'd0;
    11'b10100001010: data <= 32'd0;
    11'b10100001011: data <= 32'd0;
    11'b10100001100: data <= 32'd0;
    11'b10100001101: data <= 32'd0;
    11'b10100001110: data <= 32'd0;
    11'b10100001111: data <= 32'd0;
    11'b10100010000: data <= 32'd0;
    11'b10100010001: data <= 32'd0;
    11'b10100010010: data <= 32'd0;
    11'b10100010011: data <= 32'd0;
    11'b10100010100: data <= 32'd0;
    11'b10100010101: data <= 32'd0;
    11'b10100010110: data <= 32'd0;
    11'b10100010111: data <= 32'd0;
    11'b10100011000: data <= 32'd0;
    11'b10100011001: data <= 32'd0;
    11'b10100011010: data <= 32'd0;
    11'b10100011011: data <= 32'd0;
    11'b10100011100: data <= 32'd0;
    11'b10100011101: data <= 32'd0;
    11'b10100011110: data <= 32'd0;
    11'b10100011111: data <= 32'd0;
    11'b10100100000: data <= 32'd0;
    11'b10100100001: data <= 32'd0;
    11'b10100100010: data <= 32'd0;
    11'b10100100011: data <= 32'd0;
    11'b10100100100: data <= 32'd0;
    11'b10100100101: data <= 32'd0;
    11'b10100100110: data <= 32'd0;
    11'b10100100111: data <= 32'd0;
    11'b10100101000: data <= 32'd0;
    11'b10100101001: data <= 32'd0;
    11'b10100101010: data <= 32'd0;
    11'b10100101011: data <= 32'd0;
    11'b10100101100: data <= 32'd0;
    11'b10100101101: data <= 32'd0;
    11'b10100101110: data <= 32'd0;
    11'b10100101111: data <= 32'd0;
    11'b10100110000: data <= 32'd0;
    11'b10100110001: data <= 32'd0;
    11'b10100110010: data <= 32'd0;
    11'b10100110011: data <= 32'd0;
    11'b10100110100: data <= 32'd0;
    11'b10100110101: data <= 32'd0;
    11'b10100110110: data <= 32'd0;
    11'b10100110111: data <= 32'd0;
    11'b10100111000: data <= 32'd0;
    11'b10100111001: data <= 32'd0;
    11'b10100111010: data <= 32'd0;
    11'b10100111011: data <= 32'd0;
    11'b10100111100: data <= 32'd0;
    11'b10100111101: data <= 32'd0;
    11'b10100111110: data <= 32'd0;
    11'b10100111111: data <= 32'd0;
    11'b10101000000: data <= 32'd0;
    11'b10101000001: data <= 32'd0;
    11'b10101000010: data <= 32'd0;
    11'b10101000011: data <= 32'd0;
    11'b10101000100: data <= 32'd0;
    11'b10101000101: data <= 32'd0;
    11'b10101000110: data <= 32'd0;
    11'b10101000111: data <= 32'd0;
    11'b10101001000: data <= 32'd0;
    11'b10101001001: data <= 32'd0;
    11'b10101001010: data <= 32'd0;
    11'b10101001011: data <= 32'd0;
    11'b10101001100: data <= 32'd0;
    11'b10101001101: data <= 32'd0;
    11'b10101001110: data <= 32'd0;
    11'b10101001111: data <= 32'd0;
    11'b10101010000: data <= 32'd0;
    11'b10101010001: data <= 32'd0;
    11'b10101010010: data <= 32'd0;
    11'b10101010011: data <= 32'd0;
    11'b10101010100: data <= 32'd0;
    11'b10101010101: data <= 32'd0;
    11'b10101010110: data <= 32'd0;
    11'b10101010111: data <= 32'd0;
    11'b10101011000: data <= 32'd0;
    11'b10101011001: data <= 32'd0;
    11'b10101011010: data <= 32'd0;
    11'b10101011011: data <= 32'd0;
    11'b10101011100: data <= 32'd0;
    11'b10101011101: data <= 32'd0;
    11'b10101011110: data <= 32'd0;
    11'b10101011111: data <= 32'd0;
    11'b10101100000: data <= 32'd0;
    11'b10101100001: data <= 32'd0;
    11'b10101100010: data <= 32'd0;
    11'b10101100011: data <= 32'd0;
    11'b10101100100: data <= 32'd0;
    11'b10101100101: data <= 32'd0;
    11'b10101100110: data <= 32'd0;
    11'b10101100111: data <= 32'd0;
    11'b10101101000: data <= 32'd0;
    11'b10101101001: data <= 32'd0;
    11'b10101101010: data <= 32'd0;
    11'b10101101011: data <= 32'd0;
    11'b10101101100: data <= 32'd0;
    11'b10101101101: data <= 32'd0;
    11'b10101101110: data <= 32'd0;
    11'b10101101111: data <= 32'd0;
    11'b10101110000: data <= 32'd0;
    11'b10101110001: data <= 32'd0;
    11'b10101110010: data <= 32'd0;
    11'b10101110011: data <= 32'd0;
    11'b10101110100: data <= 32'd0;
    11'b10101110101: data <= 32'd0;
    11'b10101110110: data <= 32'd0;
    11'b10101110111: data <= 32'd0;
    11'b10101111000: data <= 32'd0;
    11'b10101111001: data <= 32'd0;
    11'b10101111010: data <= 32'd0;
    11'b10101111011: data <= 32'd0;
    11'b10101111100: data <= 32'd0;
    11'b10101111101: data <= 32'd0;
    11'b10101111110: data <= 32'd0;
    11'b10101111111: data <= 32'd0;
    11'b10110000000: data <= 32'd0;
    11'b10110000001: data <= 32'd0;
    11'b10110000010: data <= 32'd0;
    11'b10110000011: data <= 32'd0;
    11'b10110000100: data <= 32'd0;
    11'b10110000101: data <= 32'd0;
    11'b10110000110: data <= 32'd0;
    11'b10110000111: data <= 32'd0;
    11'b10110001000: data <= 32'd0;
    11'b10110001001: data <= 32'd0;
    11'b10110001010: data <= 32'd0;
    11'b10110001011: data <= 32'd0;
    11'b10110001100: data <= 32'd0;
    11'b10110001101: data <= 32'd0;
    11'b10110001110: data <= 32'd0;
    11'b10110001111: data <= 32'd0;
    11'b10110010000: data <= 32'd0;
    11'b10110010001: data <= 32'd0;
    11'b10110010010: data <= 32'd0;
    11'b10110010011: data <= 32'd0;
    11'b10110010100: data <= 32'd0;
    11'b10110010101: data <= 32'd0;
    11'b10110010110: data <= 32'd0;
    11'b10110010111: data <= 32'd0;
    11'b10110011000: data <= 32'd0;
    11'b10110011001: data <= 32'd0;
    11'b10110011010: data <= 32'd0;
    11'b10110011011: data <= 32'd0;
    11'b10110011100: data <= 32'd0;
    11'b10110011101: data <= 32'd0;
    11'b10110011110: data <= 32'd0;
    11'b10110011111: data <= 32'd0;
    11'b10110100000: data <= 32'd0;
    11'b10110100001: data <= 32'd0;
    11'b10110100010: data <= 32'd0;
    11'b10110100011: data <= 32'd0;
    11'b10110100100: data <= 32'd0;
    11'b10110100101: data <= 32'd0;
    11'b10110100110: data <= 32'd0;
    11'b10110100111: data <= 32'd0;
    11'b10110101000: data <= 32'd0;
    11'b10110101001: data <= 32'd0;
    11'b10110101010: data <= 32'd0;
    11'b10110101011: data <= 32'd0;
    11'b10110101100: data <= 32'd0;
    11'b10110101101: data <= 32'd0;
    11'b10110101110: data <= 32'd0;
    11'b10110101111: data <= 32'd0;
    11'b10110110000: data <= 32'd0;
    11'b10110110001: data <= 32'd0;
    11'b10110110010: data <= 32'd0;
    11'b10110110011: data <= 32'd0;
    11'b10110110100: data <= 32'd0;
    11'b10110110101: data <= 32'd0;
    11'b10110110110: data <= 32'd0;
    11'b10110110111: data <= 32'd0;
    11'b10110111000: data <= 32'd0;
    11'b10110111001: data <= 32'd0;
    11'b10110111010: data <= 32'd0;
    11'b10110111011: data <= 32'd0;
    11'b10110111100: data <= 32'd0;
    11'b10110111101: data <= 32'd0;
    11'b10110111110: data <= 32'd0;
    11'b10110111111: data <= 32'd0;
    11'b10111000000: data <= 32'd0;
    11'b10111000001: data <= 32'd0;
    11'b10111000010: data <= 32'd0;
    11'b10111000011: data <= 32'd0;
    11'b10111000100: data <= 32'd0;
    11'b10111000101: data <= 32'd0;
    11'b10111000110: data <= 32'd0;
    11'b10111000111: data <= 32'd0;
    11'b10111001000: data <= 32'd0;
    11'b10111001001: data <= 32'd0;
    11'b10111001010: data <= 32'd0;
    11'b10111001011: data <= 32'd0;
    11'b10111001100: data <= 32'd0;
    11'b10111001101: data <= 32'd0;
    11'b10111001110: data <= 32'd0;
    11'b10111001111: data <= 32'd0;
    11'b10111010000: data <= 32'd0;
    11'b10111010001: data <= 32'd0;
    11'b10111010010: data <= 32'd0;
    11'b10111010011: data <= 32'd0;
    11'b10111010100: data <= 32'd0;
    11'b10111010101: data <= 32'd0;
    11'b10111010110: data <= 32'd0;
    11'b10111010111: data <= 32'd0;
    11'b10111011000: data <= 32'd0;
    11'b10111011001: data <= 32'd0;
    11'b10111011010: data <= 32'd0;
    11'b10111011011: data <= 32'd0;
    11'b10111011100: data <= 32'd0;
    11'b10111011101: data <= 32'd0;
    11'b10111011110: data <= 32'd0;
    11'b10111011111: data <= 32'd0;
    11'b10111100000: data <= 32'd0;
    11'b10111100001: data <= 32'd0;
    11'b10111100010: data <= 32'd0;
    11'b10111100011: data <= 32'd0;
    11'b10111100100: data <= 32'd0;
    11'b10111100101: data <= 32'd0;
    11'b10111100110: data <= 32'd0;
    11'b10111100111: data <= 32'd0;
    11'b10111101000: data <= 32'd0;
    11'b10111101001: data <= 32'd0;
    11'b10111101010: data <= 32'd0;
    11'b10111101011: data <= 32'd0;
    11'b10111101100: data <= 32'd0;
    11'b10111101101: data <= 32'd0;
    11'b10111101110: data <= 32'd0;
    11'b10111101111: data <= 32'd0;
    11'b10111110000: data <= 32'd0;
    11'b10111110001: data <= 32'd0;
    11'b10111110010: data <= 32'd0;
    11'b10111110011: data <= 32'd0;
    11'b10111110100: data <= 32'd0;
    11'b10111110101: data <= 32'd0;
    11'b10111110110: data <= 32'd0;
    11'b10111110111: data <= 32'd0;
    11'b10111111000: data <= 32'd0;
    11'b10111111001: data <= 32'd0;
    11'b10111111010: data <= 32'd0;
    11'b10111111011: data <= 32'd0;
    11'b10111111100: data <= 32'd0;
    11'b10111111101: data <= 32'd0;
    11'b10111111110: data <= 32'd0;
    11'b10111111111: data <= 32'd0;
    11'b11000000000: data <= 32'd0;
    11'b11000000001: data <= 32'd0;
    11'b11000000010: data <= 32'd0;
    11'b11000000011: data <= 32'd0;
    11'b11000000100: data <= 32'd0;
    11'b11000000101: data <= 32'd0;
    11'b11000000110: data <= 32'd0;
    11'b11000000111: data <= 32'd0;
    11'b11000001000: data <= 32'd0;
    11'b11000001001: data <= 32'd0;
    11'b11000001010: data <= 32'd0;
    11'b11000001011: data <= 32'd0;
    11'b11000001100: data <= 32'd0;
    11'b11000001101: data <= 32'd0;
    11'b11000001110: data <= 32'd0;
    11'b11000001111: data <= 32'd0;
    11'b11000010000: data <= 32'd0;
    11'b11000010001: data <= 32'd0;
    11'b11000010010: data <= 32'd0;
    11'b11000010011: data <= 32'd0;
    11'b11000010100: data <= 32'd0;
    11'b11000010101: data <= 32'd0;
    11'b11000010110: data <= 32'd0;
    11'b11000010111: data <= 32'd0;
    11'b11000011000: data <= 32'd0;
    11'b11000011001: data <= 32'd0;
    11'b11000011010: data <= 32'd0;
    11'b11000011011: data <= 32'd0;
    11'b11000011100: data <= 32'd0;
    11'b11000011101: data <= 32'd0;
    11'b11000011110: data <= 32'd0;
    11'b11000011111: data <= 32'd0;
    11'b11000100000: data <= 32'd0;
    11'b11000100001: data <= 32'd0;
    11'b11000100010: data <= 32'd0;
    11'b11000100011: data <= 32'd0;
    11'b11000100100: data <= 32'd0;
    11'b11000100101: data <= 32'd0;
    11'b11000100110: data <= 32'd0;
    11'b11000100111: data <= 32'd0;
    11'b11000101000: data <= 32'd0;
    11'b11000101001: data <= 32'd0;
    11'b11000101010: data <= 32'd0;
    11'b11000101011: data <= 32'd0;
    11'b11000101100: data <= 32'd0;
    11'b11000101101: data <= 32'd0;
    11'b11000101110: data <= 32'd0;
    11'b11000101111: data <= 32'd0;
    11'b11000110000: data <= 32'd0;
    11'b11000110001: data <= 32'd0;
    11'b11000110010: data <= 32'd0;
    11'b11000110011: data <= 32'd0;
    11'b11000110100: data <= 32'd0;
    11'b11000110101: data <= 32'd0;
    11'b11000110110: data <= 32'd0;
    11'b11000110111: data <= 32'd0;
    11'b11000111000: data <= 32'd0;
    11'b11000111001: data <= 32'd0;
    11'b11000111010: data <= 32'd0;
    11'b11000111011: data <= 32'd0;
    11'b11000111100: data <= 32'd0;
    11'b11000111101: data <= 32'd0;
    11'b11000111110: data <= 32'd0;
    11'b11000111111: data <= 32'd0;
    11'b11001000000: data <= 32'd0;
    11'b11001000001: data <= 32'd0;
    11'b11001000010: data <= 32'd0;
    11'b11001000011: data <= 32'd0;
    11'b11001000100: data <= 32'd0;
    11'b11001000101: data <= 32'd0;
    11'b11001000110: data <= 32'd0;
    11'b11001000111: data <= 32'd0;
    11'b11001001000: data <= 32'd0;
    11'b11001001001: data <= 32'd0;
    11'b11001001010: data <= 32'd0;
    11'b11001001011: data <= 32'd0;
    11'b11001001100: data <= 32'd0;
    11'b11001001101: data <= 32'd0;
    11'b11001001110: data <= 32'd0;
    11'b11001001111: data <= 32'd0;
    11'b11001010000: data <= 32'd0;
    11'b11001010001: data <= 32'd0;
    11'b11001010010: data <= 32'd0;
    11'b11001010011: data <= 32'd0;
    11'b11001010100: data <= 32'd0;
    11'b11001010101: data <= 32'd0;
    11'b11001010110: data <= 32'd0;
    11'b11001010111: data <= 32'd0;
    11'b11001011000: data <= 32'd0;
    11'b11001011001: data <= 32'd0;
    11'b11001011010: data <= 32'd0;
    11'b11001011011: data <= 32'd0;
    11'b11001011100: data <= 32'd0;
    11'b11001011101: data <= 32'd0;
    11'b11001011110: data <= 32'd0;
    11'b11001011111: data <= 32'd0;
    11'b11001100000: data <= 32'd0;
    11'b11001100001: data <= 32'd0;
    11'b11001100010: data <= 32'd0;
    11'b11001100011: data <= 32'd0;
    11'b11001100100: data <= 32'd0;
    11'b11001100101: data <= 32'd0;
    11'b11001100110: data <= 32'd0;
    11'b11001100111: data <= 32'd0;
    11'b11001101000: data <= 32'd0;
    11'b11001101001: data <= 32'd0;
    11'b11001101010: data <= 32'd0;
    11'b11001101011: data <= 32'd0;
    11'b11001101100: data <= 32'd0;
    11'b11001101101: data <= 32'd0;
    11'b11001101110: data <= 32'd0;
    11'b11001101111: data <= 32'd0;
    11'b11001110000: data <= 32'd0;
    11'b11001110001: data <= 32'd0;
    11'b11001110010: data <= 32'd0;
    11'b11001110011: data <= 32'd0;
    11'b11001110100: data <= 32'd0;
    11'b11001110101: data <= 32'd0;
    11'b11001110110: data <= 32'd0;
    11'b11001110111: data <= 32'd0;
    11'b11001111000: data <= 32'd0;
    11'b11001111001: data <= 32'd0;
    11'b11001111010: data <= 32'd0;
    11'b11001111011: data <= 32'd0;
    11'b11001111100: data <= 32'd0;
    11'b11001111101: data <= 32'd0;
    11'b11001111110: data <= 32'd0;
    11'b11001111111: data <= 32'd0;
    11'b11010000000: data <= 32'd0;
    11'b11010000001: data <= 32'd0;
    11'b11010000010: data <= 32'd0;
    11'b11010000011: data <= 32'd0;
    11'b11010000100: data <= 32'd0;
    11'b11010000101: data <= 32'd0;
    11'b11010000110: data <= 32'd0;
    11'b11010000111: data <= 32'd0;
    11'b11010001000: data <= 32'd0;
    11'b11010001001: data <= 32'd0;
    11'b11010001010: data <= 32'd0;
    11'b11010001011: data <= 32'd0;
    11'b11010001100: data <= 32'd0;
    11'b11010001101: data <= 32'd0;
    11'b11010001110: data <= 32'd0;
    11'b11010001111: data <= 32'd0;
    11'b11010010000: data <= 32'd0;
    11'b11010010001: data <= 32'd0;
    11'b11010010010: data <= 32'd0;
    11'b11010010011: data <= 32'd0;
    11'b11010010100: data <= 32'd0;
    11'b11010010101: data <= 32'd0;
    11'b11010010110: data <= 32'd0;
    11'b11010010111: data <= 32'd0;
    11'b11010011000: data <= 32'd0;
    11'b11010011001: data <= 32'd0;
    11'b11010011010: data <= 32'd0;
    11'b11010011011: data <= 32'd0;
    11'b11010011100: data <= 32'd0;
    11'b11010011101: data <= 32'd0;
    11'b11010011110: data <= 32'd0;
    11'b11010011111: data <= 32'd0;
    11'b11010100000: data <= 32'd0;
    11'b11010100001: data <= 32'd0;
    11'b11010100010: data <= 32'd0;
    11'b11010100011: data <= 32'd0;
    11'b11010100100: data <= 32'd0;
    11'b11010100101: data <= 32'd0;
    11'b11010100110: data <= 32'd0;
    11'b11010100111: data <= 32'd0;
    11'b11010101000: data <= 32'd0;
    11'b11010101001: data <= 32'd0;
    11'b11010101010: data <= 32'd0;
    11'b11010101011: data <= 32'd0;
    11'b11010101100: data <= 32'd0;
    11'b11010101101: data <= 32'd0;
    11'b11010101110: data <= 32'd0;
    11'b11010101111: data <= 32'd0;
    11'b11010110000: data <= 32'd0;
    11'b11010110001: data <= 32'd0;
    11'b11010110010: data <= 32'd0;
    11'b11010110011: data <= 32'd0;
    11'b11010110100: data <= 32'd0;
    11'b11010110101: data <= 32'd0;
    11'b11010110110: data <= 32'd0;
    11'b11010110111: data <= 32'd0;
    11'b11010111000: data <= 32'd0;
    11'b11010111001: data <= 32'd0;
    11'b11010111010: data <= 32'd0;
    11'b11010111011: data <= 32'd0;
    11'b11010111100: data <= 32'd0;
    11'b11010111101: data <= 32'd0;
    11'b11010111110: data <= 32'd0;
    11'b11010111111: data <= 32'd0;
    11'b11011000000: data <= 32'd0;
    11'b11011000001: data <= 32'd0;
    11'b11011000010: data <= 32'd0;
    11'b11011000011: data <= 32'd0;
    11'b11011000100: data <= 32'd0;
    11'b11011000101: data <= 32'd0;
    11'b11011000110: data <= 32'd0;
    11'b11011000111: data <= 32'd0;
    11'b11011001000: data <= 32'd0;
    11'b11011001001: data <= 32'd0;
    11'b11011001010: data <= 32'd0;
    11'b11011001011: data <= 32'd0;
    11'b11011001100: data <= 32'd0;
    11'b11011001101: data <= 32'd0;
    11'b11011001110: data <= 32'd0;
    11'b11011001111: data <= 32'd0;
    11'b11011010000: data <= 32'd0;
    11'b11011010001: data <= 32'd0;
    11'b11011010010: data <= 32'd0;
    11'b11011010011: data <= 32'd0;
    11'b11011010100: data <= 32'd0;
    11'b11011010101: data <= 32'd0;
    11'b11011010110: data <= 32'd0;
    11'b11011010111: data <= 32'd0;
    11'b11011011000: data <= 32'd0;
    11'b11011011001: data <= 32'd0;
    11'b11011011010: data <= 32'd0;
    11'b11011011011: data <= 32'd0;
    11'b11011011100: data <= 32'd0;
    11'b11011011101: data <= 32'd0;
    11'b11011011110: data <= 32'd0;
    11'b11011011111: data <= 32'd0;
    11'b11011100000: data <= 32'd0;
    11'b11011100001: data <= 32'd0;
    11'b11011100010: data <= 32'd0;
    11'b11011100011: data <= 32'd0;
    11'b11011100100: data <= 32'd0;
    11'b11011100101: data <= 32'd0;
    11'b11011100110: data <= 32'd0;
    11'b11011100111: data <= 32'd0;
    11'b11011101000: data <= 32'd0;
    11'b11011101001: data <= 32'd0;
    11'b11011101010: data <= 32'd0;
    11'b11011101011: data <= 32'd0;
    11'b11011101100: data <= 32'd0;
    11'b11011101101: data <= 32'd0;
    11'b11011101110: data <= 32'd0;
    11'b11011101111: data <= 32'd0;
    11'b11011110000: data <= 32'd0;
    11'b11011110001: data <= 32'd0;
    11'b11011110010: data <= 32'd0;
    11'b11011110011: data <= 32'd0;
    11'b11011110100: data <= 32'd0;
    11'b11011110101: data <= 32'd0;
    11'b11011110110: data <= 32'd0;
    11'b11011110111: data <= 32'd0;
    11'b11011111000: data <= 32'd0;
    11'b11011111001: data <= 32'd0;
    11'b11011111010: data <= 32'd0;
    11'b11011111011: data <= 32'd0;
    11'b11011111100: data <= 32'd0;
    11'b11011111101: data <= 32'd0;
    11'b11011111110: data <= 32'd0;
    11'b11011111111: data <= 32'd0;
    11'b11100000000: data <= 32'd0;
    11'b11100000001: data <= 32'd0;
    11'b11100000010: data <= 32'd0;
    11'b11100000011: data <= 32'd0;
    11'b11100000100: data <= 32'd0;
    11'b11100000101: data <= 32'd0;
    11'b11100000110: data <= 32'd0;
    11'b11100000111: data <= 32'd0;
    11'b11100001000: data <= 32'd0;
    11'b11100001001: data <= 32'd0;
    11'b11100001010: data <= 32'd0;
    11'b11100001011: data <= 32'd0;
    11'b11100001100: data <= 32'd0;
    11'b11100001101: data <= 32'd0;
    11'b11100001110: data <= 32'd0;
    11'b11100001111: data <= 32'd0;
    11'b11100010000: data <= 32'd0;
    11'b11100010001: data <= 32'd0;
    11'b11100010010: data <= 32'd0;
    11'b11100010011: data <= 32'd0;
    11'b11100010100: data <= 32'd0;
    11'b11100010101: data <= 32'd0;
    11'b11100010110: data <= 32'd0;
    11'b11100010111: data <= 32'd0;
    11'b11100011000: data <= 32'd0;
    11'b11100011001: data <= 32'd0;
    11'b11100011010: data <= 32'd0;
    11'b11100011011: data <= 32'd0;
    11'b11100011100: data <= 32'd0;
    11'b11100011101: data <= 32'd0;
    11'b11100011110: data <= 32'd0;
    11'b11100011111: data <= 32'd0;
    11'b11100100000: data <= 32'd0;
    11'b11100100001: data <= 32'd0;
    11'b11100100010: data <= 32'd0;
    11'b11100100011: data <= 32'd0;
    11'b11100100100: data <= 32'd0;
    11'b11100100101: data <= 32'd0;
    11'b11100100110: data <= 32'd0;
    11'b11100100111: data <= 32'd0;
    11'b11100101000: data <= 32'd0;
    11'b11100101001: data <= 32'd0;
    11'b11100101010: data <= 32'd0;
    11'b11100101011: data <= 32'd0;
    11'b11100101100: data <= 32'd0;
    11'b11100101101: data <= 32'd0;
    11'b11100101110: data <= 32'd0;
    11'b11100101111: data <= 32'd0;
    11'b11100110000: data <= 32'd0;
    11'b11100110001: data <= 32'd0;
    11'b11100110010: data <= 32'd0;
    11'b11100110011: data <= 32'd0;
    11'b11100110100: data <= 32'd0;
    11'b11100110101: data <= 32'd0;
    11'b11100110110: data <= 32'd0;
    11'b11100110111: data <= 32'd0;
    11'b11100111000: data <= 32'd0;
    11'b11100111001: data <= 32'd0;
    11'b11100111010: data <= 32'd0;
    11'b11100111011: data <= 32'd0;
    11'b11100111100: data <= 32'd0;
    11'b11100111101: data <= 32'd0;
    11'b11100111110: data <= 32'd0;
    11'b11100111111: data <= 32'd0;
    11'b11101000000: data <= 32'd0;
    11'b11101000001: data <= 32'd0;
    11'b11101000010: data <= 32'd0;
    11'b11101000011: data <= 32'd0;
    11'b11101000100: data <= 32'd0;
    11'b11101000101: data <= 32'd0;
    11'b11101000110: data <= 32'd0;
    11'b11101000111: data <= 32'd0;
    11'b11101001000: data <= 32'd0;
    11'b11101001001: data <= 32'd0;
    11'b11101001010: data <= 32'd0;
    11'b11101001011: data <= 32'd0;
    11'b11101001100: data <= 32'd0;
    11'b11101001101: data <= 32'd0;
    11'b11101001110: data <= 32'd0;
    11'b11101001111: data <= 32'd0;
    11'b11101010000: data <= 32'd0;
    11'b11101010001: data <= 32'd0;
    11'b11101010010: data <= 32'd0;
    11'b11101010011: data <= 32'd0;
    11'b11101010100: data <= 32'd0;
    11'b11101010101: data <= 32'd0;
    11'b11101010110: data <= 32'd0;
    11'b11101010111: data <= 32'd0;
    11'b11101011000: data <= 32'd0;
    11'b11101011001: data <= 32'd0;
    11'b11101011010: data <= 32'd0;
    11'b11101011011: data <= 32'd0;
    11'b11101011100: data <= 32'd0;
    11'b11101011101: data <= 32'd0;
    11'b11101011110: data <= 32'd0;
    11'b11101011111: data <= 32'd0;
    11'b11101100000: data <= 32'd0;
    11'b11101100001: data <= 32'd0;
    11'b11101100010: data <= 32'd0;
    11'b11101100011: data <= 32'd0;
    11'b11101100100: data <= 32'd0;
    11'b11101100101: data <= 32'd0;
    11'b11101100110: data <= 32'd0;
    11'b11101100111: data <= 32'd0;
    11'b11101101000: data <= 32'd0;
    11'b11101101001: data <= 32'd0;
    11'b11101101010: data <= 32'd0;
    11'b11101101011: data <= 32'd0;
    11'b11101101100: data <= 32'd0;
    11'b11101101101: data <= 32'd0;
    11'b11101101110: data <= 32'd0;
    11'b11101101111: data <= 32'd0;
    11'b11101110000: data <= 32'd0;
    11'b11101110001: data <= 32'd0;
    11'b11101110010: data <= 32'd0;
    11'b11101110011: data <= 32'd0;
    11'b11101110100: data <= 32'd0;
    11'b11101110101: data <= 32'd0;
    11'b11101110110: data <= 32'd0;
    11'b11101110111: data <= 32'd0;
    11'b11101111000: data <= 32'd0;
    11'b11101111001: data <= 32'd0;
    11'b11101111010: data <= 32'd0;
    11'b11101111011: data <= 32'd0;
    11'b11101111100: data <= 32'd0;
    11'b11101111101: data <= 32'd0;
    11'b11101111110: data <= 32'd0;
    11'b11101111111: data <= 32'd0;
    11'b11110000000: data <= 32'd0;
    11'b11110000001: data <= 32'd0;
    11'b11110000010: data <= 32'd0;
    11'b11110000011: data <= 32'd0;
    11'b11110000100: data <= 32'd0;
    11'b11110000101: data <= 32'd0;
    11'b11110000110: data <= 32'd0;
    11'b11110000111: data <= 32'd0;
    11'b11110001000: data <= 32'd0;
    11'b11110001001: data <= 32'd0;
    11'b11110001010: data <= 32'd0;
    11'b11110001011: data <= 32'd0;
    11'b11110001100: data <= 32'd0;
    11'b11110001101: data <= 32'd0;
    11'b11110001110: data <= 32'd0;
    11'b11110001111: data <= 32'd0;
    11'b11110010000: data <= 32'd0;
    11'b11110010001: data <= 32'd0;
    11'b11110010010: data <= 32'd0;
    11'b11110010011: data <= 32'd0;
    11'b11110010100: data <= 32'd0;
    11'b11110010101: data <= 32'd0;
    11'b11110010110: data <= 32'd0;
    11'b11110010111: data <= 32'd0;
    11'b11110011000: data <= 32'd0;
    11'b11110011001: data <= 32'd0;
    11'b11110011010: data <= 32'd0;
    11'b11110011011: data <= 32'd0;
    11'b11110011100: data <= 32'd0;
    11'b11110011101: data <= 32'd0;
    11'b11110011110: data <= 32'd0;
    11'b11110011111: data <= 32'd0;
    11'b11110100000: data <= 32'd0;
    11'b11110100001: data <= 32'd0;
    11'b11110100010: data <= 32'd0;
    11'b11110100011: data <= 32'd0;
    11'b11110100100: data <= 32'd0;
    11'b11110100101: data <= 32'd0;
    11'b11110100110: data <= 32'd0;
    11'b11110100111: data <= 32'd0;
    11'b11110101000: data <= 32'd0;
    11'b11110101001: data <= 32'd0;
    11'b11110101010: data <= 32'd0;
    11'b11110101011: data <= 32'd0;
    11'b11110101100: data <= 32'd0;
    11'b11110101101: data <= 32'd0;
    11'b11110101110: data <= 32'd0;
    11'b11110101111: data <= 32'd0;
    11'b11110110000: data <= 32'd0;
    11'b11110110001: data <= 32'd0;
    11'b11110110010: data <= 32'd0;
    11'b11110110011: data <= 32'd0;
    11'b11110110100: data <= 32'd0;
    11'b11110110101: data <= 32'd0;
    11'b11110110110: data <= 32'd0;
    11'b11110110111: data <= 32'd0;
    11'b11110111000: data <= 32'd0;
    11'b11110111001: data <= 32'd0;
    11'b11110111010: data <= 32'd0;
    11'b11110111011: data <= 32'd0;
    11'b11110111100: data <= 32'd0;
    11'b11110111101: data <= 32'd0;
    11'b11110111110: data <= 32'd0;
    11'b11110111111: data <= 32'd0;
    11'b11111000000: data <= 32'd0;
    11'b11111000001: data <= 32'd0;
    11'b11111000010: data <= 32'd0;
    11'b11111000011: data <= 32'd0;
    11'b11111000100: data <= 32'd0;
    11'b11111000101: data <= 32'd0;
    11'b11111000110: data <= 32'd0;
    11'b11111000111: data <= 32'd0;
    11'b11111001000: data <= 32'd0;
    11'b11111001001: data <= 32'd0;
    11'b11111001010: data <= 32'd0;
    11'b11111001011: data <= 32'd0;
    11'b11111001100: data <= 32'd0;
    11'b11111001101: data <= 32'd0;
    11'b11111001110: data <= 32'd0;
    11'b11111001111: data <= 32'd0;
    11'b11111010000: data <= 32'd0;
    11'b11111010001: data <= 32'd0;
    11'b11111010010: data <= 32'd0;
    11'b11111010011: data <= 32'd0;
    11'b11111010100: data <= 32'd0;
    11'b11111010101: data <= 32'd0;
    11'b11111010110: data <= 32'd0;
    11'b11111010111: data <= 32'd0;
    11'b11111011000: data <= 32'd0;
    11'b11111011001: data <= 32'd0;
    11'b11111011010: data <= 32'd0;
    11'b11111011011: data <= 32'd0;
    11'b11111011100: data <= 32'd0;
    11'b11111011101: data <= 32'd0;
    11'b11111011110: data <= 32'd0;
    11'b11111011111: data <= 32'd0;
    11'b11111100000: data <= 32'd0;
    11'b11111100001: data <= 32'd0;
    11'b11111100010: data <= 32'd0;
    11'b11111100011: data <= 32'd0;
    11'b11111100100: data <= 32'd0;
    11'b11111100101: data <= 32'd0;
    11'b11111100110: data <= 32'd0;
    11'b11111100111: data <= 32'd0;
    11'b11111101000: data <= 32'd0;
    11'b11111101001: data <= 32'd0;
    11'b11111101010: data <= 32'd0;
    11'b11111101011: data <= 32'd0;
    11'b11111101100: data <= 32'd0;
    11'b11111101101: data <= 32'd0;
    11'b11111101110: data <= 32'd0;
    11'b11111101111: data <= 32'd0;
    11'b11111110000: data <= 32'd0;
    11'b11111110001: data <= 32'd0;
    11'b11111110010: data <= 32'd0;
    11'b11111110011: data <= 32'd0;
    11'b11111110100: data <= 32'd0;
    11'b11111110101: data <= 32'd0;
    11'b11111110110: data <= 32'd0;
    11'b11111110111: data <= 32'd0;
    11'b11111111000: data <= 32'd0;
    11'b11111111001: data <= 32'd0;
    11'b11111111010: data <= 32'd0;
    11'b11111111011: data <= 32'd0;
    11'b11111111100: data <= 32'd0;
    11'b11111111101: data <= 32'd0;
    11'b11111111110: data <= 32'd0;
    11'b11111111111: data <= 32'd0;
    
endcase
end
end

assign Q = data;

endmodule

    